* NGSPICE file created from digital_top.ext - technology: sky130A

.subckt sky130_fd_sc_hs__or2b_4 VNB VPB VPWR VGND A B_N X a_676_48# a_489_392# a_81_296#
X0 VPWR a_81_296# X VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X1 X a_81_296# VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X2 a_81_296# a_676_48# VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X3 VPWR a_81_296# X VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X4 X a_81_296# VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X5 a_81_296# A VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X6 a_676_48# B_N VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 X a_81_296# VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X8 VGND A a_81_296# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X9 X a_81_296# VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X10 a_676_48# B_N VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X11 VGND a_81_296# X VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X12 VPWR A a_489_392# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13 a_489_392# A VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14 VGND a_676_48# a_81_296# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X15 a_489_392# a_676_48# a_81_296# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16 a_81_296# a_676_48# a_489_392# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17 VGND a_81_296# X VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
.ends

.subckt sky130_fd_sc_hs__buf_2 VNB VPB VPWR VGND A X a_21_260#
X0 a_21_260# A VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 VPWR a_21_260# X VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X2 VGND a_21_260# X VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X3 X a_21_260# VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X4 a_21_260# A VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X5 X a_21_260# VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
.ends

.subckt sky130_fd_sc_hs__clkbuf_4 VNB VPB VPWR VGND A X a_83_270#
X0 X a_83_270# VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1 a_83_270# A VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X2 a_83_270# A VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3 VPWR a_83_270# X VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X4 X a_83_270# VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X5 VPWR a_83_270# X VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X6 VGND a_83_270# X VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7 VGND a_83_270# X VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8 X a_83_270# VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9 X a_83_270# VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
.ends

.subckt sky130_fd_sc_hs__einvp_2 VNB VPB VPWR VGND Z A TE a_263_323# a_36_74# a_27_368#
X0 VGND TE a_36_74# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X1 VPWR TE a_263_323# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X2 a_36_74# A Z VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X3 VGND TE a_263_323# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4 Z A a_36_74# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X5 a_27_368# a_263_323# VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X6 VPWR a_263_323# a_27_368# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X7 a_27_368# A Z VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X8 a_36_74# TE VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X9 Z A a_27_368# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
.ends

.subckt sky130_fd_sc_hs__clkinv_4 VNB VPB VPWR VGND Y A
X0 VGND A Y VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1 VPWR A Y VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X2 Y A VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X3 VPWR A Y VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X4 Y A VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X5 VPWR A Y VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X6 Y A VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7 VGND A Y VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8 Y A VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9 Y A VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
.ends

.subckt sky130_fd_sc_hs__and2_2 VNB VPB VPWR VGND A B X a_31_74# a_118_74#
X0 a_118_74# A a_31_74# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X1 VPWR a_31_74# X VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X2 X a_31_74# VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X3 VGND B a_118_74# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X4 VPWR B a_31_74# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 VGND a_31_74# X VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X6 a_31_74# A VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 X a_31_74# VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
.ends

.subckt sky130_fd_sc_hs__conb_1 VNB VPB VPWR VGND LO HI a_165_290# a_21_290#
R0 HI VPWR sky130_fd_pr__res_generic_po w=510000u l=45000u
R1 VGND LO sky130_fd_pr__res_generic_po w=510000u l=45000u
.ends

.subckt sky130_fd_sc_hs__dlrtp_1 VNB VPB VPWR VGND Q GATE RESET_B D a_216_424# a_759_508#
+ a_565_74# a_27_424# a_1045_74# a_643_74# a_817_48# a_568_392# a_363_74# a_769_74#
X0 Q a_817_48# VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X1 a_1045_74# a_643_74# a_817_48# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X2 VGND a_216_424# a_363_74# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X3 a_769_74# a_216_424# a_643_74# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4 Q a_817_48# VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X5 a_643_74# a_363_74# a_565_74# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X6 VPWR a_216_424# a_363_74# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X7 VGND D a_27_424# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=550000u l=150000u
X8 a_216_424# GATE VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X9 VGND RESET_B a_1045_74# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X10 VPWR D a_27_424# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X11 VPWR RESET_B a_817_48# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 VGND a_817_48# a_769_74# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13 a_643_74# a_216_424# a_568_392# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14 a_565_74# a_27_424# VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X15 a_568_392# a_27_424# VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16 a_759_508# a_363_74# a_643_74# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17 a_817_48# a_643_74# VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X18 a_216_424# GATE VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X19 VPWR a_817_48# a_759_508# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
.ends

.subckt sky130_fd_sc_hs__inv_4 VNB VPB VPWR VGND Y A
X0 Y A VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X1 Y A VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X2 Y A VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X3 VPWR A Y VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X4 VGND A Y VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X5 Y A VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X6 VGND A Y VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X7 VPWR A Y VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
.ends

.subckt sky130_fd_sc_hs__clkbuf_2 VNB VPB VPWR VGND X A a_43_192#
X0 a_43_192# A VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X1 VPWR a_43_192# X VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X2 X a_43_192# VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3 a_43_192# A VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4 X a_43_192# VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X5 VGND a_43_192# X VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
.ends

.subckt sky130_fd_sc_hs__clkinv_2 VNB VPB VPWR VGND Y A
X0 VPWR A Y VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X1 Y A VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 VPWR A Y VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X3 Y A VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X4 VGND A Y VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
.ends

.subckt sky130_fd_sc_hs__o21bai_2 VNB VPB VPWR VGND A1 A2 B1_N Y a_27_74# a_225_74#
+ a_507_368#
X0 VGND A2 a_225_74# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X1 VGND B1_N a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X2 a_225_74# A1 VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X3 VGND A1 a_225_74# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X4 Y a_27_74# a_225_74# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X5 a_225_74# A2 VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X6 VPWR B1_N a_27_74# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 a_225_74# a_27_74# Y VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X8 VPWR a_27_74# Y VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X9 a_507_368# A2 Y VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X10 Y a_27_74# VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X11 Y A2 a_507_368# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X12 a_507_368# A1 VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X13 VPWR A1 a_507_368# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
.ends

.subckt sky130_fd_sc_hs__o21bai_4 VNB VPB VPWR VGND Y A1 A2 B1_N a_28_368# a_27_74#
+ a_828_48#
X0 VGND A1 a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X1 Y a_828_48# a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X2 VPWR A1 a_28_368# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X3 a_28_368# A2 Y VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X4 VGND A1 a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X5 Y a_828_48# VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X6 VGND A2 a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X7 a_27_74# a_828_48# Y VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X8 Y A2 a_28_368# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X9 a_28_368# A2 Y VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X10 VPWR B1_N a_828_48# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X11 VGND B1_N a_828_48# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X12 a_828_48# B1_N VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X13 a_27_74# A2 VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X14 Y A2 a_28_368# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X15 a_28_368# A1 VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X16 Y a_828_48# a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X17 VPWR A1 a_28_368# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X18 a_27_74# A1 VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X19 a_28_368# A1 VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X20 VPWR a_828_48# Y VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X21 a_27_74# a_828_48# Y VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X22 a_27_74# A1 VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X23 VGND A2 a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X24 a_27_74# A2 VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
.ends

.subckt sky130_fd_sc_hs__clkbuf_8 VNB VPB VPWR VGND X A a_125_368#
X0 VGND a_125_368# X VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1 VGND a_125_368# X VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 X a_125_368# VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X3 a_125_368# A VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4 VPWR A a_125_368# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X5 X a_125_368# VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 X a_125_368# VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7 a_125_368# A VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X8 VPWR a_125_368# X VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X9 VGND a_125_368# X VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10 X a_125_368# VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X11 VPWR a_125_368# X VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X12 X a_125_368# VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13 X a_125_368# VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X14 VGND A a_125_368# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15 VGND a_125_368# X VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16 VPWR a_125_368# X VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X17 X a_125_368# VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X18 VPWR a_125_368# X VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X19 X a_125_368# VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
.ends

.subckt sky130_fd_sc_hs__nand2_2 VNB VPB VPWR VGND Y B A a_27_74#
X0 VPWR A Y VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X1 Y A a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X2 Y A VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X3 Y B VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X4 VGND B a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X5 VPWR B Y VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X6 a_27_74# B VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X7 a_27_74# A Y VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
.ends

.subckt sky130_fd_sc_hs__xnor2_1 VNB VPB VPWR VGND A Y B a_376_368# a_112_119# a_138_385#
+ a_293_74#
X0 a_138_385# A VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X1 a_138_385# B a_112_119# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X2 VGND A a_293_74# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X3 Y B a_376_368# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X4 a_293_74# B VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X5 a_376_368# A VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X6 VPWR B a_138_385# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X7 VPWR a_138_385# Y VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X8 Y a_138_385# a_293_74# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X9 a_112_119# A VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
.ends

.subckt sky130_fd_sc_hs__nor2b_1 VNB VPB VPWR VGND B_N Y A a_278_368# a_27_112#
X0 Y A VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X1 Y a_27_112# a_278_368# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X2 a_278_368# A VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X3 VGND B_N a_27_112# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=550000u l=150000u
X4 VGND a_27_112# Y VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X5 VPWR B_N a_27_112# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
.ends

.subckt sky130_fd_sc_hs__a22o_1 VNB VPB VPWR VGND X B2 B1 A2 A1 a_222_392# a_230_79#
+ a_52_123# a_132_392#
X0 a_222_392# B1 a_230_79# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1 a_52_123# A1 a_222_392# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X2 a_222_392# B2 a_132_392# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 a_132_392# B1 a_222_392# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 X a_222_392# VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X5 VGND A2 a_52_123# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X6 X a_222_392# VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X7 VPWR A1 a_132_392# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 a_132_392# A2 VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 a_230_79# B2 VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
.ends

.subckt sky130_fd_sc_hs__nand2_1 VNB VPB VPWR VGND B Y A a_117_74#
X0 a_117_74# B VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X1 VPWR A Y VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X2 Y A a_117_74# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X3 Y B VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
.ends

.subckt sky130_fd_sc_hs__dfxtp_4 VNB VPB VPWR VGND Q D CLK a_1226_296# a_735_102#
+ a_1141_508# a_206_368# a_437_503# a_27_74# a_651_503# a_696_458# a_544_485# a_1178_124#
+ a_1034_424#
X0 a_651_503# a_27_74# a_544_485# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1 VPWR a_1226_296# Q VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X2 Q a_1226_296# VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X3 VPWR a_1226_296# Q VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X4 Q a_1226_296# VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X5 a_437_503# D VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 a_544_485# a_27_74# a_437_503# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7 VGND a_1034_424# a_1226_296# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X8 Q a_1226_296# VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X9 Q a_1226_296# VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X10 VGND CLK a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X11 a_1034_424# a_206_368# a_696_458# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=550000u l=150000u
X12 a_696_458# a_544_485# VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=550000u l=150000u
X13 a_1178_124# a_27_74# a_1034_424# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14 VGND a_696_458# a_735_102# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15 a_1141_508# a_206_368# a_1034_424# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16 a_206_368# a_27_74# VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X17 a_544_485# a_206_368# a_437_503# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18 VPWR a_696_458# a_651_503# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19 VPWR a_1226_296# a_1141_508# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20 a_696_458# a_544_485# VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X21 VGND a_1226_296# Q VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X22 VPWR a_1034_424# a_1226_296# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X23 a_206_368# a_27_74# VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X24 a_1226_296# a_1034_424# VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X25 VGND a_1226_296# a_1178_124# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X26 a_437_503# D VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X27 a_735_102# a_206_368# a_544_485# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X28 VGND a_1226_296# Q VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X29 VPWR CLK a_27_74# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X30 a_1034_424# a_27_74# a_696_458# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
.ends

.subckt sky130_fd_sc_hs__sdlclkp_2 VNB VPB VPWR VGND GCLK CLK GATE SCE a_114_112#
+ a_706_317# a_685_81# a_580_74# a_288_48# a_114_424# a_1195_374# a_708_451# a_1198_74#
+ a_318_74#
X0 a_708_451# a_288_48# a_580_74# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1 a_1195_374# CLK VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 a_706_317# a_580_74# VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X3 VPWR a_1195_374# GCLK VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X4 VGND a_1195_374# GCLK VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X5 GCLK a_1195_374# VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X6 a_114_424# SCE VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X7 a_1195_374# a_706_317# a_1198_74# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X8 a_580_74# a_288_48# a_114_112# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=550000u l=150000u
X9 a_318_74# a_288_48# VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X10 GCLK a_1195_374# VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X11 a_706_317# a_580_74# VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X12 VPWR a_706_317# a_1195_374# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13 a_685_81# a_318_74# a_580_74# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14 a_1198_74# CLK VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X15 VPWR CLK a_288_48# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X16 a_114_112# GATE a_114_424# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X17 VGND GATE a_114_112# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=550000u l=150000u
X18 a_318_74# a_288_48# VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X19 a_114_112# SCE VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=550000u l=150000u
X20 VGND CLK a_288_48# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X21 a_580_74# a_318_74# a_114_112# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X22 VPWR a_706_317# a_708_451# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23 VGND a_706_317# a_685_81# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
.ends

.subckt sky130_fd_sc_hs__and2b_2 VNB VPB VPWR VGND X B A_N a_505_74# a_27_74# a_198_48#
X0 a_198_48# a_27_74# a_505_74# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X1 VGND A_N a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=550000u l=150000u
X2 VGND a_198_48# X VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X3 VPWR a_27_74# a_198_48# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 a_198_48# B VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 VPWR a_198_48# X VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X6 a_505_74# B VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X7 X a_198_48# VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X8 X a_198_48# VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X9 VPWR A_N a_27_74# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
.ends

.subckt sky130_fd_sc_hs__clkbuf_16 VNB VPB VPWR VGND X A a_114_74#
X0 VGND a_114_74# X VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1 X a_114_74# VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 X a_114_74# VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3 a_114_74# A VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X4 X a_114_74# VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 a_114_74# A VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 VPWR a_114_74# X VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X7 a_114_74# A VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8 X a_114_74# VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X9 VPWR a_114_74# X VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X10 X a_114_74# VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X11 VGND a_114_74# X VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12 VPWR a_114_74# X VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X13 VGND A a_114_74# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14 X a_114_74# VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15 X a_114_74# VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X16 X a_114_74# VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X17 VPWR a_114_74# X VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X18 VPWR a_114_74# X VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X19 X a_114_74# VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20 X a_114_74# VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21 VPWR A a_114_74# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X22 VGND A a_114_74# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23 VGND a_114_74# X VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24 X a_114_74# VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X25 a_114_74# A VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X26 VPWR A a_114_74# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X27 VGND a_114_74# X VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X28 X a_114_74# VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X29 VGND a_114_74# X VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X30 X a_114_74# VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X31 VPWR a_114_74# X VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X32 VPWR a_114_74# X VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X33 VGND a_114_74# X VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X34 VGND a_114_74# X VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X35 X a_114_74# VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X36 X a_114_74# VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X37 VPWR a_114_74# X VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X38 VGND a_114_74# X VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X39 X a_114_74# VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
.ends

.subckt sky130_fd_sc_hs__or2_1 VNB VPB VPWR VGND B A X a_152_368# a_63_368#
X0 VPWR A a_152_368# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X1 a_152_368# B a_63_368# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X2 X a_63_368# VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X3 X a_63_368# VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X4 a_63_368# B VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=550000u l=150000u
X5 VGND A a_63_368# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=550000u l=150000u
.ends

.subckt prbs_generator_syn clk rst cke init_val[31] init_val[30] init_val[29] init_val[28]
+ init_val[27] init_val[26] init_val[25] init_val[24] init_val[23] init_val[22] init_val[21]
+ init_val[20] init_val[19] init_val[18] init_val[17] init_val[16] init_val[15] init_val[14]
+ init_val[13] init_val[12] init_val[11] init_val[10] init_val[9] init_val[8] init_val[7]
+ init_val[6] init_val[5] init_val[4] init_val[3] init_val[2] init_val[1] init_val[0]
+ eqn[31] eqn[30] eqn[29] eqn[28] eqn[27] eqn[26] eqn[25] eqn[24] eqn[23] eqn[22]
+ eqn[21] eqn[20] eqn[19] eqn[18] eqn[17] eqn[16] eqn[15] eqn[14] eqn[13] eqn[12]
+ eqn[11] eqn[10] eqn[9] eqn[8] eqn[7] eqn[6] eqn[5] eqn[4] eqn[3] eqn[2] eqn[1] eqn[0]
+ inj_err inv_chicken[1] inv_chicken[0] out DVSS DVDD sky130_fd_sc_hs__xnor2_1_1/a_293_74#
+ sky130_fd_sc_hs__a22o_1_15/X sky130_fd_sc_hs__nand2_1_35/B sky130_fd_sc_hs__xnor2_1_51/Y
+ sky130_fd_sc_hs__xnor2_1_9/A sky130_fd_sc_hs__dfxtp_4_9/CLK sky130_fd_sc_hs__dfxtp_4_47/a_27_74#
+ sky130_fd_sc_hs__dfxtp_4_37/a_1226_296# sky130_fd_sc_hs__xnor2_1_3/B sky130_fd_sc_hs__nor2b_1_7/a_27_112#
+ sky130_fd_sc_hs__xnor2_1_29/B sky130_fd_sc_hs__sdlclkp_2_1/a_580_74# sky130_fd_sc_hs__dfxtp_4_1/a_1141_508#
+ sky130_fd_sc_hs__xnor2_1_5/Y sky130_fd_sc_hs__a22o_1_41/a_230_79# sky130_fd_sc_hs__xnor2_1_61/a_138_385#
+ sky130_fd_sc_hs__a22o_1_43/a_132_392# sky130_fd_sc_hs__a22o_1_3/a_222_392# sky130_fd_sc_hs__nor2b_1_9/a_27_112#
+ sky130_fd_sc_hs__dfxtp_4_61/a_27_74# sky130_fd_sc_hs__dfxtp_4_35/a_206_368# sky130_fd_sc_hs__nand2_2_3/Y
+ sky130_fd_sc_hs__xnor2_1_25/B sky130_fd_sc_hs__nand2_1_11/a_117_74# sky130_fd_sc_hs__dfxtp_4_67/a_651_503#
+ sky130_fd_sc_hs__a22o_1_45/X sky130_fd_sc_hs__dfxtp_4_39/a_696_458# sky130_fd_sc_hs__sdlclkp_2_1/a_1198_74#
+ sky130_fd_sc_hs__dfxtp_4_45/a_1034_424# sky130_fd_sc_hs__a22o_1_17/a_222_392# sky130_fd_sc_hs__a22o_1_55/a_222_392#
+ sky130_fd_sc_hs__xnor2_1_53/Y sky130_fd_sc_hs__xnor2_1_35/A m3_13600_1651# sky130_fd_sc_hs__a22o_1_59/a_52_123#
+ sky130_fd_sc_hs__xnor2_1_5/a_293_74# sky130_fd_sc_hs__dfxtp_4_35/a_1226_296# sky130_fd_sc_hs__nand2_1_51/B
+ sky130_fd_sc_hs__dfxtp_4_5/a_651_503# sky130_fd_sc_hs__nand2_1_21/B sky130_fd_sc_hs__dfxtp_4_8/a_27_74#
+ sky130_fd_sc_hs__dfxtp_4_15/a_27_74# sky130_fd_sc_hs__and2b_2_1/X sky130_fd_sc_hs__a22o_1_13/X
+ sky130_fd_sc_hs__nand2_2_3/a_27_74# sky130_fd_sc_hs__xnor2_1_50/a_138_385# sky130_fd_sc_hs__a22o_1_33/a_132_392#
+ sky130_fd_sc_hs__xnor2_1_1/a_376_368# sky130_fd_sc_hs__dfxtp_4_25/a_206_368# sky130_fd_sc_hs__dfxtp_4_35/a_437_503#
+ sky130_fd_sc_hs__sdlclkp_2_1/a_708_451# sky130_fd_sc_hs__a22o_1_45/a_230_79# sky130_fd_sc_hs__dfxtp_4_29/a_696_458#
+ sky130_fd_sc_hs__dfxtp_4_32/a_27_74# sky130_fd_sc_hs__nor2b_1_4/Y sky130_fd_sc_hs__xnor2_1_59/a_293_74#
+ sky130_fd_sc_hs__nand2_1_47/a_117_74# sky130_fd_sc_hs__dfxtp_4_73/a_735_102# sky130_fd_sc_hs__xnor2_1_21/a_112_119#
+ sky130_fd_sc_hs__dfxtp_4_23/a_1141_508# sky130_fd_sc_hs__xnor2_1_25/a_293_74# sky130_fd_sc_hs__dfxtp_4_7/Q
+ sky130_fd_sc_hs__xnor2_1_3/a_112_119# sky130_fd_sc_hs__xnor2_1_35/B sky130_fd_sc_hs__a22o_1_51/X
+ sky130_fd_sc_hs__dfxtp_4_53/a_1178_124# sky130_fd_sc_hs__a22o_1_23/a_132_392# sky130_fd_sc_hs__nand2_1_3/B
+ sky130_fd_sc_hs__dfxtp_4_15/a_206_368# sky130_fd_sc_hs__a22o_1_63/a_132_392# sky130_fd_sc_hs__dfxtp_4_55/a_27_74#
+ sky130_fd_sc_hs__dfxtp_4_25/a_437_503# sky130_fd_sc_hs__a22o_1_41/a_52_123# sky130_fd_sc_hs__dfxtp_4_47/a_651_503#
+ sky130_fd_sc_hs__dfxtp_4_73/a_1141_508# sky130_fd_sc_hs__dfxtp_4_19/a_696_458# sky130_fd_sc_hs__dfxtp_4_57/a_696_458#
+ sky130_fd_sc_hs__a22o_1_7/X sky130_fd_sc_hs__dfxtp_4_43/a_1034_424# sky130_fd_sc_hs__xnor2_1_55/A
+ sky130_fd_sc_hs__xnor2_1_11/a_112_119# sky130_fd_sc_hs__dfxtp_4_21/a_1141_508# sky130_fd_sc_hs__a22o_1_35/a_222_392#
+ sky130_fd_sc_hs__a22o_1_49/a_230_79# sky130_fd_sc_hs__xnor2_1_67/Y sky130_fd_sc_hs__dfxtp_4_71/a_27_74#
+ sky130_fd_sc_hs__nand2_1_33/B sky130_fd_sc_hs__conb_1_1/LO sky130_fd_sc_hs__nand2_1_19/a_117_74#
+ sky130_fd_sc_hs__dfxtp_4_51/a_1178_124# sky130_fd_sc_hs__a22o_1_33/X sky130_fd_sc_hs__nand2_1_29/B
+ sky130_fd_sc_hs__xnor2_1_41/Y sky130_fd_sc_hs__a22o_1_53/a_132_392# sky130_fd_sc_hs__dfxtp_4_45/a_206_368#
+ sky130_fd_sc_hs__dfxtp_4_15/a_437_503# sky130_fd_sc_hs__dfxtp_4_37/a_651_503# sky130_fd_sc_hs__dfxtp_4_39/a_544_485#
+ sky130_fd_sc_hs__dfxtp_4_53/a_735_102# sky130_fd_sc_hs__a22o_1_45/a_52_123# sky130_fd_sc_hs__xnor2_1_1/B
+ sky130_fd_sc_hs__nand2_2_3/B sky130_fd_sc_hs__clkbuf_16_1/A sky130_fd_sc_hs__a22o_1_21/X
+ sky130_fd_sc_hs__nand2_1_25/B sky130_fd_sc_hs__xnor2_1_39/a_376_368# sky130_fd_sc_hs__a22o_1_63/X
+ m3_13600_3481# sky130_fd_sc_hs__dfxtp_4_69/a_1178_124# sky130_fd_sc_hs__xnor2_1_21/a_138_385#
+ sky130_fd_sc_hs__nor2b_1_8/Y sky130_fd_sc_hs__dfxtp_4_19/a_1178_124# sky130_fd_sc_hs__dfxtp_4_49/a_27_74#
+ sky130_fd_sc_hs__dfxtp_4_45/a_437_503# sky130_fd_sc_hs__dfxtp_4_27/a_651_503# sky130_fd_sc_hs__dfxtp_4_71/a_1141_508#
+ sky130_fd_sc_hs__dfxtp_4_65/a_651_503# sky130_fd_sc_hs__dfxtp_4_29/a_544_485# sky130_fd_sc_hs__xnor2_1_3/a_138_385#
+ sky130_fd_sc_hs__a22o_1_55/X sky130_fd_sc_hs__dfxtp_4_43/a_735_102# sky130_fd_sc_hs__dfxtp_4_41/a_1034_424#
+ sky130_fd_sc_hs__nand2_1_9/B sky130_fd_sc_hs__nor2b_1_9/Y sky130_fd_sc_hs__dfxtp_4_59/a_1034_424#
+ sky130_fd_sc_hs__dfxtp_4_39/a_1141_508# sky130_fd_sc_hs__dfxtp_4_33/a_1226_296#
+ sky130_fd_sc_hs__a22o_1_49/a_52_123# sky130_fd_sc_hs__xnor2_1_47/Y sky130_fd_sc_hs__xnor2_1_43/Y
+ sky130_fd_sc_hs__dfxtp_4_4/a_651_503# sky130_fd_sc_hs__nand2_1_49/B sky130_fd_sc_hs__xnor2_1_19/A
+ sky130_fd_sc_hs__xnor2_1_11/a_138_385# sky130_fd_sc_hs__a22o_1_5/X sky130_fd_sc_hs__dfxtp_4_63/a_206_368#
+ sky130_fd_sc_hs__dfxtp_4_17/a_651_503# sky130_fd_sc_hs__dfxtp_4_19/a_544_485# sky130_fd_sc_hs__dfxtp_4_55/a_651_503#
+ sky130_fd_sc_hs__xnor2_1_9/Y sky130_fd_sc_hs__nand2_1_17/B sky130_fd_sc_hs__dfxtp_4_57/a_544_485#
+ sky130_fd_sc_hs__dfxtp_4_67/a_696_458# sky130_fd_sc_hs__a22o_1_35/X sky130_fd_sc_hs__dfxtp_4_19/a_27_74#
+ sky130_fd_sc_hs__a22o_1_45/a_222_392# sky130_fd_sc_hs__dfxtp_4_32/a_1226_296# sky130_fd_sc_hs__nand2_1_43/B
+ sky130_fd_sc_hs__xnor2_1_25/A sky130_fd_sc_hs__dfxtp_4_1/a_206_368# sky130_fd_sc_hs__dfxtp_4_49/a_1226_296#
+ sky130_fd_sc_hs__xnor2_1_1/a_112_119# sky130_fd_sc_hs__or2_1_1/X sky130_fd_sc_hs__xnor2_1_59/a_376_368#
+ sky130_fd_sc_hs__nand2_1_19/B sky130_fd_sc_hs__dfxtp_4_5/a_696_458# sky130_fd_sc_hs__nor2b_1_1/Y
+ sky130_fd_sc_hs__nor2b_1_5/a_278_368# sky130_fd_sc_hs__dfxtp_4_17/a_1178_124# sky130_fd_sc_hs__a22o_1_39/X
+ m3_13600_5433# sky130_fd_sc_hs__dfxtp_4_63/a_437_503# sky130_fd_sc_hs__nand2_2_5/B
+ sky130_fd_sc_hs__dfxtp_4_23/a_735_102# sky130_fd_sc_hs__xnor2_1_53/A sky130_fd_sc_hs__dfxtp_4_61/a_735_102#
+ sky130_fd_sc_hs__dfxtp_4_57/a_1034_424# sky130_fd_sc_hs__xnor2_1_63/B sky130_fd_sc_hs__dfxtp_4_37/a_1141_508#
+ sky130_fd_sc_hs__nand2_1_47/B sky130_fd_sc_hs__a22o_1_29/X sky130_fd_sc_hs__xnor2_1_65/Y
+ m3_13600_4701# sky130_fd_sc_hs__dfxtp_4_1/a_437_503# sky130_fd_sc_hs__dfxtp_4_67/a_1178_124#
+ sky130_fd_sc_hs__dfxtp_4_9/a_735_102# sky130_fd_sc_hs__a22o_1_13/a_132_392# sky130_fd_sc_hs__dfxtp_4_15/a_1178_124#
+ sky130_fd_sc_hs__xnor2_1_15/A sky130_fd_sc_hs__nand2_1_1/B sky130_fd_sc_hs__xnor2_1_43/B
+ sky130_fd_sc_hs__dfxtp_4_35/a_651_503# sky130_fd_sc_hs__dfxtp_4_8/D sky130_fd_sc_hs__xnor2_1_29/A
+ sky130_fd_sc_hs__nand2_1_7/B sky130_fd_sc_hs__dfxtp_4_13/a_735_102# sky130_fd_sc_hs__dfxtp_4_47/a_696_458#
+ sky130_fd_sc_hs__nand2_1_31/B sky130_fd_sc_hs__dfxtp_4_51/a_735_102# sky130_fd_sc_hs__a22o_1_59/X
+ sky130_fd_sc_hs__dfxtp_4_35/a_1141_508# sky130_fd_sc_hs__a22o_1_25/a_222_392# sky130_fd_sc_hs__sdlclkp_2_1/a_288_48#
+ sky130_fd_sc_hs__xnor2_1_55/B sky130_fd_sc_hs__xnor2_1_17/B sky130_fd_sc_hs__xnor2_1_43/A
+ sky130_fd_sc_hs__xnor2_1_7/A sky130_fd_sc_hs__dfxtp_4_65/a_1178_124# sky130_fd_sc_hs__xnor2_1_59/Y
+ sky130_fd_sc_hs__a22o_1_41/X sky130_fd_sc_hs__a22o_1_21/a_230_79# sky130_fd_sc_hs__nand2_1_57/a_117_74#
+ sky130_fd_sc_hs__a22o_1_1/a_222_392# sky130_fd_sc_hs__xnor2_1_19/B sky130_fd_sc_hs__xnor2_1_35/a_293_74#
+ sky130_fd_sc_hs__nand2_1_23/a_117_74# sky130_fd_sc_hs__dfxtp_4_73/a_206_368# sky130_fd_sc_hs__dfxtp_4_25/a_651_503#
+ sky130_fd_sc_hs__xnor2_1_1/a_138_385# sky130_fd_sc_hs__dfxtp_4_37/a_696_458# sky130_fd_sc_hs__dfxtp_4_67/a_544_485#
+ sky130_fd_sc_hs__dfxtp_4_43/a_27_74# sky130_fd_sc_hs__a22o_1_9/X sky130_fd_sc_hs__dfxtp_4_55/a_1034_424#
+ sky130_fd_sc_hs__xnor2_1_39/a_112_119# sky130_fd_sc_hs__a22o_1_15/a_222_392# sky130_fd_sc_hs__conb_1_1/HI
+ sky130_fd_sc_hs__nand2_1_23/B sky130_fd_sc_hs__nand2_1_53/B sky130_fd_sc_hs__dfxtp_4_9/a_1178_124#
+ sky130_fd_sc_hs__nor2b_1_4/A sky130_fd_sc_hs__dfxtp_4_47/a_1226_296# m3_13600_11045#
+ sky130_fd_sc_hs__a22o_1_17/X sky130_fd_sc_hs__xnor2_1_29/a_376_368# sky130_fd_sc_hs__dfxtp_4_5/a_544_485#
+ sky130_fd_sc_hs__a22o_1_3/X sky130_fd_sc_hs__a22o_1_31/a_132_392# sky130_fd_sc_hs__xnor2_1_61/A
+ sky130_fd_sc_hs__dfxtp_4_15/a_651_503# sky130_fd_sc_hs__dfxtp_4_73/a_437_503# sky130_fd_sc_hs__a22o_1_25/a_230_79#
+ sky130_fd_sc_hs__dfxtp_4_27/a_696_458# sky130_fd_sc_hs__dfxtp_4_65/a_696_458# sky130_fd_sc_hs__dfxtp_4_33/a_735_102#
+ sky130_fd_sc_hs__dfxtp_4_71/a_735_102# m3_13600_7263# sky130_fd_sc_hs__a22o_1_43/a_222_392#
+ sky130_fd_sc_hs__xnor2_1_50/Y sky130_fd_sc_hs__dfxtp_4_8/a_1178_124# sky130_fd_sc_hs__xnor2_1_53/B
+ sky130_fd_sc_hs__xnor2_1_19/a_376_368# sky130_fd_sc_hs__dfxtp_4_63/a_1178_124# sky130_fd_sc_hs__dfxtp_4_4/a_696_458#
+ sky130_fd_sc_hs__nor2b_1_4/a_278_368# sky130_fd_sc_hs__dfxtp_4_13/a_1178_124# sky130_fd_sc_hs__a22o_1_61/a_132_392#
+ sky130_fd_sc_hs__dfxtp_4_53/a_206_368# sky130_fd_sc_hs__a22o_1_21/a_52_123# sky130_fd_sc_hs__dfxtp_4_45/a_651_503#
+ sky130_fd_sc_hs__dfxtp_4_17/a_696_458# sky130_fd_sc_hs__dfxtp_4_47/a_544_485# sky130_fd_sc_hs__dfxtp_4_55/a_696_458#
+ sky130_fd_sc_hs__dfxtp_4_21/a_735_102# sky130_fd_sc_hs__dfxtp_4_37/a_27_74# sky130_fd_sc_hs__xnor2_1_61/B
+ sky130_fd_sc_hs__a22o_1_61/X sky130_fd_sc_hs__xnor2_1_59/a_112_119# sky130_fd_sc_hs__xnor2_1_31/A
+ sky130_fd_sc_hs__a22o_1_33/a_222_392# sky130_fd_sc_hs__a22o_1_29/a_230_79# sky130_fd_sc_hs__dfxtp_4_45/a_1226_296#
+ sky130_fd_sc_hs__a22o_1_9/a_132_392# sky130_fd_sc_hs__xnor2_1_5/A sky130_fd_sc_hs__xnor2_1_57/Y
+ sky130_fd_sc_hs__a22o_1_31/X sky130_fd_sc_hs__dfxtp_4_51/a_27_74# sky130_fd_sc_hs__nor2b_1_8/a_27_112#
+ sky130_fd_sc_hs__xnor2_1_47/a_376_368# sky130_fd_sc_hs__xnor2_1_53/a_293_74# sky130_fd_sc_hs__nand2_1_43/a_117_74#
+ sky130_fd_sc_hs__dfxtp_4_8/a_735_102# sky130_fd_sc_hs__xnor2_1_21/a_293_74# sky130_fd_sc_hs__xnor2_1_39/a_138_385#
+ sky130_fd_sc_hs__xnor2_1_63/Y sky130_fd_sc_hs__a22o_1_51/a_132_392# sky130_fd_sc_hs__dfxtp_4_43/a_206_368#
+ sky130_fd_sc_hs__dfxtp_4_53/a_437_503# sky130_fd_sc_hs__dfxtp_4_37/a_544_485# sky130_fd_sc_hs__a22o_1_57/X
+ sky130_fd_sc_hs__dfxtp_4_53/a_1034_424# sky130_fd_sc_hs__a22o_1_25/a_52_123# sky130_fd_sc_hs__dfxtp_4_33/a_1141_508#
+ sky130_fd_sc_hs__dfxtp_4_63/Q sky130_fd_sc_hs__a22o_1_23/a_222_392# sky130_fd_sc_hs__a22o_1_63/a_222_392#
+ sky130_fd_sc_hs__dfxtp_4_7/a_1178_124# sky130_fd_sc_hs__a22o_1_53/X sky130_fd_sc_hs__nand2_2_5/Y
+ sky130_fd_sc_hs__dfxtp_4_61/a_1178_124# sky130_fd_sc_hs__a22o_1_1/a_230_79# sky130_fd_sc_hs__a22o_1_43/a_230_79#
+ sky130_fd_sc_hs__a22o_1_11/a_230_79# sky130_fd_sc_hs__a22o_1_41/a_132_392# sky130_fd_sc_hs__nand2_1_13/a_117_74#
+ sky130_fd_sc_hs__dfxtp_4_43/a_437_503# sky130_fd_sc_hs__dfxtp_4_27/a_544_485# sky130_fd_sc_hs__dfxtp_4_63/a_651_503#
+ sky130_fd_sc_hs__nand2_1_7/a_117_74# sky130_fd_sc_hs__dfxtp_4_35/a_696_458# sky130_fd_sc_hs__dfxtp_4_65/a_544_485#
+ sky130_fd_sc_hs__dfxtp_4_51/a_1034_424# sky130_fd_sc_hs__dfxtp_4_41/a_735_102# sky130_fd_sc_hs__dfxtp_4_32/a_1141_508#
+ sky130_fd_sc_hs__dfxtp_4_49/a_1141_508# sky130_fd_sc_hs__nand2_1_55/B sky130_fd_sc_hs__a22o_1_53/a_222_392#
+ sky130_fd_sc_hs__sdlclkp_2_1/a_114_112# sky130_fd_sc_hs__xnor2_1_9/a_293_74# sky130_fd_sc_hs__dfxtp_4_43/a_1226_296#
+ sky130_fd_sc_hs__a22o_1_29/a_52_123# sky130_fd_sc_hs__nand2_1_37/B sky130_fd_sc_hs__dfxtp_4_1/a_651_503#
+ sky130_fd_sc_hs__xnor2_1_27/a_376_368# sky130_fd_sc_hs__dfxtp_4_4/a_544_485# sky130_fd_sc_hs__xnor2_1_67/a_376_368#
+ sky130_fd_sc_hs__a22o_1_27/X sky130_fd_sc_hs__a22o_1_1/X sky130_fd_sc_hs__xnor2_1_59/a_138_385#
+ sky130_fd_sc_hs__dfxtp_4_29/a_1178_124# m3_13600_2871# sky130_fd_sc_hs__a22o_1_5/a_230_79#
+ sky130_fd_sc_hs__dfxtp_4_23/a_206_368# sky130_fd_sc_hs__dfxtp_4_61/a_206_368# sky130_fd_sc_hs__dfxtp_4_17/a_544_485#
+ sky130_fd_sc_hs__a22o_1_15/a_230_79# sky130_fd_sc_hs__dfxtp_4_25/a_696_458# sky130_fd_sc_hs__dfxtp_4_55/a_544_485#
+ sky130_fd_sc_hs__dfxtp_4_32/a_735_102# sky130_fd_sc_hs__xnor2_1_29/a_293_74# sky130_fd_sc_hs__nand2_1_17/a_117_74#
+ sky130_fd_sc_hs__dfxtp_4_69/a_1034_424# sky130_fd_sc_hs__xnor2_1_29/a_112_119# sky130_fd_sc_hs__a22o_1_37/X
+ sky130_fd_sc_hs__xnor2_1_31/B sky130_fd_sc_hs__dfxtp_4_19/a_1034_424# sky130_fd_sc_hs__xnor2_1_33/A
+ sky130_fd_sc_hs__dfxtp_4_9/a_206_368# sky130_fd_sc_hs__xnor2_1_57/a_376_368# sky130_fd_sc_hs__sdlclkp_2_1/a_706_317#
+ sky130_fd_sc_hs__xnor2_1_11/B sky130_fd_sc_hs__a22o_1_1/a_52_123# sky130_fd_sc_hs__xnor2_1_39/B
+ sky130_fd_sc_hs__a22o_1_21/a_132_392# sky130_fd_sc_hs__dfxtp_4_13/a_206_368# sky130_fd_sc_hs__a22o_1_43/a_52_123#
+ sky130_fd_sc_hs__dfxtp_4_51/a_206_368# sky130_fd_sc_hs__a22o_1_47/X sky130_fd_sc_hs__dfxtp_4_23/a_437_503#
+ sky130_fd_sc_hs__a22o_1_11/a_52_123# sky130_fd_sc_hs__dfxtp_4_61/a_437_503# sky130_fd_sc_hs__nor2b_1_7/Y
+ sky130_fd_sc_hs__xnor2_1_51/A sky130_fd_sc_hs__dfxtp_4_15/a_696_458# sky130_fd_sc_hs__nor2b_1_5/Y
+ sky130_fd_sc_hs__a22o_1_9/a_230_79# sky130_fd_sc_hs__a22o_1_25/X sky130_fd_sc_hs__xnor2_1_19/a_112_119#
+ sky130_fd_sc_hs__nand2_1_45/B sky130_fd_sc_hs__dfxtp_4_5/a_1178_124# sky130_fd_sc_hs__a22o_1_19/a_230_79#
+ sky130_fd_sc_hs__dfxtp_4_41/a_1226_296# sky130_fd_sc_hs__dfxtp_4_59/a_1226_296#
+ sky130_fd_sc_hs__a22o_1_63/a_230_79# sky130_fd_sc_hs__dfxtp_4_51/Q sky130_fd_sc_hs__a22o_1_7/a_132_392#
+ sky130_fd_sc_hs__dfxtp_4_9/a_437_503# sky130_fd_sc_hs__xnor2_1_46/a_376_368# sky130_fd_sc_hs__nand2_1_33/a_117_74#
+ sky130_fd_sc_hs__xnor2_1_11/a_293_74# sky130_fd_sc_hs__dfxtp_4_27/a_1178_124# sky130_fd_sc_hs__a22o_1_11/a_132_392#
+ sky130_fd_sc_hs__dfxtp_4_13/a_437_503# sky130_fd_sc_hs__dfxtp_4_51/a_437_503# sky130_fd_sc_hs__a22o_1_5/a_52_123#
+ sky130_fd_sc_hs__dfxtp_4_35/a_544_485# sky130_fd_sc_hs__dfxtp_4_73/a_651_503# sky130_fd_sc_hs__dfxtp_4_45/a_696_458#
+ sky130_fd_sc_hs__a22o_1_15/a_52_123# sky130_fd_sc_hs__dfxtp_4_47/a_1141_508# sky130_fd_sc_hs__xnor2_1_47/a_112_119#
+ sky130_fd_sc_hs__dfxtp_4_4/a_1178_124# sky130_fd_sc_hs__dfxtp_4_17/a_1034_424# sky130_fd_sc_hs__xnor2_1_23/B
+ sky130_fd_sc_hs__xnor2_1_37/a_376_368# sky130_fd_sc_hs__xnor2_1_15/B sky130_fd_sc_hs__xnor2_1_7/Y
+ sky130_fd_sc_hs__xnor2_1_29/a_138_385# sky130_fd_sc_hs__a22o_1_33/a_230_79# sky130_fd_sc_hs__dfxtp_4_25/a_1178_124#
+ sky130_fd_sc_hs__xnor2_1_47/a_293_74# sky130_fd_sc_hs__nand2_1_37/a_117_74# sky130_fd_sc_hs__dfxtp_4_33/a_206_368#
+ sky130_fd_sc_hs__xnor2_1_15/a_293_74# sky130_fd_sc_hs__dfxtp_4_71/a_206_368# sky130_fd_sc_hs__dfxtp_4_25/a_544_485#
+ sky130_fd_sc_hs__dfxtp_4_67/a_1034_424# sky130_fd_sc_hs__a22o_1_13/a_222_392# sky130_fd_sc_hs__a22o_1_9/a_52_123#
+ sky130_fd_sc_hs__dfxtp_4_15/a_1034_424# sky130_fd_sc_hs__dfxtp_4_57/a_1226_296#
+ sky130_fd_sc_hs__a22o_1_19/a_52_123# sky130_fd_sc_hs__a22o_1_23/X sky130_fd_sc_hs__a22o_1_63/a_52_123#
+ sky130_fd_sc_hs__xnor2_1_19/a_138_385# sky130_fd_sc_hs__xnor2_1_9/a_376_368# sky130_fd_sc_hs__dfxtp_4_21/a_206_368#
+ sky130_fd_sc_hs__dfxtp_4_33/a_437_503# sky130_fd_sc_hs__dfxtp_4_71/a_437_503# sky130_fd_sc_hs__dfxtp_4_53/a_651_503#
+ sky130_fd_sc_hs__dfxtp_4_15/a_544_485# sky130_fd_sc_hs__dfxtp_4_63/a_696_458# sky130_fd_sc_hs__dfxtp_4_65/a_1034_424#
+ sky130_fd_sc_hs__xnor2_1_19/a_293_74# sky130_fd_sc_hs__dfxtp_4_45/a_1141_508# sky130_fd_sc_hs__xnor2_1_27/a_112_119#
+ sky130_fd_sc_hs__xnor2_1_67/a_112_119# sky130_fd_sc_hs__dfxtp_4_1/a_1178_124# sky130_fd_sc_hs__conb_1_1/a_21_290#
+ sky130_fd_sc_hs__xnor2_1_63/a_293_74# sky130_fd_sc_hs__dfxtp_4_8/a_206_368# sky130_fd_sc_hs__xnor2_1_17/a_376_368#
+ sky130_fd_sc_hs__dfxtp_4_63/a_27_74# sky130_fd_sc_hs__xnor2_1_21/A sky130_fd_sc_hs__xnor2_1_55/a_376_368#
+ sky130_fd_sc_hs__dfxtp_4_1/a_696_458# sky130_fd_sc_hs__nor2b_1_1/a_278_368# sky130_fd_sc_hs__xnor2_1_47/a_138_385#
+ sky130_fd_sc_hs__a22o_1_33/a_52_123# sky130_fd_sc_hs__dfxtp_4_9/a_1034_424# sky130_fd_sc_hs__dfxtp_4_21/a_437_503#
+ sky130_fd_sc_hs__dfxtp_4_1/a_27_74# sky130_fd_sc_hs__dfxtp_4_43/a_651_503# sky130_fd_sc_hs__dfxtp_4_1/Q
+ sky130_fd_sc_hs__dfxtp_4_45/a_544_485# sky130_fd_sc_hs__dfxtp_4_69/a_735_102# sky130_fd_sc_hs__xnor2_1_57/a_112_119#
+ sky130_fd_sc_hs__a22o_1_31/a_222_392# sky130_fd_sc_hs__xnor2_1_13/A sky130_fd_sc_hs__dfxtp_4_55/a_1226_296#
+ sky130_fd_sc_hs__nand2_2_5/a_27_74# sky130_fd_sc_hs__a22o_1_53/a_230_79# sky130_fd_sc_hs__dfxtp_4_8/a_437_503#
+ sky130_fd_sc_hs__xnor2_1_67/a_293_74# sky130_fd_sc_hs__xnor2_1_33/a_293_74# sky130_fd_sc_hs__dfxtp_4_7/a_735_102#
+ sky130_fd_sc_hs__dfxtp_4_23/a_1178_124# sky130_fd_sc_hs__dfxtp_4_41/a_206_368# sky130_fd_sc_hs__dfxtp_4_8/a_1034_424#
+ sky130_fd_sc_hs__dfxtp_4_63/a_1034_424# sky130_fd_sc_hs__dfxtp_4_59/a_735_102# sky130_fd_sc_hs__nand2_1_5/B
+ sky130_fd_sc_hs__dfxtp_4_43/a_1141_508# sky130_fd_sc_hs__xnor2_1_46/a_112_119# sky130_fd_sc_hs__a22o_1_61/a_222_392#
+ sky130_fd_sc_hs__dfxtp_4_13/a_1034_424# sky130_fd_sc_hs__dfxtp_4_73/a_1178_124#
+ sky130_fd_sc_hs__nand2_1_27/B sky130_fd_sc_hs__xnor2_1_13/B sky130_fd_sc_hs__dfxtp_4_57/a_27_74#
+ sky130_fd_sc_hs__a22o_1_57/a_230_79# sky130_fd_sc_hs__dfxtp_4_21/a_1178_124# sky130_fd_sc_hs__nor2b_1_1/a_27_112#
+ sky130_fd_sc_hs__xnor2_1_27/a_138_385# sky130_fd_sc_hs__a22o_1_23/a_230_79# sky130_fd_sc_hs__xnor2_1_67/a_138_385#
+ sky130_fd_sc_hs__nand2_1_41/B sky130_fd_sc_hs__a22o_1_9/a_222_392# sky130_fd_sc_hs__nand2_1_27/a_117_74#
+ sky130_fd_sc_hs__dfxtp_4_32/a_206_368# sky130_fd_sc_hs__dfxtp_4_23/a_651_503# sky130_fd_sc_hs__dfxtp_4_41/a_437_503#
+ sky130_fd_sc_hs__dfxtp_4_73/a_27_74# sky130_fd_sc_hs__dfxtp_4_61/a_651_503# sky130_fd_sc_hs__dfxtp_4_63/a_544_485#
+ sky130_fd_sc_hs__dfxtp_4_49/a_735_102# sky130_fd_sc_hs__dfxtp_4_73/a_696_458# sky130_fd_sc_hs__xnor2_1_37/a_112_119#
+ sky130_fd_sc_hs__a22o_1_51/a_222_392# sky130_fd_sc_hs__a22o_1_43/X sky130_fd_sc_hs__nand2_2_1/B
+ sky130_fd_sc_hs__dfxtp_4_9/a_651_503# sky130_fd_sc_hs__a22o_1_53/a_52_123# sky130_fd_sc_hs__a22o_1_49/X
+ sky130_fd_sc_hs__xnor2_1_25/a_376_368# sky130_fd_sc_hs__dfxtp_4_1/a_544_485# sky130_fd_sc_hs__xnor2_1_65/a_376_368#
+ sky130_fd_sc_hs__xnor2_1_57/a_138_385# sky130_fd_sc_hs__dfxtp_4_27/a_27_74# sky130_fd_sc_hs__a22o_1_39/a_132_392#
+ sky130_fd_sc_hs__dfxtp_4_7/a_1034_424# sky130_fd_sc_hs__dfxtp_4_13/a_651_503# sky130_fd_sc_hs__dfxtp_4_32/a_437_503#
+ sky130_fd_sc_hs__a22o_1_27/a_230_79# m3_13600_12265# sky130_fd_sc_hs__dfxtp_4_51/a_651_503#
+ sky130_fd_sc_hs__xnor2_1_59/B sky130_fd_sc_hs__xnor2_1_47/A sky130_fd_sc_hs__dfxtp_4_61/a_1034_424#
+ sky130_fd_sc_hs__dfxtp_4_41/a_1141_508# sky130_fd_sc_hs__dfxtp_4_59/a_1141_508#
+ sky130_fd_sc_hs__a22o_1_41/a_222_392# sky130_fd_sc_hs__dfxtp_4_53/a_1226_296# sky130_fd_sc_hs__xnor2_1_3/A
+ sky130_fd_sc_hs__dfxtp_4_71/a_1178_124# sky130_fd_sc_hs__xnor2_1_9/a_112_119# sky130_fd_sc_hs__nand2_1_3/a_117_74#
+ m3_13600_8483# sky130_fd_sc_hs__dfxtp_4_39/a_1178_124# sky130_fd_sc_hs__a22o_1_57/a_52_123#
+ sky130_fd_sc_hs__xnor2_1_46/a_138_385# sky130_fd_sc_hs__a22o_1_23/a_52_123# sky130_fd_sc_hs__dfxtp_4_67/a_27_74#
+ sky130_fd_sc_hs__dfxtp_4_53/a_696_458# sky130_fd_sc_hs__xnor2_1_17/a_112_119# sky130_fd_sc_hs__xnor2_1_11/A
+ sky130_fd_sc_hs__xnor2_1_55/a_112_119# sky130_fd_sc_hs__xnor2_1_1/A sky130_fd_sc_hs__dfxtp_4_51/a_1226_296#
+ sky130_fd_sc_hs__dfxtp_4_29/a_1034_424# sky130_fd_sc_hs__xnor2_1_59/A sky130_fd_sc_hs__xnor2_1_23/A
+ sky130_fd_sc_hs__nand2_1_39/B sky130_fd_sc_hs__dfxtp_4_5/a_27_74# sky130_fd_sc_hs__xnor2_1_57/a_293_74#
+ sky130_fd_sc_hs__xnor2_1_37/a_138_385# sky130_fd_sc_hs__a22o_1_59/a_132_392# sky130_fd_sc_hs__dfxtp_4_33/a_651_503#
+ sky130_fd_sc_hs__dfxtp_4_71/a_651_503# sky130_fd_sc_hs__dfxtp_4_43/a_696_458# sky130_fd_sc_hs__dfxtp_4_73/a_544_485#
+ sky130_fd_sc_hs__a22o_1_27/a_52_123# sky130_fd_sc_hs__dfxtp_4_57/a_1141_508# sky130_fd_sc_hs__a22o_1_21/a_222_392#
+ sky130_fd_sc_hs__dfxtp_4_35/a_27_74# sky130_fd_sc_hs__dfxtp_4_69/a_1226_296# sky130_fd_sc_hs__xnor2_1_37/B
+ sky130_fd_sc_hs__dfxtp_4_19/a_1226_296# sky130_fd_sc_hs__xnor2_1_35/a_376_368# sky130_fd_sc_hs__a22o_1_47/a_230_79#
+ sky130_fd_sc_hs__dfxtp_4_37/a_1178_124# sky130_fd_sc_hs__dfxtp_4_5/a_1034_424# sky130_fd_sc_hs__a22o_1_49/a_132_392#
+ sky130_fd_sc_hs__a22o_1_7/a_222_392# sky130_fd_sc_hs__xnor2_1_27/a_293_74# sky130_fd_sc_hs__dfxtp_4_21/a_651_503#
+ sky130_fd_sc_hs__xnor2_1_9/a_138_385# sky130_fd_sc_hs__a22o_1_11/a_222_392# m3_13600_14095#
+ sky130_fd_sc_hs__xnor2_1_50/A sky130_fd_sc_hs__dfxtp_4_27/a_1034_424# sky130_fd_sc_hs__nand2_1_13/B
+ sky130_fd_sc_hs__dfxtp_4_8/a_651_503# m3_13600_9703# sky130_fd_sc_hs__dfxtp_4_35/a_1178_124#
+ sky130_fd_sc_hs__xnor2_1_17/a_138_385# sky130_fd_sc_hs__xnor2_1_55/a_138_385# sky130_fd_sc_hs__a22o_1_7/a_230_79#
+ sky130_fd_sc_hs__dfxtp_4_4/a_1034_424# sky130_fd_sc_hs__xnor2_1_7/a_376_368# sky130_fd_sc_hs__dfxtp_4_69/a_206_368#
+ sky130_fd_sc_hs__dfxtp_4_23/a_696_458# sky130_fd_sc_hs__dfxtp_4_53/a_544_485# sky130_fd_sc_hs__dfxtp_4_39/a_735_102#
+ sky130_fd_sc_hs__dfxtp_4_61/a_696_458# sky130_fd_sc_hs__dfxtp_4_55/a_1141_508# sky130_fd_sc_hs__xnor2_1_25/a_112_119#
+ sky130_fd_sc_hs__xnor2_1_65/a_112_119# sky130_fd_sc_hs__xnor2_1_43/a_293_74# sky130_fd_sc_hs__nand2_1_57/B
+ sky130_fd_sc_hs__dfxtp_4_25/a_1034_424# sky130_fd_sc_hs__dfxtp_4_7/a_206_368# sky130_fd_sc_hs__dfxtp_4_17/a_1226_296#
+ sky130_fd_sc_hs__xnor2_1_15/a_376_368# sky130_fd_sc_hs__xnor2_1_53/a_376_368# sky130_fd_sc_hs__dfxtp_4_9/a_696_458#
+ m3_13600_431# sky130_fd_sc_hs__dfxtp_4_45/a_27_74# sky130_fd_sc_hs__a22o_1_47/a_52_123#
+ sky130_fd_sc_hs__a22o_1_29/a_132_392# sky130_fd_sc_hs__dfxtp_4_59/a_206_368# sky130_fd_sc_hs__dfxtp_4_69/a_437_503#
+ sky130_fd_sc_hs__dfxtp_4_41/a_651_503# sky130_fd_sc_hs__dfxtp_4_43/a_544_485# sky130_fd_sc_hs__dfxtp_4_13/a_696_458#
+ sky130_fd_sc_hs__dfxtp_4_29/a_735_102# sky130_fd_sc_hs__dfxtp_4_51/a_696_458# sky130_fd_sc_hs__xnor2_1_61/Y
+ sky130_fd_sc_hs__dfxtp_4_67/a_1226_296# sky130_fd_sc_hs__a22o_1_5/a_132_392# sky130_fd_sc_hs__and2b_2_1/a_198_48#
+ sky130_fd_sc_hs__dfxtp_4_7/a_437_503# sky130_fd_sc_hs__dfxtp_4_15/a_1226_296# sky130_fd_sc_hs__dfxtp_4_69/a_27_74#
+ sky130_fd_sc_hs__xnor2_1_46/a_293_74# sky130_fd_sc_hs__dfxtp_4_1/a_1034_424# sky130_fd_sc_hs__a22o_1_19/a_132_392#
+ sky130_fd_sc_hs__dfxtp_4_49/a_206_368# sky130_fd_sc_hs__a22o_1_7/a_52_123# sky130_fd_sc_hs__dfxtp_4_59/a_437_503#
+ sky130_fd_sc_hs__dfxtp_4_32/a_651_503# sky130_fd_sc_hs__dfxtp_4_7/a_27_74# sky130_fd_sc_hs__nand2_2_1/a_27_74#
+ sky130_fd_sc_hs__dfxtp_4_19/a_735_102# sky130_fd_sc_hs__dfxtp_4_57/a_735_102# sky130_fd_sc_hs__dfxtp_4_65/a_1226_296#
+ sky130_fd_sc_hs__xnor2_1_37/A sky130_fd_sc_hs__xnor2_1_33/a_376_368# sky130_fd_sc_hs__a22o_1_37/a_230_79#
+ sky130_fd_sc_hs__xnor2_1_25/a_138_385# sky130_fd_sc_hs__dfxtp_4_39/a_27_74# sky130_fd_sc_hs__xnor2_1_65/a_138_385#
+ sky130_fd_sc_hs__nor2b_1_9/a_278_368# sky130_fd_sc_hs__dfxtp_4_49/a_437_503# sky130_fd_sc_hs__and2b_2_1/a_505_74#
+ sky130_fd_sc_hs__nand2_1_51/a_117_74# sky130_fd_sc_hs__dfxtp_4_23/a_544_485# sky130_fd_sc_hs__dfxtp_4_33/a_696_458#
+ sky130_fd_sc_hs__dfxtp_4_61/a_544_485# sky130_fd_sc_hs__dfxtp_4_9/a_1226_296# sky130_fd_sc_hs__dfxtp_4_53/a_1141_508#
+ sky130_fd_sc_hs__dfxtp_4_71/a_696_458# sky130_fd_sc_hs__xnor2_1_35/a_112_119# sky130_fd_sc_hs__dfxtp_4_23/a_1034_424#
+ sky130_fd_sc_hs__dfxtp_4_9/a_544_485# sky130_fd_sc_hs__xnor2_1_63/a_376_368# sky130_fd_sc_hs__dfxtp_4_33/a_1178_124#
+ sky130_fd_sc_hs__xnor2_1_5/a_376_368# sky130_fd_sc_hs__dfxtp_4_13/a_544_485# sky130_fd_sc_hs__dfxtp_4_73/a_1034_424#
+ sky130_fd_sc_hs__dfxtp_4_21/a_696_458# sky130_fd_sc_hs__dfxtp_4_51/a_544_485# sky130_fd_sc_hs__dfxtp_4_8/a_1226_296#
+ sky130_fd_sc_hs__dfxtp_4_51/a_1141_508# sky130_fd_sc_hs__nand2_1_55/a_117_74# sky130_fd_sc_hs__dfxtp_4_21/a_1034_424#
+ sky130_fd_sc_hs__dfxtp_4_63/a_1226_296# sky130_fd_sc_hs__dfxtp_4_23/a_27_74# sky130_fd_sc_hs__xnor2_1_7/a_112_119#
+ sky130_fd_sc_hs__dfxtp_4_13/a_1226_296# sky130_fd_sc_hs__dfxtp_4_8/a_696_458# sky130_fd_sc_hs__dfxtp_4_32/a_1178_124#
+ sky130_fd_sc_hs__dfxtp_4_49/a_1178_124# sky130_fd_sc_hs__a22o_1_37/a_52_123# sky130_fd_sc_hs__a22o_1_27/a_132_392#
+ sky130_fd_sc_hs__dfxtp_4_71/Q sky130_fd_sc_hs__dfxtp_4_67/a_735_102# sky130_fd_sc_hs__dfxtp_4_69/a_1141_508#
+ sky130_fd_sc_hs__xnor2_1_15/a_112_119# sky130_fd_sc_hs__xnor2_1_53/a_112_119# sky130_fd_sc_hs__a22o_1_39/a_222_392#
+ sky130_fd_sc_hs__a22o_1_55/a_230_79# sky130_fd_sc_hs__dfxtp_4_19/a_1141_508# sky130_fd_sc_hs__xnor2_1_37/a_293_74#
+ sky130_fd_sc_hs__xnor2_1_43/a_376_368# sky130_fd_sc_hs__dfxtp_4_5/a_735_102# sky130_fd_sc_hs__xnor2_1_35/a_138_385#
+ sky130_fd_sc_hs__sdlclkp_2_1/a_114_424# sky130_fd_sc_hs__a22o_1_57/a_132_392# sky130_fd_sc_hs__dfxtp_4_71/a_1034_424#
+ sky130_fd_sc_hs__dfxtp_4_7/a_1226_296# sky130_fd_sc_hs__dfxtp_4_33/a_544_485# sky130_fd_sc_hs__dfxtp_4_41/a_696_458#
+ sky130_fd_sc_hs__dfxtp_4_71/a_544_485# sky130_fd_sc_hs__xnor2_1_21/B sky130_fd_sc_hs__dfxtp_4_61/a_1226_296#
+ sky130_fd_sc_hs__dfxtp_4_39/a_1034_424# sky130_fd_sc_hs__dfxtp_4_17/a_27_74# sky130_fd_sc_hs__dfxtp_4_9/a_27_74#
+ sky130_fd_sc_hs__nor2b_1_5/a_27_112# sky130_fd_sc_hs__a22o_1_47/a_132_392# sky130_fd_sc_hs__nor2b_1_8/a_278_368#
+ sky130_fd_sc_hs__xnor2_1_9/B sky130_fd_sc_hs__dfxtp_4_39/a_206_368# sky130_fd_sc_hs__dfxtp_4_33/a_27_74#
+ sky130_fd_sc_hs__nand2_1_41/a_117_74# sky130_fd_sc_hs__dfxtp_4_69/a_651_503# sky130_fd_sc_hs__xnor2_1_51/a_293_74#
+ sky130_fd_sc_hs__dfxtp_4_21/a_544_485# sky130_fd_sc_hs__xnor2_1_7/a_138_385# sky130_fd_sc_hs__dfxtp_4_32/a_696_458#
+ sky130_fd_sc_hs__dfxtp_4_47/a_735_102# sky130_fd_sc_hs__xnor2_1_33/a_112_119# sky130_fd_sc_hs__a22o_1_59/a_222_392#
+ sky130_fd_sc_hs__dfxtp_4_17/a_1141_508# sky130_fd_sc_hs__a22o_1_55/a_52_123# sky130_fd_sc_hs__xnor2_1_3/a_293_74#
+ sky130_fd_sc_hs__dfxtp_4_7/a_651_503# sky130_fd_sc_hs__dfxtp_4_29/a_1226_296# sky130_fd_sc_hs__xnor2_1_23/a_376_368#
+ sky130_fd_sc_hs__dfxtp_4_8/a_544_485# sky130_fd_sc_hs__xnor2_1_47/B sky130_fd_sc_hs__dfxtp_4_47/a_1178_124#
+ sky130_fd_sc_hs__xnor2_1_15/a_138_385# sky130_fd_sc_hs__sdlclkp_2_1/a_1195_374#
+ sky130_fd_sc_hs__xnor2_1_53/a_138_385# sky130_fd_sc_hs__a22o_1_37/a_132_392# sky130_fd_sc_hs__dfxtp_4_29/a_206_368#
+ sky130_fd_sc_hs__dfxtp_4_39/a_437_503# sky130_fd_sc_hs__dfxtp_4_59/a_651_503# sky130_fd_sc_hs__dfxtp_4_37/a_735_102#
+ sky130_fd_sc_hs__dfxtp_4_67/a_1141_508# sky130_fd_sc_hs__and2b_2_1/a_27_74# sky130_fd_sc_hs__conb_1_1/a_165_290#
+ sky130_fd_sc_hs__xnor2_1_55/a_293_74# sky130_fd_sc_hs__nand2_1_45/a_117_74# sky130_fd_sc_hs__xnor2_1_63/a_112_119#
+ sky130_fd_sc_hs__a22o_1_49/a_222_392# sky130_fd_sc_hs__dfxtp_4_37/a_1034_424# sky130_fd_sc_hs__xnor2_1_23/a_293_74#
+ sky130_fd_sc_hs__dfxtp_4_15/a_1141_508# sky130_fd_sc_hs__nand2_1_5/a_117_74# m3_13600_13485#
+ sky130_fd_sc_hs__xnor2_1_5/a_112_119# sky130_fd_sc_hs__xnor2_1_13/a_376_368# sky130_fd_sc_hs__xnor2_1_51/a_376_368#
+ sky130_fd_sc_hs__xnor2_1_7/a_293_74# sky130_fd_sc_hs__dfxtp_4_19/a_206_368# sky130_fd_sc_hs__dfxtp_4_57/a_206_368#
+ sky130_fd_sc_hs__sdlclkp_2_1/a_318_74# sky130_fd_sc_hs__dfxtp_4_29/a_437_503# sky130_fd_sc_hs__dfxtp_4_49/a_651_503#
+ sky130_fd_sc_hs__dfxtp_4_25/a_27_74# sky130_fd_sc_hs__dfxtp_4_5/a_1226_296# sky130_fd_sc_hs__dfxtp_4_41/a_544_485#
+ sky130_fd_sc_hs__dfxtp_4_27/a_735_102# sky130_fd_sc_hs__dfxtp_4_65/a_1141_508# sky130_fd_sc_hs__dfxtp_4_65/a_735_102#
+ sky130_fd_sc_hs__a22o_1_3/a_230_79# sky130_fd_sc_hs__dfxtp_4_35/a_1034_424# sky130_fd_sc_hs__a22o_1_13/a_230_79#
+ sky130_fd_sc_hs__dfxtp_4_41/a_27_74# sky130_fd_sc_hs__a22o_1_3/a_132_392# sky130_fd_sc_hs__nand2_1_49/a_117_74#
+ sky130_fd_sc_hs__dfxtp_4_27/a_1226_296# sky130_fd_sc_hs__nand2_1_15/a_117_74# sky130_fd_sc_hs__xnor2_1_41/a_376_368#
+ sky130_fd_sc_hs__dfxtp_4_45/a_1178_124# sky130_fd_sc_hs__dfxtp_4_4/a_735_102# sky130_fd_sc_hs__nand2_1_9/a_117_74#
+ sky130_fd_sc_hs__xnor2_1_33/a_138_385# sky130_fd_sc_hs__a22o_1_17/a_132_392# sky130_fd_sc_hs__a22o_1_55/a_132_392#
+ sky130_fd_sc_hs__dfxtp_4_9/a_1141_508# sky130_fd_sc_hs__dfxtp_4_19/a_437_503# sky130_fd_sc_hs__dfxtp_4_57/a_437_503#
+ sky130_fd_sc_hs__dfxtp_4_4/a_1226_296# sky130_fd_sc_hs__dfxtp_4_32/a_544_485# sky130_fd_sc_hs__dfxtp_4_17/a_735_102#
+ sky130_fd_sc_hs__dfxtp_4_55/a_735_102# m3_13600_2261# sky130_fd_sc_hs__dfxtp_4_65/a_27_74#
+ sky130_fd_sc_hs__a22o_1_29/a_222_392# sky130_fd_sc_hs__xnor2_1_43/a_112_119# sky130_fd_sc_hs__a22o_1_19/X
+ sky130_fd_sc_hs__dfxtp_4_25/a_1226_296# sky130_fd_sc_hs__xnor2_1_31/a_376_368# sky130_fd_sc_hs__or2_1_1/a_63_368#
+ sky130_fd_sc_hs__a22o_1_17/a_230_79# sky130_fd_sc_hs__dfxtp_4_4/a_27_74# sky130_fd_sc_hs__a22o_1_61/a_230_79#
+ sky130_fd_sc_hs__xnor2_1_63/a_138_385# sky130_fd_sc_hs__a22o_1_5/a_222_392# sky130_fd_sc_hs__dfxtp_4_8/a_1141_508#
+ sky130_fd_sc_hs__xnor2_1_41/a_293_74# sky130_fd_sc_hs__nand2_1_31/a_117_74# sky130_fd_sc_hs__xnor2_1_5/a_138_385#
+ sky130_fd_sc_hs__dfxtp_4_63/a_1141_508# sky130_fd_sc_hs__a22o_1_19/a_222_392# sky130_fd_sc_hs__dfxtp_4_13/a_1141_508#
+ sky130_fd_sc_hs__a22o_1_3/a_52_123# sky130_fd_sc_hs__a22o_1_13/a_52_123# sky130_fd_sc_hs__dfxtp_4_43/a_1178_124#
+ sky130_fd_sc_hs__xnor2_1_61/a_376_368# sky130_fd_sc_hs__a22o_1_35/a_132_392# sky130_fd_sc_hs__dfxtp_4_67/a_206_368#
+ sky130_fd_sc_hs__dfxtp_4_1/a_1226_296# sky130_fd_sc_hs__dfxtp_4_69/a_696_458# sky130_fd_sc_hs__a22o_1_31/a_230_79#
+ sky130_fd_sc_hs__dfxtp_4_35/a_735_102# sky130_fd_sc_hs__xnor2_1_23/a_112_119# sky130_fd_sc_hs__nand2_1_35/a_117_74#
+ sky130_fd_sc_hs__dfxtp_4_59/a_27_74# sky130_fd_sc_hs__xnor2_1_13/a_293_74# sky130_fd_sc_hs__dfxtp_4_5/a_206_368#
+ sky130_fd_sc_hs__xnor2_1_50/a_376_368# sky130_fd_sc_hs__dfxtp_4_7/a_696_458# sky130_fd_sc_hs__nor2b_1_7/a_278_368#
+ sky130_fd_sc_hs__a22o_1_17/a_52_123# sky130_fd_sc_hs__xnor2_1_43/a_138_385# sky130_fd_sc_hs__dfxtp_4_7/a_1141_508#
+ sky130_fd_sc_hs__a22o_1_61/a_52_123# sky130_fd_sc_hs__dfxtp_4_67/a_437_503# sky130_fd_sc_hs__dfxtp_4_61/a_1141_508#
+ sky130_fd_sc_hs__dfxtp_4_25/a_735_102# sky130_fd_sc_hs__dfxtp_4_59/a_696_458# sky130_fd_sc_hs__xnor2_1_13/a_112_119#
+ sky130_fd_sc_hs__dfxtp_4_33/a_1034_424# sky130_fd_sc_hs__xnor2_1_51/a_112_119# sky130_fd_sc_hs__a22o_1_35/a_230_79#
+ m3_13600_4091# sky130_fd_sc_hs__dfxtp_4_23/a_1226_296# sky130_fd_sc_hs__nand2_1_39/a_117_74#
+ sky130_fd_sc_hs__dfxtp_4_29/a_27_74# sky130_fd_sc_hs__dfxtp_4_5/a_437_503# sky130_fd_sc_hs__xnor2_1_17/a_293_74#
+ sky130_fd_sc_hs__dfxtp_4_41/a_1178_124# sky130_fd_sc_hs__or2_1_1/a_152_368# sky130_fd_sc_hs__dfxtp_4_59/a_1178_124#
+ sky130_fd_sc_hs__xnor2_1_61/a_293_74# sky130_fd_sc_hs__dfxtp_4_47/a_206_368# sky130_fd_sc_hs__dfxtp_4_39/a_651_503#
+ sky130_fd_sc_hs__dfxtp_4_49/a_696_458# sky130_fd_sc_hs__dfxtp_4_15/a_735_102# sky130_fd_sc_hs__dfxtp_4_32/a_1034_424#
+ sky130_fd_sc_hs__dfxtp_4_73/a_1226_296# sky130_fd_sc_hs__a22o_1_27/a_222_392# sky130_fd_sc_hs__xnor2_1_41/a_112_119#
+ sky130_fd_sc_hs__a22o_1_31/a_52_123# sky130_fd_sc_hs__dfxtp_4_49/a_1034_424# sky130_fd_sc_hs__dfxtp_4_29/a_1141_508#
+ sky130_fd_sc_hs__dfxtp_4_21/a_1226_296# sky130_fd_sc_hs__a22o_1_39/a_230_79# sky130_fd_sc_hs__xnor2_1_23/a_138_385#
+ sky130_fd_sc_hs__a22o_1_51/a_230_79# sky130_fd_sc_hs__a22o_1_45/a_132_392# sky130_fd_sc_hs__dfxtp_4_37/a_206_368#
+ sky130_fd_sc_hs__xnor2_1_65/a_293_74# sky130_fd_sc_hs__nand2_1_53/a_117_74# sky130_fd_sc_hs__dfxtp_4_47/a_437_503#
+ sky130_fd_sc_hs__dfxtp_4_29/a_651_503# sky130_fd_sc_hs__xnor2_1_31/a_293_74# sky130_fd_sc_hs__nand2_1_21/a_117_74#
+ sky130_fd_sc_hs__dfxtp_4_69/a_544_485# sky130_fd_sc_hs__clkbuf_16_1/a_114_74# sky130_fd_sc_hs__dfxtp_4_45/a_735_102#
+ sky130_fd_sc_hs__dfxtp_4_13/a_27_74# sky130_fd_sc_hs__xnor2_1_31/a_112_119# sky130_fd_sc_hs__a22o_1_57/a_222_392#
+ sky130_fd_sc_hs__a22o_1_35/a_52_123# sky130_fd_sc_hs__xnor2_1_21/a_376_368# sky130_fd_sc_hs__dfxtp_4_7/a_544_485#
+ sky130_fd_sc_hs__dfxtp_4_57/a_1178_124# m3_13600_6043# sky130_fd_sc_hs__xnor2_1_13/a_138_385#
+ sky130_fd_sc_hs__xnor2_1_51/a_138_385# sky130_fd_sc_hs__dfxtp_4_5/a_1141_508# sky130_fd_sc_hs__xnor2_1_3/a_376_368#
+ sky130_fd_sc_hs__dfxtp_4_27/a_206_368# sky130_fd_sc_hs__dfxtp_4_65/a_206_368# sky130_fd_sc_hs__dfxtp_4_37/a_437_503#
+ sky130_fd_sc_hs__dfxtp_4_19/a_651_503# sky130_fd_sc_hs__dfxtp_4_57/a_651_503# sky130_fd_sc_hs__dfxtp_4_59/a_544_485#
+ sky130_fd_sc_hs__dfxtp_4_71/a_1226_296# sky130_fd_sc_hs__nand2_1_25/a_117_74# sky130_fd_sc_hs__xnor2_1_61/a_112_119#
+ sky130_fd_sc_hs__a22o_1_47/a_222_392# sky130_fd_sc_hs__dfxtp_4_27/a_1141_508# sky130_fd_sc_hs__dfxtp_4_53/a_27_74#
+ sky130_fd_sc_hs__dfxtp_4_4/a_206_368# sky130_fd_sc_hs__dfxtp_4_39/a_1226_296# sky130_fd_sc_hs__xnor2_1_11/a_376_368#
+ sky130_fd_sc_hs__a22o_1_39/a_52_123# sky130_fd_sc_hs__xnor2_1_41/a_138_385# sky130_fd_sc_hs__dfxtp_4_4/a_1141_508#
+ sky130_fd_sc_hs__a22o_1_25/a_132_392# sky130_fd_sc_hs__dfxtp_4_17/a_206_368# sky130_fd_sc_hs__xnor2_1_41/A
+ sky130_fd_sc_hs__dfxtp_4_55/a_206_368# sky130_fd_sc_hs__a22o_1_51/a_52_123# sky130_fd_sc_hs__dfxtp_4_27/a_437_503#
+ sky130_fd_sc_hs__dfxtp_4_65/a_437_503# sky130_fd_sc_hs__dfxtp_4_49/a_544_485# sky130_fd_sc_hs__dfxtp_4_63/a_735_102#
+ sky130_fd_sc_hs__dfxtp_4_47/a_1034_424# sky130_fd_sc_hs__xnor2_1_50/a_112_119# sky130_fd_sc_hs__a22o_1_37/a_222_392#
+ sky130_fd_sc_hs__a22o_1_59/a_230_79# sky130_fd_sc_hs__dfxtp_4_25/a_1141_508# sky130_fd_sc_hs__nor2b_1_4/a_27_112#
+ sky130_fd_sc_hs__sdlclkp_2_1/a_685_81# sky130_fd_sc_hs__a22o_1_1/a_132_392# sky130_fd_sc_hs__xnor2_1_39/a_293_74#
+ sky130_fd_sc_hs__nand2_1_29/a_117_74# sky130_fd_sc_hs__dfxtp_4_4/a_437_503# sky130_fd_sc_hs__dfxtp_4_55/a_1178_124#
+ sky130_fd_sc_hs__dfxtp_4_21/a_27_74# m3_13600_12875# sky130_fd_sc_hs__xnor2_1_50/a_293_74#
+ sky130_fd_sc_hs__dfxtp_4_1/a_735_102# sky130_fd_sc_hs__xnor2_1_31/a_138_385# sky130_fd_sc_hs__a22o_1_15/a_132_392#
+ sky130_fd_sc_hs__nand2_1_1/a_117_74# sky130_fd_sc_hs__dfxtp_4_17/a_437_503# sky130_fd_sc_hs__dfxtp_4_55/a_437_503#
+
Xsky130_fd_sc_hs__xnor2_1_7 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__xnor2_1_7/A sky130_fd_sc_hs__xnor2_1_7/Y
+ sky130_fd_sc_hs__xnor2_1_9/Y sky130_fd_sc_hs__xnor2_1_7/a_376_368# sky130_fd_sc_hs__xnor2_1_7/a_112_119#
+ sky130_fd_sc_hs__xnor2_1_7/a_138_385# sky130_fd_sc_hs__xnor2_1_7/a_293_74# sky130_fd_sc_hs__xnor2_1
Xsky130_fd_sc_hs__nor2b_1_10 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__dfxtp_4_71/Q sky130_fd_sc_hs__nor2b_1_8/Y
+ rst sky130_fd_sc_hs__nor2b_1_8/a_278_368# sky130_fd_sc_hs__nor2b_1_8/a_27_112# sky130_fd_sc_hs__nor2b_1
Xsky130_fd_sc_hs__a22o_1_14 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__a22o_1_15/X sky130_fd_sc_hs__nand2_1_29/B
+ sky130_fd_sc_hs__and2b_2_1/X init_val[7] rst sky130_fd_sc_hs__a22o_1_15/a_222_392#
+ sky130_fd_sc_hs__a22o_1_15/a_230_79# sky130_fd_sc_hs__a22o_1_15/a_52_123# sky130_fd_sc_hs__a22o_1_15/a_132_392#
+ sky130_fd_sc_hs__a22o_1
Xsky130_fd_sc_hs__a22o_1_25 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__a22o_1_25/X sky130_fd_sc_hs__nand2_1_9/B
+ sky130_fd_sc_hs__and2b_2_1/X init_val[5] rst sky130_fd_sc_hs__a22o_1_25/a_222_392#
+ sky130_fd_sc_hs__a22o_1_25/a_230_79# sky130_fd_sc_hs__a22o_1_25/a_52_123# sky130_fd_sc_hs__a22o_1_25/a_132_392#
+ sky130_fd_sc_hs__a22o_1
Xsky130_fd_sc_hs__a22o_1_58 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__a22o_1_59/X sky130_fd_sc_hs__nand2_2_3/B
+ sky130_fd_sc_hs__and2b_2_1/X init_val[26] rst sky130_fd_sc_hs__a22o_1_59/a_222_392#
+ sky130_fd_sc_hs__a22o_1_59/a_230_79# sky130_fd_sc_hs__a22o_1_59/a_52_123# sky130_fd_sc_hs__a22o_1_59/a_132_392#
+ sky130_fd_sc_hs__a22o_1
Xsky130_fd_sc_hs__a22o_1_47 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__a22o_1_47/X sky130_fd_sc_hs__nand2_1_49/B
+ sky130_fd_sc_hs__and2b_2_1/X init_val[29] rst sky130_fd_sc_hs__a22o_1_47/a_222_392#
+ sky130_fd_sc_hs__a22o_1_47/a_230_79# sky130_fd_sc_hs__a22o_1_47/a_52_123# sky130_fd_sc_hs__a22o_1_47/a_132_392#
+ sky130_fd_sc_hs__a22o_1
Xsky130_fd_sc_hs__a22o_1_36 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__a22o_1_37/X sky130_fd_sc_hs__xnor2_1_43/Y
+ sky130_fd_sc_hs__and2b_2_1/X init_val[0] rst sky130_fd_sc_hs__a22o_1_37/a_222_392#
+ sky130_fd_sc_hs__a22o_1_37/a_230_79# sky130_fd_sc_hs__a22o_1_37/a_52_123# sky130_fd_sc_hs__a22o_1_37/a_132_392#
+ sky130_fd_sc_hs__a22o_1
Xsky130_fd_sc_hs__nand2_1_14 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__dfxtp_4_1/Q sky130_fd_sc_hs__xnor2_1_15/A
+ eqn[13] sky130_fd_sc_hs__nand2_1_15/a_117_74# sky130_fd_sc_hs__nand2_1
Xsky130_fd_sc_hs__nand2_1_25 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_1_25/B sky130_fd_sc_hs__xnor2_1_31/A
+ eqn[14] sky130_fd_sc_hs__nand2_1_25/a_117_74# sky130_fd_sc_hs__nand2_1
Xsky130_fd_sc_hs__nand2_1_36 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_1_37/B sky130_fd_sc_hs__xnor2_1_37/B
+ eqn[24] sky130_fd_sc_hs__nand2_1_37/a_117_74# sky130_fd_sc_hs__nand2_1
Xsky130_fd_sc_hs__nand2_1_47 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_1_47/B sky130_fd_sc_hs__xnor2_1_55/B
+ eqn[19] sky130_fd_sc_hs__nand2_1_47/a_117_74# sky130_fd_sc_hs__nand2_1
Xsky130_fd_sc_hs__dfxtp_4_4 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_2_1/B sky130_fd_sc_hs__a22o_1_5/X
+ sky130_fd_sc_hs__dfxtp_4_9/CLK sky130_fd_sc_hs__dfxtp_4_4/a_1226_296# sky130_fd_sc_hs__dfxtp_4_4/a_735_102#
+ sky130_fd_sc_hs__dfxtp_4_4/a_1141_508# sky130_fd_sc_hs__dfxtp_4_4/a_206_368# sky130_fd_sc_hs__dfxtp_4_4/a_437_503#
+ sky130_fd_sc_hs__dfxtp_4_4/a_27_74# sky130_fd_sc_hs__dfxtp_4_4/a_651_503# sky130_fd_sc_hs__dfxtp_4_4/a_696_458#
+ sky130_fd_sc_hs__dfxtp_4_4/a_544_485# sky130_fd_sc_hs__dfxtp_4_4/a_1178_124# sky130_fd_sc_hs__dfxtp_4_4/a_1034_424#
+ sky130_fd_sc_hs__dfxtp_4
Xsky130_fd_sc_hs__xnor2_1_8 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__xnor2_1_9/A sky130_fd_sc_hs__xnor2_1_9/Y
+ sky130_fd_sc_hs__xnor2_1_9/B sky130_fd_sc_hs__xnor2_1_9/a_376_368# sky130_fd_sc_hs__xnor2_1_9/a_112_119#
+ sky130_fd_sc_hs__xnor2_1_9/a_138_385# sky130_fd_sc_hs__xnor2_1_9/a_293_74# sky130_fd_sc_hs__xnor2_1
Xsky130_fd_sc_hs__nor2b_1_11 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__dfxtp_4_63/Q sky130_fd_sc_hs__nor2b_1_9/Y
+ rst sky130_fd_sc_hs__nor2b_1_9/a_278_368# sky130_fd_sc_hs__nor2b_1_9/a_27_112# sky130_fd_sc_hs__nor2b_1
Xsky130_fd_sc_hs__a22o_1_15 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__a22o_1_15/X sky130_fd_sc_hs__nand2_1_29/B
+ sky130_fd_sc_hs__and2b_2_1/X init_val[7] rst sky130_fd_sc_hs__a22o_1_15/a_222_392#
+ sky130_fd_sc_hs__a22o_1_15/a_230_79# sky130_fd_sc_hs__a22o_1_15/a_52_123# sky130_fd_sc_hs__a22o_1_15/a_132_392#
+ sky130_fd_sc_hs__a22o_1
Xsky130_fd_sc_hs__a22o_1_26 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__a22o_1_27/X sky130_fd_sc_hs__nand2_1_17/B
+ sky130_fd_sc_hs__and2b_2_1/X init_val[4] rst sky130_fd_sc_hs__a22o_1_27/a_222_392#
+ sky130_fd_sc_hs__a22o_1_27/a_230_79# sky130_fd_sc_hs__a22o_1_27/a_52_123# sky130_fd_sc_hs__a22o_1_27/a_132_392#
+ sky130_fd_sc_hs__a22o_1
Xsky130_fd_sc_hs__a22o_1_59 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__a22o_1_59/X sky130_fd_sc_hs__nand2_2_3/B
+ sky130_fd_sc_hs__and2b_2_1/X init_val[26] rst sky130_fd_sc_hs__a22o_1_59/a_222_392#
+ sky130_fd_sc_hs__a22o_1_59/a_230_79# sky130_fd_sc_hs__a22o_1_59/a_52_123# sky130_fd_sc_hs__a22o_1_59/a_132_392#
+ sky130_fd_sc_hs__a22o_1
Xsky130_fd_sc_hs__a22o_1_48 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__a22o_1_49/X sky130_fd_sc_hs__nand2_1_27/B
+ sky130_fd_sc_hs__and2b_2_1/X init_val[22] rst sky130_fd_sc_hs__a22o_1_49/a_222_392#
+ sky130_fd_sc_hs__a22o_1_49/a_230_79# sky130_fd_sc_hs__a22o_1_49/a_52_123# sky130_fd_sc_hs__a22o_1_49/a_132_392#
+ sky130_fd_sc_hs__a22o_1
Xsky130_fd_sc_hs__a22o_1_37 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__a22o_1_37/X sky130_fd_sc_hs__xnor2_1_43/Y
+ sky130_fd_sc_hs__and2b_2_1/X init_val[0] rst sky130_fd_sc_hs__a22o_1_37/a_222_392#
+ sky130_fd_sc_hs__a22o_1_37/a_230_79# sky130_fd_sc_hs__a22o_1_37/a_52_123# sky130_fd_sc_hs__a22o_1_37/a_132_392#
+ sky130_fd_sc_hs__a22o_1
Xsky130_fd_sc_hs__nand2_1_15 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__dfxtp_4_1/Q sky130_fd_sc_hs__xnor2_1_15/A
+ eqn[13] sky130_fd_sc_hs__nand2_1_15/a_117_74# sky130_fd_sc_hs__nand2_1
Xsky130_fd_sc_hs__nand2_1_26 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_1_27/B sky130_fd_sc_hs__xnor2_1_19/B
+ eqn[21] sky130_fd_sc_hs__nand2_1_27/a_117_74# sky130_fd_sc_hs__nand2_1
Xsky130_fd_sc_hs__nand2_1_37 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_1_37/B sky130_fd_sc_hs__xnor2_1_37/B
+ eqn[24] sky130_fd_sc_hs__nand2_1_37/a_117_74# sky130_fd_sc_hs__nand2_1
Xsky130_fd_sc_hs__nand2_1_48 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_1_49/B sky130_fd_sc_hs__xnor2_1_59/A
+ eqn[28] sky130_fd_sc_hs__nand2_1_49/a_117_74# sky130_fd_sc_hs__nand2_1
Xsky130_fd_sc_hs__dfxtp_4_5 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_1_3/B sky130_fd_sc_hs__a22o_1_3/X
+ sky130_fd_sc_hs__dfxtp_4_9/CLK sky130_fd_sc_hs__dfxtp_4_5/a_1226_296# sky130_fd_sc_hs__dfxtp_4_5/a_735_102#
+ sky130_fd_sc_hs__dfxtp_4_5/a_1141_508# sky130_fd_sc_hs__dfxtp_4_5/a_206_368# sky130_fd_sc_hs__dfxtp_4_5/a_437_503#
+ sky130_fd_sc_hs__dfxtp_4_5/a_27_74# sky130_fd_sc_hs__dfxtp_4_5/a_651_503# sky130_fd_sc_hs__dfxtp_4_5/a_696_458#
+ sky130_fd_sc_hs__dfxtp_4_5/a_544_485# sky130_fd_sc_hs__dfxtp_4_5/a_1178_124# sky130_fd_sc_hs__dfxtp_4_5/a_1034_424#
+ sky130_fd_sc_hs__dfxtp_4
Xsky130_fd_sc_hs__xnor2_1_9 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__xnor2_1_9/A sky130_fd_sc_hs__xnor2_1_9/Y
+ sky130_fd_sc_hs__xnor2_1_9/B sky130_fd_sc_hs__xnor2_1_9/a_376_368# sky130_fd_sc_hs__xnor2_1_9/a_112_119#
+ sky130_fd_sc_hs__xnor2_1_9/a_138_385# sky130_fd_sc_hs__xnor2_1_9/a_293_74# sky130_fd_sc_hs__xnor2_1
Xsky130_fd_sc_hs__conb_1_0 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__conb_1_1/LO sky130_fd_sc_hs__conb_1_1/HI
+ sky130_fd_sc_hs__conb_1_1/a_165_290# sky130_fd_sc_hs__conb_1_1/a_21_290# sky130_fd_sc_hs__conb_1
Xsky130_fd_sc_hs__a22o_1_16 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__a22o_1_17/X sky130_fd_sc_hs__nand2_1_25/B
+ sky130_fd_sc_hs__and2b_2_1/X init_val[15] rst sky130_fd_sc_hs__a22o_1_17/a_222_392#
+ sky130_fd_sc_hs__a22o_1_17/a_230_79# sky130_fd_sc_hs__a22o_1_17/a_52_123# sky130_fd_sc_hs__a22o_1_17/a_132_392#
+ sky130_fd_sc_hs__a22o_1
Xsky130_fd_sc_hs__a22o_1_27 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__a22o_1_27/X sky130_fd_sc_hs__nand2_1_17/B
+ sky130_fd_sc_hs__and2b_2_1/X init_val[4] rst sky130_fd_sc_hs__a22o_1_27/a_222_392#
+ sky130_fd_sc_hs__a22o_1_27/a_230_79# sky130_fd_sc_hs__a22o_1_27/a_52_123# sky130_fd_sc_hs__a22o_1_27/a_132_392#
+ sky130_fd_sc_hs__a22o_1
Xsky130_fd_sc_hs__a22o_1_49 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__a22o_1_49/X sky130_fd_sc_hs__nand2_1_27/B
+ sky130_fd_sc_hs__and2b_2_1/X init_val[22] rst sky130_fd_sc_hs__a22o_1_49/a_222_392#
+ sky130_fd_sc_hs__a22o_1_49/a_230_79# sky130_fd_sc_hs__a22o_1_49/a_52_123# sky130_fd_sc_hs__a22o_1_49/a_132_392#
+ sky130_fd_sc_hs__a22o_1
Xsky130_fd_sc_hs__a22o_1_38 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__a22o_1_39/X sky130_fd_sc_hs__nand2_1_55/B
+ sky130_fd_sc_hs__and2b_2_1/X init_val[30] rst sky130_fd_sc_hs__a22o_1_39/a_222_392#
+ sky130_fd_sc_hs__a22o_1_39/a_230_79# sky130_fd_sc_hs__a22o_1_39/a_52_123# sky130_fd_sc_hs__a22o_1_39/a_132_392#
+ sky130_fd_sc_hs__a22o_1
Xsky130_fd_sc_hs__nand2_1_16 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_1_17/B sky130_fd_sc_hs__xnor2_1_11/B
+ eqn[3] sky130_fd_sc_hs__nand2_1_17/a_117_74# sky130_fd_sc_hs__nand2_1
Xsky130_fd_sc_hs__nand2_1_27 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_1_27/B sky130_fd_sc_hs__xnor2_1_19/B
+ eqn[21] sky130_fd_sc_hs__nand2_1_27/a_117_74# sky130_fd_sc_hs__nand2_1
Xsky130_fd_sc_hs__nand2_1_38 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_1_39/B sky130_fd_sc_hs__xnor2_1_35/A
+ eqn[26] sky130_fd_sc_hs__nand2_1_39/a_117_74# sky130_fd_sc_hs__nand2_1
Xsky130_fd_sc_hs__nand2_1_49 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_1_49/B sky130_fd_sc_hs__xnor2_1_59/A
+ eqn[28] sky130_fd_sc_hs__nand2_1_49/a_117_74# sky130_fd_sc_hs__nand2_1
Xsky130_fd_sc_hs__dfxtp_4_6 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__dfxtp_4_7/Q sky130_fd_sc_hs__a22o_1_7/X
+ sky130_fd_sc_hs__dfxtp_4_9/CLK sky130_fd_sc_hs__dfxtp_4_7/a_1226_296# sky130_fd_sc_hs__dfxtp_4_7/a_735_102#
+ sky130_fd_sc_hs__dfxtp_4_7/a_1141_508# sky130_fd_sc_hs__dfxtp_4_7/a_206_368# sky130_fd_sc_hs__dfxtp_4_7/a_437_503#
+ sky130_fd_sc_hs__dfxtp_4_7/a_27_74# sky130_fd_sc_hs__dfxtp_4_7/a_651_503# sky130_fd_sc_hs__dfxtp_4_7/a_696_458#
+ sky130_fd_sc_hs__dfxtp_4_7/a_544_485# sky130_fd_sc_hs__dfxtp_4_7/a_1178_124# sky130_fd_sc_hs__dfxtp_4_7/a_1034_424#
+ sky130_fd_sc_hs__dfxtp_4
Xsky130_fd_sc_hs__conb_1_1 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__conb_1_1/LO sky130_fd_sc_hs__conb_1_1/HI
+ sky130_fd_sc_hs__conb_1_1/a_165_290# sky130_fd_sc_hs__conb_1_1/a_21_290# sky130_fd_sc_hs__conb_1
Xsky130_fd_sc_hs__a22o_1_17 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__a22o_1_17/X sky130_fd_sc_hs__nand2_1_25/B
+ sky130_fd_sc_hs__and2b_2_1/X init_val[15] rst sky130_fd_sc_hs__a22o_1_17/a_222_392#
+ sky130_fd_sc_hs__a22o_1_17/a_230_79# sky130_fd_sc_hs__a22o_1_17/a_52_123# sky130_fd_sc_hs__a22o_1_17/a_132_392#
+ sky130_fd_sc_hs__a22o_1
Xsky130_fd_sc_hs__a22o_1_28 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__a22o_1_29/X sky130_fd_sc_hs__nand2_1_23/B
+ sky130_fd_sc_hs__and2b_2_1/X init_val[3] rst sky130_fd_sc_hs__a22o_1_29/a_222_392#
+ sky130_fd_sc_hs__a22o_1_29/a_230_79# sky130_fd_sc_hs__a22o_1_29/a_52_123# sky130_fd_sc_hs__a22o_1_29/a_132_392#
+ sky130_fd_sc_hs__a22o_1
Xsky130_fd_sc_hs__a22o_1_39 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__a22o_1_39/X sky130_fd_sc_hs__nand2_1_55/B
+ sky130_fd_sc_hs__and2b_2_1/X init_val[30] rst sky130_fd_sc_hs__a22o_1_39/a_222_392#
+ sky130_fd_sc_hs__a22o_1_39/a_230_79# sky130_fd_sc_hs__a22o_1_39/a_52_123# sky130_fd_sc_hs__a22o_1_39/a_132_392#
+ sky130_fd_sc_hs__a22o_1
Xsky130_fd_sc_hs__nand2_1_17 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_1_17/B sky130_fd_sc_hs__xnor2_1_11/B
+ eqn[3] sky130_fd_sc_hs__nand2_1_17/a_117_74# sky130_fd_sc_hs__nand2_1
Xsky130_fd_sc_hs__nand2_1_28 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_1_29/B sky130_fd_sc_hs__xnor2_1_19/A
+ eqn[6] sky130_fd_sc_hs__nand2_1_29/a_117_74# sky130_fd_sc_hs__nand2_1
Xsky130_fd_sc_hs__nand2_1_39 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_1_39/B sky130_fd_sc_hs__xnor2_1_35/A
+ eqn[26] sky130_fd_sc_hs__nand2_1_39/a_117_74# sky130_fd_sc_hs__nand2_1
Xsky130_fd_sc_hs__dfxtp_4_7 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__dfxtp_4_7/Q sky130_fd_sc_hs__a22o_1_7/X
+ sky130_fd_sc_hs__dfxtp_4_9/CLK sky130_fd_sc_hs__dfxtp_4_7/a_1226_296# sky130_fd_sc_hs__dfxtp_4_7/a_735_102#
+ sky130_fd_sc_hs__dfxtp_4_7/a_1141_508# sky130_fd_sc_hs__dfxtp_4_7/a_206_368# sky130_fd_sc_hs__dfxtp_4_7/a_437_503#
+ sky130_fd_sc_hs__dfxtp_4_7/a_27_74# sky130_fd_sc_hs__dfxtp_4_7/a_651_503# sky130_fd_sc_hs__dfxtp_4_7/a_696_458#
+ sky130_fd_sc_hs__dfxtp_4_7/a_544_485# sky130_fd_sc_hs__dfxtp_4_7/a_1178_124# sky130_fd_sc_hs__dfxtp_4_7/a_1034_424#
+ sky130_fd_sc_hs__dfxtp_4
Xsky130_fd_sc_hs__a22o_1_18 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__a22o_1_19/X sky130_fd_sc_hs__dfxtp_4_1/Q
+ sky130_fd_sc_hs__and2b_2_1/X init_val[14] rst sky130_fd_sc_hs__a22o_1_19/a_222_392#
+ sky130_fd_sc_hs__a22o_1_19/a_230_79# sky130_fd_sc_hs__a22o_1_19/a_52_123# sky130_fd_sc_hs__a22o_1_19/a_132_392#
+ sky130_fd_sc_hs__a22o_1
Xsky130_fd_sc_hs__a22o_1_29 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__a22o_1_29/X sky130_fd_sc_hs__nand2_1_23/B
+ sky130_fd_sc_hs__and2b_2_1/X init_val[3] rst sky130_fd_sc_hs__a22o_1_29/a_222_392#
+ sky130_fd_sc_hs__a22o_1_29/a_230_79# sky130_fd_sc_hs__a22o_1_29/a_52_123# sky130_fd_sc_hs__a22o_1_29/a_132_392#
+ sky130_fd_sc_hs__a22o_1
Xsky130_fd_sc_hs__nand2_1_18 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_1_19/B sky130_fd_sc_hs__xnor2_1_11/A
+ eqn[16] sky130_fd_sc_hs__nand2_1_19/a_117_74# sky130_fd_sc_hs__nand2_1
Xsky130_fd_sc_hs__nand2_1_29 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_1_29/B sky130_fd_sc_hs__xnor2_1_19/A
+ eqn[6] sky130_fd_sc_hs__nand2_1_29/a_117_74# sky130_fd_sc_hs__nand2_1
Xsky130_fd_sc_hs__dfxtp_4_8 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_1_1/B sky130_fd_sc_hs__dfxtp_4_8/D
+ sky130_fd_sc_hs__dfxtp_4_9/CLK sky130_fd_sc_hs__dfxtp_4_8/a_1226_296# sky130_fd_sc_hs__dfxtp_4_8/a_735_102#
+ sky130_fd_sc_hs__dfxtp_4_8/a_1141_508# sky130_fd_sc_hs__dfxtp_4_8/a_206_368# sky130_fd_sc_hs__dfxtp_4_8/a_437_503#
+ sky130_fd_sc_hs__dfxtp_4_8/a_27_74# sky130_fd_sc_hs__dfxtp_4_8/a_651_503# sky130_fd_sc_hs__dfxtp_4_8/a_696_458#
+ sky130_fd_sc_hs__dfxtp_4_8/a_544_485# sky130_fd_sc_hs__dfxtp_4_8/a_1178_124# sky130_fd_sc_hs__dfxtp_4_8/a_1034_424#
+ sky130_fd_sc_hs__dfxtp_4
Xsky130_fd_sc_hs__xnor2_1_60 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__xnor2_1_61/A sky130_fd_sc_hs__xnor2_1_61/Y
+ sky130_fd_sc_hs__xnor2_1_61/B sky130_fd_sc_hs__xnor2_1_61/a_376_368# sky130_fd_sc_hs__xnor2_1_61/a_112_119#
+ sky130_fd_sc_hs__xnor2_1_61/a_138_385# sky130_fd_sc_hs__xnor2_1_61/a_293_74# sky130_fd_sc_hs__xnor2_1
Xsky130_fd_sc_hs__a22o_1_19 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__a22o_1_19/X sky130_fd_sc_hs__dfxtp_4_1/Q
+ sky130_fd_sc_hs__and2b_2_1/X init_val[14] rst sky130_fd_sc_hs__a22o_1_19/a_222_392#
+ sky130_fd_sc_hs__a22o_1_19/a_230_79# sky130_fd_sc_hs__a22o_1_19/a_52_123# sky130_fd_sc_hs__a22o_1_19/a_132_392#
+ sky130_fd_sc_hs__a22o_1
Xsky130_fd_sc_hs__nand2_1_19 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_1_19/B sky130_fd_sc_hs__xnor2_1_11/A
+ eqn[16] sky130_fd_sc_hs__nand2_1_19/a_117_74# sky130_fd_sc_hs__nand2_1
Xsky130_fd_sc_hs__xnor2_1_50 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__xnor2_1_50/A sky130_fd_sc_hs__xnor2_1_50/Y
+ sky130_fd_sc_hs__xnor2_1_51/Y sky130_fd_sc_hs__xnor2_1_50/a_376_368# sky130_fd_sc_hs__xnor2_1_50/a_112_119#
+ sky130_fd_sc_hs__xnor2_1_50/a_138_385# sky130_fd_sc_hs__xnor2_1_50/a_293_74# sky130_fd_sc_hs__xnor2_1
Xsky130_fd_sc_hs__xnor2_1_61 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__xnor2_1_61/A sky130_fd_sc_hs__xnor2_1_61/Y
+ sky130_fd_sc_hs__xnor2_1_61/B sky130_fd_sc_hs__xnor2_1_61/a_376_368# sky130_fd_sc_hs__xnor2_1_61/a_112_119#
+ sky130_fd_sc_hs__xnor2_1_61/a_138_385# sky130_fd_sc_hs__xnor2_1_61/a_293_74# sky130_fd_sc_hs__xnor2_1
Xsky130_fd_sc_hs__dfxtp_4_9 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_1_7/B sky130_fd_sc_hs__a22o_1_9/X
+ sky130_fd_sc_hs__dfxtp_4_9/CLK sky130_fd_sc_hs__dfxtp_4_9/a_1226_296# sky130_fd_sc_hs__dfxtp_4_9/a_735_102#
+ sky130_fd_sc_hs__dfxtp_4_9/a_1141_508# sky130_fd_sc_hs__dfxtp_4_9/a_206_368# sky130_fd_sc_hs__dfxtp_4_9/a_437_503#
+ sky130_fd_sc_hs__dfxtp_4_9/a_27_74# sky130_fd_sc_hs__dfxtp_4_9/a_651_503# sky130_fd_sc_hs__dfxtp_4_9/a_696_458#
+ sky130_fd_sc_hs__dfxtp_4_9/a_544_485# sky130_fd_sc_hs__dfxtp_4_9/a_1178_124# sky130_fd_sc_hs__dfxtp_4_9/a_1034_424#
+ sky130_fd_sc_hs__dfxtp_4
Xsky130_fd_sc_hs__xnor2_1_40 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__xnor2_1_41/A sky130_fd_sc_hs__xnor2_1_41/Y
+ sky130_fd_sc_hs__xnor2_1_53/Y sky130_fd_sc_hs__xnor2_1_41/a_376_368# sky130_fd_sc_hs__xnor2_1_41/a_112_119#
+ sky130_fd_sc_hs__xnor2_1_41/a_138_385# sky130_fd_sc_hs__xnor2_1_41/a_293_74# sky130_fd_sc_hs__xnor2_1
Xsky130_fd_sc_hs__xnor2_1_51 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__xnor2_1_51/A sky130_fd_sc_hs__xnor2_1_51/Y
+ sky130_fd_sc_hs__xnor2_1_59/Y sky130_fd_sc_hs__xnor2_1_51/a_376_368# sky130_fd_sc_hs__xnor2_1_51/a_112_119#
+ sky130_fd_sc_hs__xnor2_1_51/a_138_385# sky130_fd_sc_hs__xnor2_1_51/a_293_74# sky130_fd_sc_hs__xnor2_1
Xsky130_fd_sc_hs__xnor2_1_62 DVSS DVDD DVDD DVSS inv_chicken[0] sky130_fd_sc_hs__xnor2_1_63/Y
+ sky130_fd_sc_hs__xnor2_1_63/B sky130_fd_sc_hs__xnor2_1_63/a_376_368# sky130_fd_sc_hs__xnor2_1_63/a_112_119#
+ sky130_fd_sc_hs__xnor2_1_63/a_138_385# sky130_fd_sc_hs__xnor2_1_63/a_293_74# sky130_fd_sc_hs__xnor2_1
Xsky130_fd_sc_hs__xnor2_1_30 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__xnor2_1_31/A sky130_fd_sc_hs__xnor2_1_33/A
+ sky130_fd_sc_hs__xnor2_1_31/B sky130_fd_sc_hs__xnor2_1_31/a_376_368# sky130_fd_sc_hs__xnor2_1_31/a_112_119#
+ sky130_fd_sc_hs__xnor2_1_31/a_138_385# sky130_fd_sc_hs__xnor2_1_31/a_293_74# sky130_fd_sc_hs__xnor2_1
Xsky130_fd_sc_hs__xnor2_1_41 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__xnor2_1_41/A sky130_fd_sc_hs__xnor2_1_41/Y
+ sky130_fd_sc_hs__xnor2_1_53/Y sky130_fd_sc_hs__xnor2_1_41/a_376_368# sky130_fd_sc_hs__xnor2_1_41/a_112_119#
+ sky130_fd_sc_hs__xnor2_1_41/a_138_385# sky130_fd_sc_hs__xnor2_1_41/a_293_74# sky130_fd_sc_hs__xnor2_1
Xsky130_fd_sc_hs__xnor2_1_52 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__xnor2_1_53/A sky130_fd_sc_hs__xnor2_1_53/Y
+ sky130_fd_sc_hs__xnor2_1_53/B sky130_fd_sc_hs__xnor2_1_53/a_376_368# sky130_fd_sc_hs__xnor2_1_53/a_112_119#
+ sky130_fd_sc_hs__xnor2_1_53/a_138_385# sky130_fd_sc_hs__xnor2_1_53/a_293_74# sky130_fd_sc_hs__xnor2_1
Xsky130_fd_sc_hs__xnor2_1_63 DVSS DVDD DVDD DVSS inv_chicken[0] sky130_fd_sc_hs__xnor2_1_63/Y
+ sky130_fd_sc_hs__xnor2_1_63/B sky130_fd_sc_hs__xnor2_1_63/a_376_368# sky130_fd_sc_hs__xnor2_1_63/a_112_119#
+ sky130_fd_sc_hs__xnor2_1_63/a_138_385# sky130_fd_sc_hs__xnor2_1_63/a_293_74# sky130_fd_sc_hs__xnor2_1
Xsky130_fd_sc_hs__xnor2_1_20 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__xnor2_1_21/A sky130_fd_sc_hs__xnor2_1_23/A
+ sky130_fd_sc_hs__xnor2_1_21/B sky130_fd_sc_hs__xnor2_1_21/a_376_368# sky130_fd_sc_hs__xnor2_1_21/a_112_119#
+ sky130_fd_sc_hs__xnor2_1_21/a_138_385# sky130_fd_sc_hs__xnor2_1_21/a_293_74# sky130_fd_sc_hs__xnor2_1
Xsky130_fd_sc_hs__xnor2_1_31 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__xnor2_1_31/A sky130_fd_sc_hs__xnor2_1_33/A
+ sky130_fd_sc_hs__xnor2_1_31/B sky130_fd_sc_hs__xnor2_1_31/a_376_368# sky130_fd_sc_hs__xnor2_1_31/a_112_119#
+ sky130_fd_sc_hs__xnor2_1_31/a_138_385# sky130_fd_sc_hs__xnor2_1_31/a_293_74# sky130_fd_sc_hs__xnor2_1
Xsky130_fd_sc_hs__xnor2_1_42 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__xnor2_1_43/A sky130_fd_sc_hs__xnor2_1_43/Y
+ sky130_fd_sc_hs__xnor2_1_43/B sky130_fd_sc_hs__xnor2_1_43/a_376_368# sky130_fd_sc_hs__xnor2_1_43/a_112_119#
+ sky130_fd_sc_hs__xnor2_1_43/a_138_385# sky130_fd_sc_hs__xnor2_1_43/a_293_74# sky130_fd_sc_hs__xnor2_1
Xsky130_fd_sc_hs__xnor2_1_53 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__xnor2_1_53/A sky130_fd_sc_hs__xnor2_1_53/Y
+ sky130_fd_sc_hs__xnor2_1_53/B sky130_fd_sc_hs__xnor2_1_53/a_376_368# sky130_fd_sc_hs__xnor2_1_53/a_112_119#
+ sky130_fd_sc_hs__xnor2_1_53/a_138_385# sky130_fd_sc_hs__xnor2_1_53/a_293_74# sky130_fd_sc_hs__xnor2_1
Xsky130_fd_sc_hs__xnor2_1_64 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nor2b_1_4/Y sky130_fd_sc_hs__xnor2_1_65/Y
+ sky130_fd_sc_hs__xnor2_1_67/Y sky130_fd_sc_hs__xnor2_1_65/a_376_368# sky130_fd_sc_hs__xnor2_1_65/a_112_119#
+ sky130_fd_sc_hs__xnor2_1_65/a_138_385# sky130_fd_sc_hs__xnor2_1_65/a_293_74# sky130_fd_sc_hs__xnor2_1
Xsky130_fd_sc_hs__xnor2_1_10 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__xnor2_1_11/A sky130_fd_sc_hs__xnor2_1_17/B
+ sky130_fd_sc_hs__xnor2_1_11/B sky130_fd_sc_hs__xnor2_1_11/a_376_368# sky130_fd_sc_hs__xnor2_1_11/a_112_119#
+ sky130_fd_sc_hs__xnor2_1_11/a_138_385# sky130_fd_sc_hs__xnor2_1_11/a_293_74# sky130_fd_sc_hs__xnor2_1
Xsky130_fd_sc_hs__xnor2_1_21 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__xnor2_1_21/A sky130_fd_sc_hs__xnor2_1_23/A
+ sky130_fd_sc_hs__xnor2_1_21/B sky130_fd_sc_hs__xnor2_1_21/a_376_368# sky130_fd_sc_hs__xnor2_1_21/a_112_119#
+ sky130_fd_sc_hs__xnor2_1_21/a_138_385# sky130_fd_sc_hs__xnor2_1_21/a_293_74# sky130_fd_sc_hs__xnor2_1
Xsky130_fd_sc_hs__xnor2_1_32 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__xnor2_1_33/A sky130_fd_sc_hs__xnor2_1_43/A
+ sky130_fd_sc_hs__xnor2_1_47/Y sky130_fd_sc_hs__xnor2_1_33/a_376_368# sky130_fd_sc_hs__xnor2_1_33/a_112_119#
+ sky130_fd_sc_hs__xnor2_1_33/a_138_385# sky130_fd_sc_hs__xnor2_1_33/a_293_74# sky130_fd_sc_hs__xnor2_1
Xsky130_fd_sc_hs__xnor2_1_43 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__xnor2_1_43/A sky130_fd_sc_hs__xnor2_1_43/Y
+ sky130_fd_sc_hs__xnor2_1_43/B sky130_fd_sc_hs__xnor2_1_43/a_376_368# sky130_fd_sc_hs__xnor2_1_43/a_112_119#
+ sky130_fd_sc_hs__xnor2_1_43/a_138_385# sky130_fd_sc_hs__xnor2_1_43/a_293_74# sky130_fd_sc_hs__xnor2_1
Xsky130_fd_sc_hs__xnor2_1_54 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__xnor2_1_55/A sky130_fd_sc_hs__xnor2_1_63/B
+ sky130_fd_sc_hs__xnor2_1_55/B sky130_fd_sc_hs__xnor2_1_55/a_376_368# sky130_fd_sc_hs__xnor2_1_55/a_112_119#
+ sky130_fd_sc_hs__xnor2_1_55/a_138_385# sky130_fd_sc_hs__xnor2_1_55/a_293_74# sky130_fd_sc_hs__xnor2_1
Xsky130_fd_sc_hs__xnor2_1_65 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nor2b_1_4/Y sky130_fd_sc_hs__xnor2_1_65/Y
+ sky130_fd_sc_hs__xnor2_1_67/Y sky130_fd_sc_hs__xnor2_1_65/a_376_368# sky130_fd_sc_hs__xnor2_1_65/a_112_119#
+ sky130_fd_sc_hs__xnor2_1_65/a_138_385# sky130_fd_sc_hs__xnor2_1_65/a_293_74# sky130_fd_sc_hs__xnor2_1
Xsky130_fd_sc_hs__xnor2_1_11 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__xnor2_1_11/A sky130_fd_sc_hs__xnor2_1_17/B
+ sky130_fd_sc_hs__xnor2_1_11/B sky130_fd_sc_hs__xnor2_1_11/a_376_368# sky130_fd_sc_hs__xnor2_1_11/a_112_119#
+ sky130_fd_sc_hs__xnor2_1_11/a_138_385# sky130_fd_sc_hs__xnor2_1_11/a_293_74# sky130_fd_sc_hs__xnor2_1
Xsky130_fd_sc_hs__xnor2_1_22 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__xnor2_1_23/A sky130_fd_sc_hs__xnor2_1_25/A
+ sky130_fd_sc_hs__xnor2_1_23/B sky130_fd_sc_hs__xnor2_1_23/a_376_368# sky130_fd_sc_hs__xnor2_1_23/a_112_119#
+ sky130_fd_sc_hs__xnor2_1_23/a_138_385# sky130_fd_sc_hs__xnor2_1_23/a_293_74# sky130_fd_sc_hs__xnor2_1
Xsky130_fd_sc_hs__xnor2_1_33 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__xnor2_1_33/A sky130_fd_sc_hs__xnor2_1_43/A
+ sky130_fd_sc_hs__xnor2_1_47/Y sky130_fd_sc_hs__xnor2_1_33/a_376_368# sky130_fd_sc_hs__xnor2_1_33/a_112_119#
+ sky130_fd_sc_hs__xnor2_1_33/a_138_385# sky130_fd_sc_hs__xnor2_1_33/a_293_74# sky130_fd_sc_hs__xnor2_1
Xsky130_fd_sc_hs__xnor2_1_44 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_2_5/Y sky130_fd_sc_hs__xnor2_1_47/B
+ sky130_fd_sc_hs__nand2_2_3/Y sky130_fd_sc_hs__xnor2_1_46/a_376_368# sky130_fd_sc_hs__xnor2_1_46/a_112_119#
+ sky130_fd_sc_hs__xnor2_1_46/a_138_385# sky130_fd_sc_hs__xnor2_1_46/a_293_74# sky130_fd_sc_hs__xnor2_1
Xsky130_fd_sc_hs__xnor2_1_55 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__xnor2_1_55/A sky130_fd_sc_hs__xnor2_1_63/B
+ sky130_fd_sc_hs__xnor2_1_55/B sky130_fd_sc_hs__xnor2_1_55/a_376_368# sky130_fd_sc_hs__xnor2_1_55/a_112_119#
+ sky130_fd_sc_hs__xnor2_1_55/a_138_385# sky130_fd_sc_hs__xnor2_1_55/a_293_74# sky130_fd_sc_hs__xnor2_1
Xsky130_fd_sc_hs__xnor2_1_66 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_2_5/B sky130_fd_sc_hs__xnor2_1_67/Y
+ inv_chicken[1] sky130_fd_sc_hs__xnor2_1_67/a_376_368# sky130_fd_sc_hs__xnor2_1_67/a_112_119#
+ sky130_fd_sc_hs__xnor2_1_67/a_138_385# sky130_fd_sc_hs__xnor2_1_67/a_293_74# sky130_fd_sc_hs__xnor2_1
Xsky130_fd_sc_hs__xnor2_1_12 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__xnor2_1_13/A sky130_fd_sc_hs__xnor2_1_25/B
+ sky130_fd_sc_hs__xnor2_1_13/B sky130_fd_sc_hs__xnor2_1_13/a_376_368# sky130_fd_sc_hs__xnor2_1_13/a_112_119#
+ sky130_fd_sc_hs__xnor2_1_13/a_138_385# sky130_fd_sc_hs__xnor2_1_13/a_293_74# sky130_fd_sc_hs__xnor2_1
Xsky130_fd_sc_hs__xnor2_1_23 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__xnor2_1_23/A sky130_fd_sc_hs__xnor2_1_25/A
+ sky130_fd_sc_hs__xnor2_1_23/B sky130_fd_sc_hs__xnor2_1_23/a_376_368# sky130_fd_sc_hs__xnor2_1_23/a_112_119#
+ sky130_fd_sc_hs__xnor2_1_23/a_138_385# sky130_fd_sc_hs__xnor2_1_23/a_293_74# sky130_fd_sc_hs__xnor2_1
Xsky130_fd_sc_hs__xnor2_1_34 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__xnor2_1_35/A sky130_fd_sc_hs__xnor2_1_47/A
+ sky130_fd_sc_hs__xnor2_1_35/B sky130_fd_sc_hs__xnor2_1_35/a_376_368# sky130_fd_sc_hs__xnor2_1_35/a_112_119#
+ sky130_fd_sc_hs__xnor2_1_35/a_138_385# sky130_fd_sc_hs__xnor2_1_35/a_293_74# sky130_fd_sc_hs__xnor2_1
Xsky130_fd_sc_hs__xnor2_1_45 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__xnor2_1_47/A sky130_fd_sc_hs__xnor2_1_47/Y
+ sky130_fd_sc_hs__xnor2_1_47/B sky130_fd_sc_hs__xnor2_1_47/a_376_368# sky130_fd_sc_hs__xnor2_1_47/a_112_119#
+ sky130_fd_sc_hs__xnor2_1_47/a_138_385# sky130_fd_sc_hs__xnor2_1_47/a_293_74# sky130_fd_sc_hs__xnor2_1
Xsky130_fd_sc_hs__xnor2_1_56 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__xnor2_1_61/Y sky130_fd_sc_hs__xnor2_1_57/Y
+ sky130_fd_sc_hs__xnor2_1_63/Y sky130_fd_sc_hs__xnor2_1_57/a_376_368# sky130_fd_sc_hs__xnor2_1_57/a_112_119#
+ sky130_fd_sc_hs__xnor2_1_57/a_138_385# sky130_fd_sc_hs__xnor2_1_57/a_293_74# sky130_fd_sc_hs__xnor2_1
Xsky130_fd_sc_hs__xnor2_1_67 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_2_5/B sky130_fd_sc_hs__xnor2_1_67/Y
+ inv_chicken[1] sky130_fd_sc_hs__xnor2_1_67/a_376_368# sky130_fd_sc_hs__xnor2_1_67/a_112_119#
+ sky130_fd_sc_hs__xnor2_1_67/a_138_385# sky130_fd_sc_hs__xnor2_1_67/a_293_74# sky130_fd_sc_hs__xnor2_1
Xsky130_fd_sc_hs__xnor2_1_13 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__xnor2_1_13/A sky130_fd_sc_hs__xnor2_1_25/B
+ sky130_fd_sc_hs__xnor2_1_13/B sky130_fd_sc_hs__xnor2_1_13/a_376_368# sky130_fd_sc_hs__xnor2_1_13/a_112_119#
+ sky130_fd_sc_hs__xnor2_1_13/a_138_385# sky130_fd_sc_hs__xnor2_1_13/a_293_74# sky130_fd_sc_hs__xnor2_1
Xsky130_fd_sc_hs__xnor2_1_24 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__xnor2_1_25/A sky130_fd_sc_hs__xnor2_1_39/B
+ sky130_fd_sc_hs__xnor2_1_25/B sky130_fd_sc_hs__xnor2_1_25/a_376_368# sky130_fd_sc_hs__xnor2_1_25/a_112_119#
+ sky130_fd_sc_hs__xnor2_1_25/a_138_385# sky130_fd_sc_hs__xnor2_1_25/a_293_74# sky130_fd_sc_hs__xnor2_1
Xsky130_fd_sc_hs__xnor2_1_35 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__xnor2_1_35/A sky130_fd_sc_hs__xnor2_1_47/A
+ sky130_fd_sc_hs__xnor2_1_35/B sky130_fd_sc_hs__xnor2_1_35/a_376_368# sky130_fd_sc_hs__xnor2_1_35/a_112_119#
+ sky130_fd_sc_hs__xnor2_1_35/a_138_385# sky130_fd_sc_hs__xnor2_1_35/a_293_74# sky130_fd_sc_hs__xnor2_1
Xsky130_fd_sc_hs__xnor2_1_46 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_2_5/Y sky130_fd_sc_hs__xnor2_1_47/B
+ sky130_fd_sc_hs__nand2_2_3/Y sky130_fd_sc_hs__xnor2_1_46/a_376_368# sky130_fd_sc_hs__xnor2_1_46/a_112_119#
+ sky130_fd_sc_hs__xnor2_1_46/a_138_385# sky130_fd_sc_hs__xnor2_1_46/a_293_74# sky130_fd_sc_hs__xnor2_1
Xsky130_fd_sc_hs__xnor2_1_57 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__xnor2_1_61/Y sky130_fd_sc_hs__xnor2_1_57/Y
+ sky130_fd_sc_hs__xnor2_1_63/Y sky130_fd_sc_hs__xnor2_1_57/a_376_368# sky130_fd_sc_hs__xnor2_1_57/a_112_119#
+ sky130_fd_sc_hs__xnor2_1_57/a_138_385# sky130_fd_sc_hs__xnor2_1_57/a_293_74# sky130_fd_sc_hs__xnor2_1
Xsky130_fd_sc_hs__xnor2_1_14 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__xnor2_1_15/A sky130_fd_sc_hs__xnor2_1_29/B
+ sky130_fd_sc_hs__xnor2_1_15/B sky130_fd_sc_hs__xnor2_1_15/a_376_368# sky130_fd_sc_hs__xnor2_1_15/a_112_119#
+ sky130_fd_sc_hs__xnor2_1_15/a_138_385# sky130_fd_sc_hs__xnor2_1_15/a_293_74# sky130_fd_sc_hs__xnor2_1
Xsky130_fd_sc_hs__xnor2_1_25 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__xnor2_1_25/A sky130_fd_sc_hs__xnor2_1_39/B
+ sky130_fd_sc_hs__xnor2_1_25/B sky130_fd_sc_hs__xnor2_1_25/a_376_368# sky130_fd_sc_hs__xnor2_1_25/a_112_119#
+ sky130_fd_sc_hs__xnor2_1_25/a_138_385# sky130_fd_sc_hs__xnor2_1_25/a_293_74# sky130_fd_sc_hs__xnor2_1
Xsky130_fd_sc_hs__xnor2_1_36 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__xnor2_1_37/A sky130_fd_sc_hs__xnor2_1_50/A
+ sky130_fd_sc_hs__xnor2_1_37/B sky130_fd_sc_hs__xnor2_1_37/a_376_368# sky130_fd_sc_hs__xnor2_1_37/a_112_119#
+ sky130_fd_sc_hs__xnor2_1_37/a_138_385# sky130_fd_sc_hs__xnor2_1_37/a_293_74# sky130_fd_sc_hs__xnor2_1
Xsky130_fd_sc_hs__xnor2_1_47 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__xnor2_1_47/A sky130_fd_sc_hs__xnor2_1_47/Y
+ sky130_fd_sc_hs__xnor2_1_47/B sky130_fd_sc_hs__xnor2_1_47/a_376_368# sky130_fd_sc_hs__xnor2_1_47/a_112_119#
+ sky130_fd_sc_hs__xnor2_1_47/a_138_385# sky130_fd_sc_hs__xnor2_1_47/a_293_74# sky130_fd_sc_hs__xnor2_1
Xsky130_fd_sc_hs__xnor2_1_58 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__xnor2_1_59/A sky130_fd_sc_hs__xnor2_1_59/Y
+ sky130_fd_sc_hs__xnor2_1_59/B sky130_fd_sc_hs__xnor2_1_59/a_376_368# sky130_fd_sc_hs__xnor2_1_59/a_112_119#
+ sky130_fd_sc_hs__xnor2_1_59/a_138_385# sky130_fd_sc_hs__xnor2_1_59/a_293_74# sky130_fd_sc_hs__xnor2_1
Xsky130_fd_sc_hs__sdlclkp_2_0 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__clkbuf_16_1/A clk
+ sky130_fd_sc_hs__or2_1_1/X sky130_fd_sc_hs__conb_1_1/LO sky130_fd_sc_hs__sdlclkp_2_1/a_114_112#
+ sky130_fd_sc_hs__sdlclkp_2_1/a_706_317# sky130_fd_sc_hs__sdlclkp_2_1/a_685_81# sky130_fd_sc_hs__sdlclkp_2_1/a_580_74#
+ sky130_fd_sc_hs__sdlclkp_2_1/a_288_48# sky130_fd_sc_hs__sdlclkp_2_1/a_114_424# sky130_fd_sc_hs__sdlclkp_2_1/a_1195_374#
+ sky130_fd_sc_hs__sdlclkp_2_1/a_708_451# sky130_fd_sc_hs__sdlclkp_2_1/a_1198_74#
+ sky130_fd_sc_hs__sdlclkp_2_1/a_318_74# sky130_fd_sc_hs__sdlclkp_2
Xsky130_fd_sc_hs__a22o_1_0 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__a22o_1_1/X sky130_fd_sc_hs__nand2_1_3/B
+ sky130_fd_sc_hs__and2b_2_1/X init_val[13] rst sky130_fd_sc_hs__a22o_1_1/a_222_392#
+ sky130_fd_sc_hs__a22o_1_1/a_230_79# sky130_fd_sc_hs__a22o_1_1/a_52_123# sky130_fd_sc_hs__a22o_1_1/a_132_392#
+ sky130_fd_sc_hs__a22o_1
Xsky130_fd_sc_hs__nand2_1_0 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_1_1/B sky130_fd_sc_hs__xnor2_1_1/A
+ eqn[8] sky130_fd_sc_hs__nand2_1_1/a_117_74# sky130_fd_sc_hs__nand2_1
Xsky130_fd_sc_hs__xnor2_1_15 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__xnor2_1_15/A sky130_fd_sc_hs__xnor2_1_29/B
+ sky130_fd_sc_hs__xnor2_1_15/B sky130_fd_sc_hs__xnor2_1_15/a_376_368# sky130_fd_sc_hs__xnor2_1_15/a_112_119#
+ sky130_fd_sc_hs__xnor2_1_15/a_138_385# sky130_fd_sc_hs__xnor2_1_15/a_293_74# sky130_fd_sc_hs__xnor2_1
Xsky130_fd_sc_hs__xnor2_1_26 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__xnor2_1_5/Y sky130_fd_sc_hs__xnor2_1_29/A
+ sky130_fd_sc_hs__xnor2_1_41/Y sky130_fd_sc_hs__xnor2_1_27/a_376_368# sky130_fd_sc_hs__xnor2_1_27/a_112_119#
+ sky130_fd_sc_hs__xnor2_1_27/a_138_385# sky130_fd_sc_hs__xnor2_1_27/a_293_74# sky130_fd_sc_hs__xnor2_1
Xsky130_fd_sc_hs__xnor2_1_37 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__xnor2_1_37/A sky130_fd_sc_hs__xnor2_1_50/A
+ sky130_fd_sc_hs__xnor2_1_37/B sky130_fd_sc_hs__xnor2_1_37/a_376_368# sky130_fd_sc_hs__xnor2_1_37/a_112_119#
+ sky130_fd_sc_hs__xnor2_1_37/a_138_385# sky130_fd_sc_hs__xnor2_1_37/a_293_74# sky130_fd_sc_hs__xnor2_1
Xsky130_fd_sc_hs__xnor2_1_48 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__xnor2_1_50/A sky130_fd_sc_hs__xnor2_1_50/Y
+ sky130_fd_sc_hs__xnor2_1_51/Y sky130_fd_sc_hs__xnor2_1_50/a_376_368# sky130_fd_sc_hs__xnor2_1_50/a_112_119#
+ sky130_fd_sc_hs__xnor2_1_50/a_138_385# sky130_fd_sc_hs__xnor2_1_50/a_293_74# sky130_fd_sc_hs__xnor2_1
Xsky130_fd_sc_hs__xnor2_1_59 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__xnor2_1_59/A sky130_fd_sc_hs__xnor2_1_59/Y
+ sky130_fd_sc_hs__xnor2_1_59/B sky130_fd_sc_hs__xnor2_1_59/a_376_368# sky130_fd_sc_hs__xnor2_1_59/a_112_119#
+ sky130_fd_sc_hs__xnor2_1_59/a_138_385# sky130_fd_sc_hs__xnor2_1_59/a_293_74# sky130_fd_sc_hs__xnor2_1
Xsky130_fd_sc_hs__sdlclkp_2_1 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__clkbuf_16_1/A clk
+ sky130_fd_sc_hs__or2_1_1/X sky130_fd_sc_hs__conb_1_1/LO sky130_fd_sc_hs__sdlclkp_2_1/a_114_112#
+ sky130_fd_sc_hs__sdlclkp_2_1/a_706_317# sky130_fd_sc_hs__sdlclkp_2_1/a_685_81# sky130_fd_sc_hs__sdlclkp_2_1/a_580_74#
+ sky130_fd_sc_hs__sdlclkp_2_1/a_288_48# sky130_fd_sc_hs__sdlclkp_2_1/a_114_424# sky130_fd_sc_hs__sdlclkp_2_1/a_1195_374#
+ sky130_fd_sc_hs__sdlclkp_2_1/a_708_451# sky130_fd_sc_hs__sdlclkp_2_1/a_1198_74#
+ sky130_fd_sc_hs__sdlclkp_2_1/a_318_74# sky130_fd_sc_hs__sdlclkp_2
Xsky130_fd_sc_hs__a22o_1_1 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__a22o_1_1/X sky130_fd_sc_hs__nand2_1_3/B
+ sky130_fd_sc_hs__and2b_2_1/X init_val[13] rst sky130_fd_sc_hs__a22o_1_1/a_222_392#
+ sky130_fd_sc_hs__a22o_1_1/a_230_79# sky130_fd_sc_hs__a22o_1_1/a_52_123# sky130_fd_sc_hs__a22o_1_1/a_132_392#
+ sky130_fd_sc_hs__a22o_1
Xsky130_fd_sc_hs__nand2_1_1 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_1_1/B sky130_fd_sc_hs__xnor2_1_1/A
+ eqn[8] sky130_fd_sc_hs__nand2_1_1/a_117_74# sky130_fd_sc_hs__nand2_1
Xsky130_fd_sc_hs__xnor2_1_16 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__xnor2_1_57/Y sky130_fd_sc_hs__xnor2_1_23/B
+ sky130_fd_sc_hs__xnor2_1_17/B sky130_fd_sc_hs__xnor2_1_17/a_376_368# sky130_fd_sc_hs__xnor2_1_17/a_112_119#
+ sky130_fd_sc_hs__xnor2_1_17/a_138_385# sky130_fd_sc_hs__xnor2_1_17/a_293_74# sky130_fd_sc_hs__xnor2_1
Xsky130_fd_sc_hs__xnor2_1_27 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__xnor2_1_5/Y sky130_fd_sc_hs__xnor2_1_29/A
+ sky130_fd_sc_hs__xnor2_1_41/Y sky130_fd_sc_hs__xnor2_1_27/a_376_368# sky130_fd_sc_hs__xnor2_1_27/a_112_119#
+ sky130_fd_sc_hs__xnor2_1_27/a_138_385# sky130_fd_sc_hs__xnor2_1_27/a_293_74# sky130_fd_sc_hs__xnor2_1
Xsky130_fd_sc_hs__xnor2_1_38 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__xnor2_1_50/Y sky130_fd_sc_hs__xnor2_1_41/A
+ sky130_fd_sc_hs__xnor2_1_39/B sky130_fd_sc_hs__xnor2_1_39/a_376_368# sky130_fd_sc_hs__xnor2_1_39/a_112_119#
+ sky130_fd_sc_hs__xnor2_1_39/a_138_385# sky130_fd_sc_hs__xnor2_1_39/a_293_74# sky130_fd_sc_hs__xnor2_1
Xsky130_fd_sc_hs__xnor2_1_49 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__xnor2_1_51/A sky130_fd_sc_hs__xnor2_1_51/Y
+ sky130_fd_sc_hs__xnor2_1_59/Y sky130_fd_sc_hs__xnor2_1_51/a_376_368# sky130_fd_sc_hs__xnor2_1_51/a_112_119#
+ sky130_fd_sc_hs__xnor2_1_51/a_138_385# sky130_fd_sc_hs__xnor2_1_51/a_293_74# sky130_fd_sc_hs__xnor2_1
Xsky130_fd_sc_hs__a22o_1_2 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__a22o_1_3/X sky130_fd_sc_hs__nand2_2_1/B
+ sky130_fd_sc_hs__and2b_2_1/X init_val[12] rst sky130_fd_sc_hs__a22o_1_3/a_222_392#
+ sky130_fd_sc_hs__a22o_1_3/a_230_79# sky130_fd_sc_hs__a22o_1_3/a_52_123# sky130_fd_sc_hs__a22o_1_3/a_132_392#
+ sky130_fd_sc_hs__a22o_1
Xsky130_fd_sc_hs__xnor2_1_17 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__xnor2_1_57/Y sky130_fd_sc_hs__xnor2_1_23/B
+ sky130_fd_sc_hs__xnor2_1_17/B sky130_fd_sc_hs__xnor2_1_17/a_376_368# sky130_fd_sc_hs__xnor2_1_17/a_112_119#
+ sky130_fd_sc_hs__xnor2_1_17/a_138_385# sky130_fd_sc_hs__xnor2_1_17/a_293_74# sky130_fd_sc_hs__xnor2_1
Xsky130_fd_sc_hs__xnor2_1_28 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__xnor2_1_29/A sky130_fd_sc_hs__xnor2_1_43/B
+ sky130_fd_sc_hs__xnor2_1_29/B sky130_fd_sc_hs__xnor2_1_29/a_376_368# sky130_fd_sc_hs__xnor2_1_29/a_112_119#
+ sky130_fd_sc_hs__xnor2_1_29/a_138_385# sky130_fd_sc_hs__xnor2_1_29/a_293_74# sky130_fd_sc_hs__xnor2_1
Xsky130_fd_sc_hs__xnor2_1_39 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__xnor2_1_50/Y sky130_fd_sc_hs__xnor2_1_41/A
+ sky130_fd_sc_hs__xnor2_1_39/B sky130_fd_sc_hs__xnor2_1_39/a_376_368# sky130_fd_sc_hs__xnor2_1_39/a_112_119#
+ sky130_fd_sc_hs__xnor2_1_39/a_138_385# sky130_fd_sc_hs__xnor2_1_39/a_293_74# sky130_fd_sc_hs__xnor2_1
Xsky130_fd_sc_hs__nor2b_1_0 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__xnor2_1_65/Y sky130_fd_sc_hs__nor2b_1_1/Y
+ rst sky130_fd_sc_hs__nor2b_1_1/a_278_368# sky130_fd_sc_hs__nor2b_1_1/a_27_112# sky130_fd_sc_hs__nor2b_1
Xsky130_fd_sc_hs__nand2_1_2 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_1_3/B sky130_fd_sc_hs__xnor2_1_3/B
+ eqn[12] sky130_fd_sc_hs__nand2_1_3/a_117_74# sky130_fd_sc_hs__nand2_1
Xsky130_fd_sc_hs__a22o_1_3 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__a22o_1_3/X sky130_fd_sc_hs__nand2_2_1/B
+ sky130_fd_sc_hs__and2b_2_1/X init_val[12] rst sky130_fd_sc_hs__a22o_1_3/a_222_392#
+ sky130_fd_sc_hs__a22o_1_3/a_230_79# sky130_fd_sc_hs__a22o_1_3/a_52_123# sky130_fd_sc_hs__a22o_1_3/a_132_392#
+ sky130_fd_sc_hs__a22o_1
Xsky130_fd_sc_hs__nor2b_1_1 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__xnor2_1_65/Y sky130_fd_sc_hs__nor2b_1_1/Y
+ rst sky130_fd_sc_hs__nor2b_1_1/a_278_368# sky130_fd_sc_hs__nor2b_1_1/a_27_112# sky130_fd_sc_hs__nor2b_1
Xsky130_fd_sc_hs__nand2_1_3 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_1_3/B sky130_fd_sc_hs__xnor2_1_3/B
+ eqn[12] sky130_fd_sc_hs__nand2_1_3/a_117_74# sky130_fd_sc_hs__nand2_1
Xsky130_fd_sc_hs__xnor2_1_18 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__xnor2_1_19/A sky130_fd_sc_hs__xnor2_1_51/A
+ sky130_fd_sc_hs__xnor2_1_19/B sky130_fd_sc_hs__xnor2_1_19/a_376_368# sky130_fd_sc_hs__xnor2_1_19/a_112_119#
+ sky130_fd_sc_hs__xnor2_1_19/a_138_385# sky130_fd_sc_hs__xnor2_1_19/a_293_74# sky130_fd_sc_hs__xnor2_1
Xsky130_fd_sc_hs__xnor2_1_29 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__xnor2_1_29/A sky130_fd_sc_hs__xnor2_1_43/B
+ sky130_fd_sc_hs__xnor2_1_29/B sky130_fd_sc_hs__xnor2_1_29/a_376_368# sky130_fd_sc_hs__xnor2_1_29/a_112_119#
+ sky130_fd_sc_hs__xnor2_1_29/a_138_385# sky130_fd_sc_hs__xnor2_1_29/a_293_74# sky130_fd_sc_hs__xnor2_1
Xsky130_fd_sc_hs__a22o_1_4 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__a22o_1_5/X sky130_fd_sc_hs__dfxtp_4_7/Q
+ sky130_fd_sc_hs__and2b_2_1/X init_val[11] rst sky130_fd_sc_hs__a22o_1_5/a_222_392#
+ sky130_fd_sc_hs__a22o_1_5/a_230_79# sky130_fd_sc_hs__a22o_1_5/a_52_123# sky130_fd_sc_hs__a22o_1_5/a_132_392#
+ sky130_fd_sc_hs__a22o_1
Xsky130_fd_sc_hs__nand2_1_4 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_1_5/B sky130_fd_sc_hs__xnor2_1_1/B
+ eqn[5] sky130_fd_sc_hs__nand2_1_5/a_117_74# sky130_fd_sc_hs__nand2_1
Xsky130_fd_sc_hs__xnor2_1_19 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__xnor2_1_19/A sky130_fd_sc_hs__xnor2_1_51/A
+ sky130_fd_sc_hs__xnor2_1_19/B sky130_fd_sc_hs__xnor2_1_19/a_376_368# sky130_fd_sc_hs__xnor2_1_19/a_112_119#
+ sky130_fd_sc_hs__xnor2_1_19/a_138_385# sky130_fd_sc_hs__xnor2_1_19/a_293_74# sky130_fd_sc_hs__xnor2_1
Xsky130_fd_sc_hs__nor2b_1_2 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__dfxtp_4_51/Q sky130_fd_sc_hs__nor2b_1_4/Y
+ sky130_fd_sc_hs__nor2b_1_4/A sky130_fd_sc_hs__nor2b_1_4/a_278_368# sky130_fd_sc_hs__nor2b_1_4/a_27_112#
+ sky130_fd_sc_hs__nor2b_1
Xsky130_fd_sc_hs__a22o_1_5 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__a22o_1_5/X sky130_fd_sc_hs__dfxtp_4_7/Q
+ sky130_fd_sc_hs__and2b_2_1/X init_val[11] rst sky130_fd_sc_hs__a22o_1_5/a_222_392#
+ sky130_fd_sc_hs__a22o_1_5/a_230_79# sky130_fd_sc_hs__a22o_1_5/a_52_123# sky130_fd_sc_hs__a22o_1_5/a_132_392#
+ sky130_fd_sc_hs__a22o_1
Xsky130_fd_sc_hs__nand2_1_5 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_1_5/B sky130_fd_sc_hs__xnor2_1_1/B
+ eqn[5] sky130_fd_sc_hs__nand2_1_5/a_117_74# sky130_fd_sc_hs__nand2_1
Xsky130_fd_sc_hs__nor2b_1_3 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__dfxtp_4_51/Q sky130_fd_sc_hs__nor2b_1_5/Y
+ rst sky130_fd_sc_hs__nor2b_1_5/a_278_368# sky130_fd_sc_hs__nor2b_1_5/a_27_112# sky130_fd_sc_hs__nor2b_1
Xsky130_fd_sc_hs__dfxtp_4_70 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__dfxtp_4_71/Q sky130_fd_sc_hs__nor2b_1_7/Y
+ sky130_fd_sc_hs__dfxtp_4_9/CLK sky130_fd_sc_hs__dfxtp_4_71/a_1226_296# sky130_fd_sc_hs__dfxtp_4_71/a_735_102#
+ sky130_fd_sc_hs__dfxtp_4_71/a_1141_508# sky130_fd_sc_hs__dfxtp_4_71/a_206_368# sky130_fd_sc_hs__dfxtp_4_71/a_437_503#
+ sky130_fd_sc_hs__dfxtp_4_71/a_27_74# sky130_fd_sc_hs__dfxtp_4_71/a_651_503# sky130_fd_sc_hs__dfxtp_4_71/a_696_458#
+ sky130_fd_sc_hs__dfxtp_4_71/a_544_485# sky130_fd_sc_hs__dfxtp_4_71/a_1178_124# sky130_fd_sc_hs__dfxtp_4_71/a_1034_424#
+ sky130_fd_sc_hs__dfxtp_4
Xsky130_fd_sc_hs__and2b_2_0 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__and2b_2_1/X cke rst
+ sky130_fd_sc_hs__and2b_2_1/a_505_74# sky130_fd_sc_hs__and2b_2_1/a_27_74# sky130_fd_sc_hs__and2b_2_1/a_198_48#
+ sky130_fd_sc_hs__and2b_2
Xsky130_fd_sc_hs__a22o_1_6 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__a22o_1_7/X sky130_fd_sc_hs__nand2_1_7/B
+ sky130_fd_sc_hs__and2b_2_1/X init_val[10] rst sky130_fd_sc_hs__a22o_1_7/a_222_392#
+ sky130_fd_sc_hs__a22o_1_7/a_230_79# sky130_fd_sc_hs__a22o_1_7/a_52_123# sky130_fd_sc_hs__a22o_1_7/a_132_392#
+ sky130_fd_sc_hs__a22o_1
Xsky130_fd_sc_hs__nand2_1_6 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_1_7/B sky130_fd_sc_hs__xnor2_1_9/A
+ eqn[9] sky130_fd_sc_hs__nand2_1_7/a_117_74# sky130_fd_sc_hs__nand2_1
Xsky130_fd_sc_hs__nor2b_1_4 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__dfxtp_4_51/Q sky130_fd_sc_hs__nor2b_1_4/Y
+ sky130_fd_sc_hs__nor2b_1_4/A sky130_fd_sc_hs__nor2b_1_4/a_278_368# sky130_fd_sc_hs__nor2b_1_4/a_27_112#
+ sky130_fd_sc_hs__nor2b_1
Xsky130_fd_sc_hs__dfxtp_4_71 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__dfxtp_4_71/Q sky130_fd_sc_hs__nor2b_1_7/Y
+ sky130_fd_sc_hs__dfxtp_4_9/CLK sky130_fd_sc_hs__dfxtp_4_71/a_1226_296# sky130_fd_sc_hs__dfxtp_4_71/a_735_102#
+ sky130_fd_sc_hs__dfxtp_4_71/a_1141_508# sky130_fd_sc_hs__dfxtp_4_71/a_206_368# sky130_fd_sc_hs__dfxtp_4_71/a_437_503#
+ sky130_fd_sc_hs__dfxtp_4_71/a_27_74# sky130_fd_sc_hs__dfxtp_4_71/a_651_503# sky130_fd_sc_hs__dfxtp_4_71/a_696_458#
+ sky130_fd_sc_hs__dfxtp_4_71/a_544_485# sky130_fd_sc_hs__dfxtp_4_71/a_1178_124# sky130_fd_sc_hs__dfxtp_4_71/a_1034_424#
+ sky130_fd_sc_hs__dfxtp_4
Xsky130_fd_sc_hs__dfxtp_4_60 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_1_39/B sky130_fd_sc_hs__a22o_1_59/X
+ sky130_fd_sc_hs__dfxtp_4_9/CLK sky130_fd_sc_hs__dfxtp_4_61/a_1226_296# sky130_fd_sc_hs__dfxtp_4_61/a_735_102#
+ sky130_fd_sc_hs__dfxtp_4_61/a_1141_508# sky130_fd_sc_hs__dfxtp_4_61/a_206_368# sky130_fd_sc_hs__dfxtp_4_61/a_437_503#
+ sky130_fd_sc_hs__dfxtp_4_61/a_27_74# sky130_fd_sc_hs__dfxtp_4_61/a_651_503# sky130_fd_sc_hs__dfxtp_4_61/a_696_458#
+ sky130_fd_sc_hs__dfxtp_4_61/a_544_485# sky130_fd_sc_hs__dfxtp_4_61/a_1178_124# sky130_fd_sc_hs__dfxtp_4_61/a_1034_424#
+ sky130_fd_sc_hs__dfxtp_4
Xsky130_fd_sc_hs__and2b_2_1 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__and2b_2_1/X cke rst
+ sky130_fd_sc_hs__and2b_2_1/a_505_74# sky130_fd_sc_hs__and2b_2_1/a_27_74# sky130_fd_sc_hs__and2b_2_1/a_198_48#
+ sky130_fd_sc_hs__and2b_2
Xsky130_fd_sc_hs__a22o_1_7 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__a22o_1_7/X sky130_fd_sc_hs__nand2_1_7/B
+ sky130_fd_sc_hs__and2b_2_1/X init_val[10] rst sky130_fd_sc_hs__a22o_1_7/a_222_392#
+ sky130_fd_sc_hs__a22o_1_7/a_230_79# sky130_fd_sc_hs__a22o_1_7/a_52_123# sky130_fd_sc_hs__a22o_1_7/a_132_392#
+ sky130_fd_sc_hs__a22o_1
Xsky130_fd_sc_hs__nor2b_1_5 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__dfxtp_4_51/Q sky130_fd_sc_hs__nor2b_1_5/Y
+ rst sky130_fd_sc_hs__nor2b_1_5/a_278_368# sky130_fd_sc_hs__nor2b_1_5/a_27_112# sky130_fd_sc_hs__nor2b_1
Xsky130_fd_sc_hs__nand2_1_7 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_1_7/B sky130_fd_sc_hs__xnor2_1_9/A
+ eqn[9] sky130_fd_sc_hs__nand2_1_7/a_117_74# sky130_fd_sc_hs__nand2_1
Xsky130_fd_sc_hs__clkbuf_16_0 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__dfxtp_4_9/CLK sky130_fd_sc_hs__clkbuf_16_1/A
+ sky130_fd_sc_hs__clkbuf_16_1/a_114_74# sky130_fd_sc_hs__clkbuf_16
Xsky130_fd_sc_hs__dfxtp_4_72 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_1_53/B sky130_fd_sc_hs__a22o_1_61/X
+ sky130_fd_sc_hs__dfxtp_4_9/CLK sky130_fd_sc_hs__dfxtp_4_73/a_1226_296# sky130_fd_sc_hs__dfxtp_4_73/a_735_102#
+ sky130_fd_sc_hs__dfxtp_4_73/a_1141_508# sky130_fd_sc_hs__dfxtp_4_73/a_206_368# sky130_fd_sc_hs__dfxtp_4_73/a_437_503#
+ sky130_fd_sc_hs__dfxtp_4_73/a_27_74# sky130_fd_sc_hs__dfxtp_4_73/a_651_503# sky130_fd_sc_hs__dfxtp_4_73/a_696_458#
+ sky130_fd_sc_hs__dfxtp_4_73/a_544_485# sky130_fd_sc_hs__dfxtp_4_73/a_1178_124# sky130_fd_sc_hs__dfxtp_4_73/a_1034_424#
+ sky130_fd_sc_hs__dfxtp_4
Xsky130_fd_sc_hs__dfxtp_4_61 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_1_39/B sky130_fd_sc_hs__a22o_1_59/X
+ sky130_fd_sc_hs__dfxtp_4_9/CLK sky130_fd_sc_hs__dfxtp_4_61/a_1226_296# sky130_fd_sc_hs__dfxtp_4_61/a_735_102#
+ sky130_fd_sc_hs__dfxtp_4_61/a_1141_508# sky130_fd_sc_hs__dfxtp_4_61/a_206_368# sky130_fd_sc_hs__dfxtp_4_61/a_437_503#
+ sky130_fd_sc_hs__dfxtp_4_61/a_27_74# sky130_fd_sc_hs__dfxtp_4_61/a_651_503# sky130_fd_sc_hs__dfxtp_4_61/a_696_458#
+ sky130_fd_sc_hs__dfxtp_4_61/a_544_485# sky130_fd_sc_hs__dfxtp_4_61/a_1178_124# sky130_fd_sc_hs__dfxtp_4_61/a_1034_424#
+ sky130_fd_sc_hs__dfxtp_4
Xsky130_fd_sc_hs__dfxtp_4_50 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__dfxtp_4_51/Q sky130_fd_sc_hs__nor2b_1_9/Y
+ sky130_fd_sc_hs__dfxtp_4_9/CLK sky130_fd_sc_hs__dfxtp_4_51/a_1226_296# sky130_fd_sc_hs__dfxtp_4_51/a_735_102#
+ sky130_fd_sc_hs__dfxtp_4_51/a_1141_508# sky130_fd_sc_hs__dfxtp_4_51/a_206_368# sky130_fd_sc_hs__dfxtp_4_51/a_437_503#
+ sky130_fd_sc_hs__dfxtp_4_51/a_27_74# sky130_fd_sc_hs__dfxtp_4_51/a_651_503# sky130_fd_sc_hs__dfxtp_4_51/a_696_458#
+ sky130_fd_sc_hs__dfxtp_4_51/a_544_485# sky130_fd_sc_hs__dfxtp_4_51/a_1178_124# sky130_fd_sc_hs__dfxtp_4_51/a_1034_424#
+ sky130_fd_sc_hs__dfxtp_4
Xsky130_fd_sc_hs__a22o_1_8 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__a22o_1_9/X sky130_fd_sc_hs__nand2_1_1/B
+ sky130_fd_sc_hs__and2b_2_1/X init_val[9] rst sky130_fd_sc_hs__a22o_1_9/a_222_392#
+ sky130_fd_sc_hs__a22o_1_9/a_230_79# sky130_fd_sc_hs__a22o_1_9/a_52_123# sky130_fd_sc_hs__a22o_1_9/a_132_392#
+ sky130_fd_sc_hs__a22o_1
Xsky130_fd_sc_hs__nor2b_1_6 DVSS DVDD DVDD DVSS inj_err sky130_fd_sc_hs__nor2b_1_7/Y
+ rst sky130_fd_sc_hs__nor2b_1_7/a_278_368# sky130_fd_sc_hs__nor2b_1_7/a_27_112# sky130_fd_sc_hs__nor2b_1
Xsky130_fd_sc_hs__nand2_1_8 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_1_9/B sky130_fd_sc_hs__xnor2_1_9/B
+ eqn[4] sky130_fd_sc_hs__nand2_1_9/a_117_74# sky130_fd_sc_hs__nand2_1
Xsky130_fd_sc_hs__clkbuf_16_1 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__dfxtp_4_9/CLK sky130_fd_sc_hs__clkbuf_16_1/A
+ sky130_fd_sc_hs__clkbuf_16_1/a_114_74# sky130_fd_sc_hs__clkbuf_16
Xsky130_fd_sc_hs__dfxtp_4_40 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_1_41/B sky130_fd_sc_hs__a22o_1_37/X
+ sky130_fd_sc_hs__dfxtp_4_9/CLK sky130_fd_sc_hs__dfxtp_4_41/a_1226_296# sky130_fd_sc_hs__dfxtp_4_41/a_735_102#
+ sky130_fd_sc_hs__dfxtp_4_41/a_1141_508# sky130_fd_sc_hs__dfxtp_4_41/a_206_368# sky130_fd_sc_hs__dfxtp_4_41/a_437_503#
+ sky130_fd_sc_hs__dfxtp_4_41/a_27_74# sky130_fd_sc_hs__dfxtp_4_41/a_651_503# sky130_fd_sc_hs__dfxtp_4_41/a_696_458#
+ sky130_fd_sc_hs__dfxtp_4_41/a_544_485# sky130_fd_sc_hs__dfxtp_4_41/a_1178_124# sky130_fd_sc_hs__dfxtp_4_41/a_1034_424#
+ sky130_fd_sc_hs__dfxtp_4
Xsky130_fd_sc_hs__dfxtp_4_73 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_1_53/B sky130_fd_sc_hs__a22o_1_61/X
+ sky130_fd_sc_hs__dfxtp_4_9/CLK sky130_fd_sc_hs__dfxtp_4_73/a_1226_296# sky130_fd_sc_hs__dfxtp_4_73/a_735_102#
+ sky130_fd_sc_hs__dfxtp_4_73/a_1141_508# sky130_fd_sc_hs__dfxtp_4_73/a_206_368# sky130_fd_sc_hs__dfxtp_4_73/a_437_503#
+ sky130_fd_sc_hs__dfxtp_4_73/a_27_74# sky130_fd_sc_hs__dfxtp_4_73/a_651_503# sky130_fd_sc_hs__dfxtp_4_73/a_696_458#
+ sky130_fd_sc_hs__dfxtp_4_73/a_544_485# sky130_fd_sc_hs__dfxtp_4_73/a_1178_124# sky130_fd_sc_hs__dfxtp_4_73/a_1034_424#
+ sky130_fd_sc_hs__dfxtp_4
Xsky130_fd_sc_hs__dfxtp_4_62 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__dfxtp_4_63/Q sky130_fd_sc_hs__nor2b_1_8/Y
+ sky130_fd_sc_hs__dfxtp_4_9/CLK sky130_fd_sc_hs__dfxtp_4_63/a_1226_296# sky130_fd_sc_hs__dfxtp_4_63/a_735_102#
+ sky130_fd_sc_hs__dfxtp_4_63/a_1141_508# sky130_fd_sc_hs__dfxtp_4_63/a_206_368# sky130_fd_sc_hs__dfxtp_4_63/a_437_503#
+ sky130_fd_sc_hs__dfxtp_4_63/a_27_74# sky130_fd_sc_hs__dfxtp_4_63/a_651_503# sky130_fd_sc_hs__dfxtp_4_63/a_696_458#
+ sky130_fd_sc_hs__dfxtp_4_63/a_544_485# sky130_fd_sc_hs__dfxtp_4_63/a_1178_124# sky130_fd_sc_hs__dfxtp_4_63/a_1034_424#
+ sky130_fd_sc_hs__dfxtp_4
Xsky130_fd_sc_hs__dfxtp_4_51 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__dfxtp_4_51/Q sky130_fd_sc_hs__nor2b_1_9/Y
+ sky130_fd_sc_hs__dfxtp_4_9/CLK sky130_fd_sc_hs__dfxtp_4_51/a_1226_296# sky130_fd_sc_hs__dfxtp_4_51/a_735_102#
+ sky130_fd_sc_hs__dfxtp_4_51/a_1141_508# sky130_fd_sc_hs__dfxtp_4_51/a_206_368# sky130_fd_sc_hs__dfxtp_4_51/a_437_503#
+ sky130_fd_sc_hs__dfxtp_4_51/a_27_74# sky130_fd_sc_hs__dfxtp_4_51/a_651_503# sky130_fd_sc_hs__dfxtp_4_51/a_696_458#
+ sky130_fd_sc_hs__dfxtp_4_51/a_544_485# sky130_fd_sc_hs__dfxtp_4_51/a_1178_124# sky130_fd_sc_hs__dfxtp_4_51/a_1034_424#
+ sky130_fd_sc_hs__dfxtp_4
Xsky130_fd_sc_hs__a22o_1_9 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__a22o_1_9/X sky130_fd_sc_hs__nand2_1_1/B
+ sky130_fd_sc_hs__and2b_2_1/X init_val[9] rst sky130_fd_sc_hs__a22o_1_9/a_222_392#
+ sky130_fd_sc_hs__a22o_1_9/a_230_79# sky130_fd_sc_hs__a22o_1_9/a_52_123# sky130_fd_sc_hs__a22o_1_9/a_132_392#
+ sky130_fd_sc_hs__a22o_1
Xsky130_fd_sc_hs__nand2_1_9 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_1_9/B sky130_fd_sc_hs__xnor2_1_9/B
+ eqn[4] sky130_fd_sc_hs__nand2_1_9/a_117_74# sky130_fd_sc_hs__nand2_1
Xsky130_fd_sc_hs__nor2b_1_7 DVSS DVDD DVDD DVSS inj_err sky130_fd_sc_hs__nor2b_1_7/Y
+ rst sky130_fd_sc_hs__nor2b_1_7/a_278_368# sky130_fd_sc_hs__nor2b_1_7/a_27_112# sky130_fd_sc_hs__nor2b_1
Xsky130_fd_sc_hs__dfxtp_4_30 DVSS DVDD DVDD DVSS out sky130_fd_sc_hs__nor2b_1_1/Y
+ sky130_fd_sc_hs__dfxtp_4_9/CLK sky130_fd_sc_hs__dfxtp_4_32/a_1226_296# sky130_fd_sc_hs__dfxtp_4_32/a_735_102#
+ sky130_fd_sc_hs__dfxtp_4_32/a_1141_508# sky130_fd_sc_hs__dfxtp_4_32/a_206_368# sky130_fd_sc_hs__dfxtp_4_32/a_437_503#
+ sky130_fd_sc_hs__dfxtp_4_32/a_27_74# sky130_fd_sc_hs__dfxtp_4_32/a_651_503# sky130_fd_sc_hs__dfxtp_4_32/a_696_458#
+ sky130_fd_sc_hs__dfxtp_4_32/a_544_485# sky130_fd_sc_hs__dfxtp_4_32/a_1178_124# sky130_fd_sc_hs__dfxtp_4_32/a_1034_424#
+ sky130_fd_sc_hs__dfxtp_4
Xsky130_fd_sc_hs__dfxtp_4_41 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_1_41/B sky130_fd_sc_hs__a22o_1_37/X
+ sky130_fd_sc_hs__dfxtp_4_9/CLK sky130_fd_sc_hs__dfxtp_4_41/a_1226_296# sky130_fd_sc_hs__dfxtp_4_41/a_735_102#
+ sky130_fd_sc_hs__dfxtp_4_41/a_1141_508# sky130_fd_sc_hs__dfxtp_4_41/a_206_368# sky130_fd_sc_hs__dfxtp_4_41/a_437_503#
+ sky130_fd_sc_hs__dfxtp_4_41/a_27_74# sky130_fd_sc_hs__dfxtp_4_41/a_651_503# sky130_fd_sc_hs__dfxtp_4_41/a_696_458#
+ sky130_fd_sc_hs__dfxtp_4_41/a_544_485# sky130_fd_sc_hs__dfxtp_4_41/a_1178_124# sky130_fd_sc_hs__dfxtp_4_41/a_1034_424#
+ sky130_fd_sc_hs__dfxtp_4
Xsky130_fd_sc_hs__dfxtp_4_63 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__dfxtp_4_63/Q sky130_fd_sc_hs__nor2b_1_8/Y
+ sky130_fd_sc_hs__dfxtp_4_9/CLK sky130_fd_sc_hs__dfxtp_4_63/a_1226_296# sky130_fd_sc_hs__dfxtp_4_63/a_735_102#
+ sky130_fd_sc_hs__dfxtp_4_63/a_1141_508# sky130_fd_sc_hs__dfxtp_4_63/a_206_368# sky130_fd_sc_hs__dfxtp_4_63/a_437_503#
+ sky130_fd_sc_hs__dfxtp_4_63/a_27_74# sky130_fd_sc_hs__dfxtp_4_63/a_651_503# sky130_fd_sc_hs__dfxtp_4_63/a_696_458#
+ sky130_fd_sc_hs__dfxtp_4_63/a_544_485# sky130_fd_sc_hs__dfxtp_4_63/a_1178_124# sky130_fd_sc_hs__dfxtp_4_63/a_1034_424#
+ sky130_fd_sc_hs__dfxtp_4
Xsky130_fd_sc_hs__dfxtp_4_52 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_1_51/B sky130_fd_sc_hs__a22o_1_49/X
+ sky130_fd_sc_hs__dfxtp_4_9/CLK sky130_fd_sc_hs__dfxtp_4_53/a_1226_296# sky130_fd_sc_hs__dfxtp_4_53/a_735_102#
+ sky130_fd_sc_hs__dfxtp_4_53/a_1141_508# sky130_fd_sc_hs__dfxtp_4_53/a_206_368# sky130_fd_sc_hs__dfxtp_4_53/a_437_503#
+ sky130_fd_sc_hs__dfxtp_4_53/a_27_74# sky130_fd_sc_hs__dfxtp_4_53/a_651_503# sky130_fd_sc_hs__dfxtp_4_53/a_696_458#
+ sky130_fd_sc_hs__dfxtp_4_53/a_544_485# sky130_fd_sc_hs__dfxtp_4_53/a_1178_124# sky130_fd_sc_hs__dfxtp_4_53/a_1034_424#
+ sky130_fd_sc_hs__dfxtp_4
Xsky130_fd_sc_hs__nor2b_1_8 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__dfxtp_4_71/Q sky130_fd_sc_hs__nor2b_1_8/Y
+ rst sky130_fd_sc_hs__nor2b_1_8/a_278_368# sky130_fd_sc_hs__nor2b_1_8/a_27_112# sky130_fd_sc_hs__nor2b_1
Xsky130_fd_sc_hs__dfxtp_4_20 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_1_31/B sky130_fd_sc_hs__a22o_1_21/X
+ sky130_fd_sc_hs__dfxtp_4_9/CLK sky130_fd_sc_hs__dfxtp_4_21/a_1226_296# sky130_fd_sc_hs__dfxtp_4_21/a_735_102#
+ sky130_fd_sc_hs__dfxtp_4_21/a_1141_508# sky130_fd_sc_hs__dfxtp_4_21/a_206_368# sky130_fd_sc_hs__dfxtp_4_21/a_437_503#
+ sky130_fd_sc_hs__dfxtp_4_21/a_27_74# sky130_fd_sc_hs__dfxtp_4_21/a_651_503# sky130_fd_sc_hs__dfxtp_4_21/a_696_458#
+ sky130_fd_sc_hs__dfxtp_4_21/a_544_485# sky130_fd_sc_hs__dfxtp_4_21/a_1178_124# sky130_fd_sc_hs__dfxtp_4_21/a_1034_424#
+ sky130_fd_sc_hs__dfxtp_4
Xsky130_fd_sc_hs__dfxtp_4_31 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_1_47/B sky130_fd_sc_hs__a22o_1_41/X
+ sky130_fd_sc_hs__dfxtp_4_9/CLK sky130_fd_sc_hs__dfxtp_4_33/a_1226_296# sky130_fd_sc_hs__dfxtp_4_33/a_735_102#
+ sky130_fd_sc_hs__dfxtp_4_33/a_1141_508# sky130_fd_sc_hs__dfxtp_4_33/a_206_368# sky130_fd_sc_hs__dfxtp_4_33/a_437_503#
+ sky130_fd_sc_hs__dfxtp_4_33/a_27_74# sky130_fd_sc_hs__dfxtp_4_33/a_651_503# sky130_fd_sc_hs__dfxtp_4_33/a_696_458#
+ sky130_fd_sc_hs__dfxtp_4_33/a_544_485# sky130_fd_sc_hs__dfxtp_4_33/a_1178_124# sky130_fd_sc_hs__dfxtp_4_33/a_1034_424#
+ sky130_fd_sc_hs__dfxtp_4
Xsky130_fd_sc_hs__dfxtp_4_42 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_1_23/B sky130_fd_sc_hs__a22o_1_33/X
+ sky130_fd_sc_hs__dfxtp_4_9/CLK sky130_fd_sc_hs__dfxtp_4_43/a_1226_296# sky130_fd_sc_hs__dfxtp_4_43/a_735_102#
+ sky130_fd_sc_hs__dfxtp_4_43/a_1141_508# sky130_fd_sc_hs__dfxtp_4_43/a_206_368# sky130_fd_sc_hs__dfxtp_4_43/a_437_503#
+ sky130_fd_sc_hs__dfxtp_4_43/a_27_74# sky130_fd_sc_hs__dfxtp_4_43/a_651_503# sky130_fd_sc_hs__dfxtp_4_43/a_696_458#
+ sky130_fd_sc_hs__dfxtp_4_43/a_544_485# sky130_fd_sc_hs__dfxtp_4_43/a_1178_124# sky130_fd_sc_hs__dfxtp_4_43/a_1034_424#
+ sky130_fd_sc_hs__dfxtp_4
Xsky130_fd_sc_hs__dfxtp_4_64 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_1_37/B sky130_fd_sc_hs__a22o_1_53/X
+ sky130_fd_sc_hs__dfxtp_4_9/CLK sky130_fd_sc_hs__dfxtp_4_65/a_1226_296# sky130_fd_sc_hs__dfxtp_4_65/a_735_102#
+ sky130_fd_sc_hs__dfxtp_4_65/a_1141_508# sky130_fd_sc_hs__dfxtp_4_65/a_206_368# sky130_fd_sc_hs__dfxtp_4_65/a_437_503#
+ sky130_fd_sc_hs__dfxtp_4_65/a_27_74# sky130_fd_sc_hs__dfxtp_4_65/a_651_503# sky130_fd_sc_hs__dfxtp_4_65/a_696_458#
+ sky130_fd_sc_hs__dfxtp_4_65/a_544_485# sky130_fd_sc_hs__dfxtp_4_65/a_1178_124# sky130_fd_sc_hs__dfxtp_4_65/a_1034_424#
+ sky130_fd_sc_hs__dfxtp_4
Xsky130_fd_sc_hs__dfxtp_4_53 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_1_51/B sky130_fd_sc_hs__a22o_1_49/X
+ sky130_fd_sc_hs__dfxtp_4_9/CLK sky130_fd_sc_hs__dfxtp_4_53/a_1226_296# sky130_fd_sc_hs__dfxtp_4_53/a_735_102#
+ sky130_fd_sc_hs__dfxtp_4_53/a_1141_508# sky130_fd_sc_hs__dfxtp_4_53/a_206_368# sky130_fd_sc_hs__dfxtp_4_53/a_437_503#
+ sky130_fd_sc_hs__dfxtp_4_53/a_27_74# sky130_fd_sc_hs__dfxtp_4_53/a_651_503# sky130_fd_sc_hs__dfxtp_4_53/a_696_458#
+ sky130_fd_sc_hs__dfxtp_4_53/a_544_485# sky130_fd_sc_hs__dfxtp_4_53/a_1178_124# sky130_fd_sc_hs__dfxtp_4_53/a_1034_424#
+ sky130_fd_sc_hs__dfxtp_4
Xsky130_fd_sc_hs__nor2b_1_9 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__dfxtp_4_63/Q sky130_fd_sc_hs__nor2b_1_9/Y
+ rst sky130_fd_sc_hs__nor2b_1_9/a_278_368# sky130_fd_sc_hs__nor2b_1_9/a_27_112# sky130_fd_sc_hs__nor2b_1
Xsky130_fd_sc_hs__dfxtp_4_10 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_1_1/B sky130_fd_sc_hs__dfxtp_4_8/D
+ sky130_fd_sc_hs__dfxtp_4_9/CLK sky130_fd_sc_hs__dfxtp_4_8/a_1226_296# sky130_fd_sc_hs__dfxtp_4_8/a_735_102#
+ sky130_fd_sc_hs__dfxtp_4_8/a_1141_508# sky130_fd_sc_hs__dfxtp_4_8/a_206_368# sky130_fd_sc_hs__dfxtp_4_8/a_437_503#
+ sky130_fd_sc_hs__dfxtp_4_8/a_27_74# sky130_fd_sc_hs__dfxtp_4_8/a_651_503# sky130_fd_sc_hs__dfxtp_4_8/a_696_458#
+ sky130_fd_sc_hs__dfxtp_4_8/a_544_485# sky130_fd_sc_hs__dfxtp_4_8/a_1178_124# sky130_fd_sc_hs__dfxtp_4_8/a_1034_424#
+ sky130_fd_sc_hs__dfxtp_4
Xsky130_fd_sc_hs__dfxtp_4_21 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_1_31/B sky130_fd_sc_hs__a22o_1_21/X
+ sky130_fd_sc_hs__dfxtp_4_9/CLK sky130_fd_sc_hs__dfxtp_4_21/a_1226_296# sky130_fd_sc_hs__dfxtp_4_21/a_735_102#
+ sky130_fd_sc_hs__dfxtp_4_21/a_1141_508# sky130_fd_sc_hs__dfxtp_4_21/a_206_368# sky130_fd_sc_hs__dfxtp_4_21/a_437_503#
+ sky130_fd_sc_hs__dfxtp_4_21/a_27_74# sky130_fd_sc_hs__dfxtp_4_21/a_651_503# sky130_fd_sc_hs__dfxtp_4_21/a_696_458#
+ sky130_fd_sc_hs__dfxtp_4_21/a_544_485# sky130_fd_sc_hs__dfxtp_4_21/a_1178_124# sky130_fd_sc_hs__dfxtp_4_21/a_1034_424#
+ sky130_fd_sc_hs__dfxtp_4
Xsky130_fd_sc_hs__dfxtp_4_32 DVSS DVDD DVDD DVSS out sky130_fd_sc_hs__nor2b_1_1/Y
+ sky130_fd_sc_hs__dfxtp_4_9/CLK sky130_fd_sc_hs__dfxtp_4_32/a_1226_296# sky130_fd_sc_hs__dfxtp_4_32/a_735_102#
+ sky130_fd_sc_hs__dfxtp_4_32/a_1141_508# sky130_fd_sc_hs__dfxtp_4_32/a_206_368# sky130_fd_sc_hs__dfxtp_4_32/a_437_503#
+ sky130_fd_sc_hs__dfxtp_4_32/a_27_74# sky130_fd_sc_hs__dfxtp_4_32/a_651_503# sky130_fd_sc_hs__dfxtp_4_32/a_696_458#
+ sky130_fd_sc_hs__dfxtp_4_32/a_544_485# sky130_fd_sc_hs__dfxtp_4_32/a_1178_124# sky130_fd_sc_hs__dfxtp_4_32/a_1034_424#
+ sky130_fd_sc_hs__dfxtp_4
Xsky130_fd_sc_hs__dfxtp_4_43 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_1_23/B sky130_fd_sc_hs__a22o_1_33/X
+ sky130_fd_sc_hs__dfxtp_4_9/CLK sky130_fd_sc_hs__dfxtp_4_43/a_1226_296# sky130_fd_sc_hs__dfxtp_4_43/a_735_102#
+ sky130_fd_sc_hs__dfxtp_4_43/a_1141_508# sky130_fd_sc_hs__dfxtp_4_43/a_206_368# sky130_fd_sc_hs__dfxtp_4_43/a_437_503#
+ sky130_fd_sc_hs__dfxtp_4_43/a_27_74# sky130_fd_sc_hs__dfxtp_4_43/a_651_503# sky130_fd_sc_hs__dfxtp_4_43/a_696_458#
+ sky130_fd_sc_hs__dfxtp_4_43/a_544_485# sky130_fd_sc_hs__dfxtp_4_43/a_1178_124# sky130_fd_sc_hs__dfxtp_4_43/a_1034_424#
+ sky130_fd_sc_hs__dfxtp_4
Xsky130_fd_sc_hs__dfxtp_4_65 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_1_37/B sky130_fd_sc_hs__a22o_1_53/X
+ sky130_fd_sc_hs__dfxtp_4_9/CLK sky130_fd_sc_hs__dfxtp_4_65/a_1226_296# sky130_fd_sc_hs__dfxtp_4_65/a_735_102#
+ sky130_fd_sc_hs__dfxtp_4_65/a_1141_508# sky130_fd_sc_hs__dfxtp_4_65/a_206_368# sky130_fd_sc_hs__dfxtp_4_65/a_437_503#
+ sky130_fd_sc_hs__dfxtp_4_65/a_27_74# sky130_fd_sc_hs__dfxtp_4_65/a_651_503# sky130_fd_sc_hs__dfxtp_4_65/a_696_458#
+ sky130_fd_sc_hs__dfxtp_4_65/a_544_485# sky130_fd_sc_hs__dfxtp_4_65/a_1178_124# sky130_fd_sc_hs__dfxtp_4_65/a_1034_424#
+ sky130_fd_sc_hs__dfxtp_4
Xsky130_fd_sc_hs__dfxtp_4_54 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_1_55/B sky130_fd_sc_hs__a22o_1_47/X
+ sky130_fd_sc_hs__dfxtp_4_9/CLK sky130_fd_sc_hs__dfxtp_4_55/a_1226_296# sky130_fd_sc_hs__dfxtp_4_55/a_735_102#
+ sky130_fd_sc_hs__dfxtp_4_55/a_1141_508# sky130_fd_sc_hs__dfxtp_4_55/a_206_368# sky130_fd_sc_hs__dfxtp_4_55/a_437_503#
+ sky130_fd_sc_hs__dfxtp_4_55/a_27_74# sky130_fd_sc_hs__dfxtp_4_55/a_651_503# sky130_fd_sc_hs__dfxtp_4_55/a_696_458#
+ sky130_fd_sc_hs__dfxtp_4_55/a_544_485# sky130_fd_sc_hs__dfxtp_4_55/a_1178_124# sky130_fd_sc_hs__dfxtp_4_55/a_1034_424#
+ sky130_fd_sc_hs__dfxtp_4
Xsky130_fd_sc_hs__dfxtp_4_11 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_1_7/B sky130_fd_sc_hs__a22o_1_9/X
+ sky130_fd_sc_hs__dfxtp_4_9/CLK sky130_fd_sc_hs__dfxtp_4_9/a_1226_296# sky130_fd_sc_hs__dfxtp_4_9/a_735_102#
+ sky130_fd_sc_hs__dfxtp_4_9/a_1141_508# sky130_fd_sc_hs__dfxtp_4_9/a_206_368# sky130_fd_sc_hs__dfxtp_4_9/a_437_503#
+ sky130_fd_sc_hs__dfxtp_4_9/a_27_74# sky130_fd_sc_hs__dfxtp_4_9/a_651_503# sky130_fd_sc_hs__dfxtp_4_9/a_696_458#
+ sky130_fd_sc_hs__dfxtp_4_9/a_544_485# sky130_fd_sc_hs__dfxtp_4_9/a_1178_124# sky130_fd_sc_hs__dfxtp_4_9/a_1034_424#
+ sky130_fd_sc_hs__dfxtp_4
Xsky130_fd_sc_hs__dfxtp_4_22 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_1_5/B sky130_fd_sc_hs__a22o_1_25/X
+ sky130_fd_sc_hs__dfxtp_4_9/CLK sky130_fd_sc_hs__dfxtp_4_23/a_1226_296# sky130_fd_sc_hs__dfxtp_4_23/a_735_102#
+ sky130_fd_sc_hs__dfxtp_4_23/a_1141_508# sky130_fd_sc_hs__dfxtp_4_23/a_206_368# sky130_fd_sc_hs__dfxtp_4_23/a_437_503#
+ sky130_fd_sc_hs__dfxtp_4_23/a_27_74# sky130_fd_sc_hs__dfxtp_4_23/a_651_503# sky130_fd_sc_hs__dfxtp_4_23/a_696_458#
+ sky130_fd_sc_hs__dfxtp_4_23/a_544_485# sky130_fd_sc_hs__dfxtp_4_23/a_1178_124# sky130_fd_sc_hs__dfxtp_4_23/a_1034_424#
+ sky130_fd_sc_hs__dfxtp_4
Xsky130_fd_sc_hs__dfxtp_4_33 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_1_47/B sky130_fd_sc_hs__a22o_1_41/X
+ sky130_fd_sc_hs__dfxtp_4_9/CLK sky130_fd_sc_hs__dfxtp_4_33/a_1226_296# sky130_fd_sc_hs__dfxtp_4_33/a_735_102#
+ sky130_fd_sc_hs__dfxtp_4_33/a_1141_508# sky130_fd_sc_hs__dfxtp_4_33/a_206_368# sky130_fd_sc_hs__dfxtp_4_33/a_437_503#
+ sky130_fd_sc_hs__dfxtp_4_33/a_27_74# sky130_fd_sc_hs__dfxtp_4_33/a_651_503# sky130_fd_sc_hs__dfxtp_4_33/a_696_458#
+ sky130_fd_sc_hs__dfxtp_4_33/a_544_485# sky130_fd_sc_hs__dfxtp_4_33/a_1178_124# sky130_fd_sc_hs__dfxtp_4_33/a_1034_424#
+ sky130_fd_sc_hs__dfxtp_4
Xsky130_fd_sc_hs__dfxtp_4_66 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_2_3/B sky130_fd_sc_hs__a22o_1_57/X
+ sky130_fd_sc_hs__dfxtp_4_9/CLK sky130_fd_sc_hs__dfxtp_4_67/a_1226_296# sky130_fd_sc_hs__dfxtp_4_67/a_735_102#
+ sky130_fd_sc_hs__dfxtp_4_67/a_1141_508# sky130_fd_sc_hs__dfxtp_4_67/a_206_368# sky130_fd_sc_hs__dfxtp_4_67/a_437_503#
+ sky130_fd_sc_hs__dfxtp_4_67/a_27_74# sky130_fd_sc_hs__dfxtp_4_67/a_651_503# sky130_fd_sc_hs__dfxtp_4_67/a_696_458#
+ sky130_fd_sc_hs__dfxtp_4_67/a_544_485# sky130_fd_sc_hs__dfxtp_4_67/a_1178_124# sky130_fd_sc_hs__dfxtp_4_67/a_1034_424#
+ sky130_fd_sc_hs__dfxtp_4
Xsky130_fd_sc_hs__dfxtp_4_55 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_1_55/B sky130_fd_sc_hs__a22o_1_47/X
+ sky130_fd_sc_hs__dfxtp_4_9/CLK sky130_fd_sc_hs__dfxtp_4_55/a_1226_296# sky130_fd_sc_hs__dfxtp_4_55/a_735_102#
+ sky130_fd_sc_hs__dfxtp_4_55/a_1141_508# sky130_fd_sc_hs__dfxtp_4_55/a_206_368# sky130_fd_sc_hs__dfxtp_4_55/a_437_503#
+ sky130_fd_sc_hs__dfxtp_4_55/a_27_74# sky130_fd_sc_hs__dfxtp_4_55/a_651_503# sky130_fd_sc_hs__dfxtp_4_55/a_696_458#
+ sky130_fd_sc_hs__dfxtp_4_55/a_544_485# sky130_fd_sc_hs__dfxtp_4_55/a_1178_124# sky130_fd_sc_hs__dfxtp_4_55/a_1034_424#
+ sky130_fd_sc_hs__dfxtp_4
Xsky130_fd_sc_hs__dfxtp_4_44 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_1_45/B sky130_fd_sc_hs__a22o_1_45/X
+ sky130_fd_sc_hs__dfxtp_4_9/CLK sky130_fd_sc_hs__dfxtp_4_45/a_1226_296# sky130_fd_sc_hs__dfxtp_4_45/a_735_102#
+ sky130_fd_sc_hs__dfxtp_4_45/a_1141_508# sky130_fd_sc_hs__dfxtp_4_45/a_206_368# sky130_fd_sc_hs__dfxtp_4_45/a_437_503#
+ sky130_fd_sc_hs__dfxtp_4_45/a_27_74# sky130_fd_sc_hs__dfxtp_4_45/a_651_503# sky130_fd_sc_hs__dfxtp_4_45/a_696_458#
+ sky130_fd_sc_hs__dfxtp_4_45/a_544_485# sky130_fd_sc_hs__dfxtp_4_45/a_1178_124# sky130_fd_sc_hs__dfxtp_4_45/a_1034_424#
+ sky130_fd_sc_hs__dfxtp_4
Xsky130_fd_sc_hs__a22o_1_60 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__a22o_1_61/X sky130_fd_sc_hs__nand2_1_39/B
+ sky130_fd_sc_hs__and2b_2_1/X init_val[27] rst sky130_fd_sc_hs__a22o_1_61/a_222_392#
+ sky130_fd_sc_hs__a22o_1_61/a_230_79# sky130_fd_sc_hs__a22o_1_61/a_52_123# sky130_fd_sc_hs__a22o_1_61/a_132_392#
+ sky130_fd_sc_hs__a22o_1
Xsky130_fd_sc_hs__dfxtp_4_12 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_1_13/B sky130_fd_sc_hs__a22o_1_17/X
+ sky130_fd_sc_hs__dfxtp_4_9/CLK sky130_fd_sc_hs__dfxtp_4_13/a_1226_296# sky130_fd_sc_hs__dfxtp_4_13/a_735_102#
+ sky130_fd_sc_hs__dfxtp_4_13/a_1141_508# sky130_fd_sc_hs__dfxtp_4_13/a_206_368# sky130_fd_sc_hs__dfxtp_4_13/a_437_503#
+ sky130_fd_sc_hs__dfxtp_4_13/a_27_74# sky130_fd_sc_hs__dfxtp_4_13/a_651_503# sky130_fd_sc_hs__dfxtp_4_13/a_696_458#
+ sky130_fd_sc_hs__dfxtp_4_13/a_544_485# sky130_fd_sc_hs__dfxtp_4_13/a_1178_124# sky130_fd_sc_hs__dfxtp_4_13/a_1034_424#
+ sky130_fd_sc_hs__dfxtp_4
Xsky130_fd_sc_hs__dfxtp_4_23 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_1_5/B sky130_fd_sc_hs__a22o_1_25/X
+ sky130_fd_sc_hs__dfxtp_4_9/CLK sky130_fd_sc_hs__dfxtp_4_23/a_1226_296# sky130_fd_sc_hs__dfxtp_4_23/a_735_102#
+ sky130_fd_sc_hs__dfxtp_4_23/a_1141_508# sky130_fd_sc_hs__dfxtp_4_23/a_206_368# sky130_fd_sc_hs__dfxtp_4_23/a_437_503#
+ sky130_fd_sc_hs__dfxtp_4_23/a_27_74# sky130_fd_sc_hs__dfxtp_4_23/a_651_503# sky130_fd_sc_hs__dfxtp_4_23/a_696_458#
+ sky130_fd_sc_hs__dfxtp_4_23/a_544_485# sky130_fd_sc_hs__dfxtp_4_23/a_1178_124# sky130_fd_sc_hs__dfxtp_4_23/a_1034_424#
+ sky130_fd_sc_hs__dfxtp_4
Xsky130_fd_sc_hs__dfxtp_4_34 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_1_43/B sky130_fd_sc_hs__a22o_1_31/X
+ sky130_fd_sc_hs__dfxtp_4_9/CLK sky130_fd_sc_hs__dfxtp_4_35/a_1226_296# sky130_fd_sc_hs__dfxtp_4_35/a_735_102#
+ sky130_fd_sc_hs__dfxtp_4_35/a_1141_508# sky130_fd_sc_hs__dfxtp_4_35/a_206_368# sky130_fd_sc_hs__dfxtp_4_35/a_437_503#
+ sky130_fd_sc_hs__dfxtp_4_35/a_27_74# sky130_fd_sc_hs__dfxtp_4_35/a_651_503# sky130_fd_sc_hs__dfxtp_4_35/a_696_458#
+ sky130_fd_sc_hs__dfxtp_4_35/a_544_485# sky130_fd_sc_hs__dfxtp_4_35/a_1178_124# sky130_fd_sc_hs__dfxtp_4_35/a_1034_424#
+ sky130_fd_sc_hs__dfxtp_4
Xsky130_fd_sc_hs__dfxtp_4_67 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_2_3/B sky130_fd_sc_hs__a22o_1_57/X
+ sky130_fd_sc_hs__dfxtp_4_9/CLK sky130_fd_sc_hs__dfxtp_4_67/a_1226_296# sky130_fd_sc_hs__dfxtp_4_67/a_735_102#
+ sky130_fd_sc_hs__dfxtp_4_67/a_1141_508# sky130_fd_sc_hs__dfxtp_4_67/a_206_368# sky130_fd_sc_hs__dfxtp_4_67/a_437_503#
+ sky130_fd_sc_hs__dfxtp_4_67/a_27_74# sky130_fd_sc_hs__dfxtp_4_67/a_651_503# sky130_fd_sc_hs__dfxtp_4_67/a_696_458#
+ sky130_fd_sc_hs__dfxtp_4_67/a_544_485# sky130_fd_sc_hs__dfxtp_4_67/a_1178_124# sky130_fd_sc_hs__dfxtp_4_67/a_1034_424#
+ sky130_fd_sc_hs__dfxtp_4
Xsky130_fd_sc_hs__dfxtp_4_56 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nor2b_1_4/A sky130_fd_sc_hs__nor2b_1_5/Y
+ sky130_fd_sc_hs__dfxtp_4_9/CLK sky130_fd_sc_hs__dfxtp_4_57/a_1226_296# sky130_fd_sc_hs__dfxtp_4_57/a_735_102#
+ sky130_fd_sc_hs__dfxtp_4_57/a_1141_508# sky130_fd_sc_hs__dfxtp_4_57/a_206_368# sky130_fd_sc_hs__dfxtp_4_57/a_437_503#
+ sky130_fd_sc_hs__dfxtp_4_57/a_27_74# sky130_fd_sc_hs__dfxtp_4_57/a_651_503# sky130_fd_sc_hs__dfxtp_4_57/a_696_458#
+ sky130_fd_sc_hs__dfxtp_4_57/a_544_485# sky130_fd_sc_hs__dfxtp_4_57/a_1178_124# sky130_fd_sc_hs__dfxtp_4_57/a_1034_424#
+ sky130_fd_sc_hs__dfxtp_4
Xsky130_fd_sc_hs__dfxtp_4_45 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_1_45/B sky130_fd_sc_hs__a22o_1_45/X
+ sky130_fd_sc_hs__dfxtp_4_9/CLK sky130_fd_sc_hs__dfxtp_4_45/a_1226_296# sky130_fd_sc_hs__dfxtp_4_45/a_735_102#
+ sky130_fd_sc_hs__dfxtp_4_45/a_1141_508# sky130_fd_sc_hs__dfxtp_4_45/a_206_368# sky130_fd_sc_hs__dfxtp_4_45/a_437_503#
+ sky130_fd_sc_hs__dfxtp_4_45/a_27_74# sky130_fd_sc_hs__dfxtp_4_45/a_651_503# sky130_fd_sc_hs__dfxtp_4_45/a_696_458#
+ sky130_fd_sc_hs__dfxtp_4_45/a_544_485# sky130_fd_sc_hs__dfxtp_4_45/a_1178_124# sky130_fd_sc_hs__dfxtp_4_45/a_1034_424#
+ sky130_fd_sc_hs__dfxtp_4
Xsky130_fd_sc_hs__a22o_1_61 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__a22o_1_61/X sky130_fd_sc_hs__nand2_1_39/B
+ sky130_fd_sc_hs__and2b_2_1/X init_val[27] rst sky130_fd_sc_hs__a22o_1_61/a_222_392#
+ sky130_fd_sc_hs__a22o_1_61/a_230_79# sky130_fd_sc_hs__a22o_1_61/a_52_123# sky130_fd_sc_hs__a22o_1_61/a_132_392#
+ sky130_fd_sc_hs__a22o_1
Xsky130_fd_sc_hs__a22o_1_50 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__a22o_1_51/X sky130_fd_sc_hs__nand2_1_57/B
+ sky130_fd_sc_hs__and2b_2_1/X init_val[31] rst sky130_fd_sc_hs__a22o_1_51/a_222_392#
+ sky130_fd_sc_hs__a22o_1_51/a_230_79# sky130_fd_sc_hs__a22o_1_51/a_52_123# sky130_fd_sc_hs__a22o_1_51/a_132_392#
+ sky130_fd_sc_hs__a22o_1
Xsky130_fd_sc_hs__nand2_1_50 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_1_51/B sky130_fd_sc_hs__xnor2_1_59/B
+ eqn[22] sky130_fd_sc_hs__nand2_1_51/a_117_74# sky130_fd_sc_hs__nand2_1
Xsky130_fd_sc_hs__dfxtp_4_13 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_1_13/B sky130_fd_sc_hs__a22o_1_17/X
+ sky130_fd_sc_hs__dfxtp_4_9/CLK sky130_fd_sc_hs__dfxtp_4_13/a_1226_296# sky130_fd_sc_hs__dfxtp_4_13/a_735_102#
+ sky130_fd_sc_hs__dfxtp_4_13/a_1141_508# sky130_fd_sc_hs__dfxtp_4_13/a_206_368# sky130_fd_sc_hs__dfxtp_4_13/a_437_503#
+ sky130_fd_sc_hs__dfxtp_4_13/a_27_74# sky130_fd_sc_hs__dfxtp_4_13/a_651_503# sky130_fd_sc_hs__dfxtp_4_13/a_696_458#
+ sky130_fd_sc_hs__dfxtp_4_13/a_544_485# sky130_fd_sc_hs__dfxtp_4_13/a_1178_124# sky130_fd_sc_hs__dfxtp_4_13/a_1034_424#
+ sky130_fd_sc_hs__dfxtp_4
Xsky130_fd_sc_hs__dfxtp_4_24 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_1_25/B sky130_fd_sc_hs__a22o_1_19/X
+ sky130_fd_sc_hs__dfxtp_4_9/CLK sky130_fd_sc_hs__dfxtp_4_25/a_1226_296# sky130_fd_sc_hs__dfxtp_4_25/a_735_102#
+ sky130_fd_sc_hs__dfxtp_4_25/a_1141_508# sky130_fd_sc_hs__dfxtp_4_25/a_206_368# sky130_fd_sc_hs__dfxtp_4_25/a_437_503#
+ sky130_fd_sc_hs__dfxtp_4_25/a_27_74# sky130_fd_sc_hs__dfxtp_4_25/a_651_503# sky130_fd_sc_hs__dfxtp_4_25/a_696_458#
+ sky130_fd_sc_hs__dfxtp_4_25/a_544_485# sky130_fd_sc_hs__dfxtp_4_25/a_1178_124# sky130_fd_sc_hs__dfxtp_4_25/a_1034_424#
+ sky130_fd_sc_hs__dfxtp_4
Xsky130_fd_sc_hs__dfxtp_4_35 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_1_43/B sky130_fd_sc_hs__a22o_1_31/X
+ sky130_fd_sc_hs__dfxtp_4_9/CLK sky130_fd_sc_hs__dfxtp_4_35/a_1226_296# sky130_fd_sc_hs__dfxtp_4_35/a_735_102#
+ sky130_fd_sc_hs__dfxtp_4_35/a_1141_508# sky130_fd_sc_hs__dfxtp_4_35/a_206_368# sky130_fd_sc_hs__dfxtp_4_35/a_437_503#
+ sky130_fd_sc_hs__dfxtp_4_35/a_27_74# sky130_fd_sc_hs__dfxtp_4_35/a_651_503# sky130_fd_sc_hs__dfxtp_4_35/a_696_458#
+ sky130_fd_sc_hs__dfxtp_4_35/a_544_485# sky130_fd_sc_hs__dfxtp_4_35/a_1178_124# sky130_fd_sc_hs__dfxtp_4_35/a_1034_424#
+ sky130_fd_sc_hs__dfxtp_4
Xsky130_fd_sc_hs__dfxtp_4_68 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_1_49/B sky130_fd_sc_hs__a22o_1_63/X
+ sky130_fd_sc_hs__dfxtp_4_9/CLK sky130_fd_sc_hs__dfxtp_4_69/a_1226_296# sky130_fd_sc_hs__dfxtp_4_69/a_735_102#
+ sky130_fd_sc_hs__dfxtp_4_69/a_1141_508# sky130_fd_sc_hs__dfxtp_4_69/a_206_368# sky130_fd_sc_hs__dfxtp_4_69/a_437_503#
+ sky130_fd_sc_hs__dfxtp_4_69/a_27_74# sky130_fd_sc_hs__dfxtp_4_69/a_651_503# sky130_fd_sc_hs__dfxtp_4_69/a_696_458#
+ sky130_fd_sc_hs__dfxtp_4_69/a_544_485# sky130_fd_sc_hs__dfxtp_4_69/a_1178_124# sky130_fd_sc_hs__dfxtp_4_69/a_1034_424#
+ sky130_fd_sc_hs__dfxtp_4
Xsky130_fd_sc_hs__dfxtp_4_57 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nor2b_1_4/A sky130_fd_sc_hs__nor2b_1_5/Y
+ sky130_fd_sc_hs__dfxtp_4_9/CLK sky130_fd_sc_hs__dfxtp_4_57/a_1226_296# sky130_fd_sc_hs__dfxtp_4_57/a_735_102#
+ sky130_fd_sc_hs__dfxtp_4_57/a_1141_508# sky130_fd_sc_hs__dfxtp_4_57/a_206_368# sky130_fd_sc_hs__dfxtp_4_57/a_437_503#
+ sky130_fd_sc_hs__dfxtp_4_57/a_27_74# sky130_fd_sc_hs__dfxtp_4_57/a_651_503# sky130_fd_sc_hs__dfxtp_4_57/a_696_458#
+ sky130_fd_sc_hs__dfxtp_4_57/a_544_485# sky130_fd_sc_hs__dfxtp_4_57/a_1178_124# sky130_fd_sc_hs__dfxtp_4_57/a_1034_424#
+ sky130_fd_sc_hs__dfxtp_4
Xsky130_fd_sc_hs__dfxtp_4_46 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_2_5/B sky130_fd_sc_hs__a22o_1_51/X
+ sky130_fd_sc_hs__dfxtp_4_9/CLK sky130_fd_sc_hs__dfxtp_4_47/a_1226_296# sky130_fd_sc_hs__dfxtp_4_47/a_735_102#
+ sky130_fd_sc_hs__dfxtp_4_47/a_1141_508# sky130_fd_sc_hs__dfxtp_4_47/a_206_368# sky130_fd_sc_hs__dfxtp_4_47/a_437_503#
+ sky130_fd_sc_hs__dfxtp_4_47/a_27_74# sky130_fd_sc_hs__dfxtp_4_47/a_651_503# sky130_fd_sc_hs__dfxtp_4_47/a_696_458#
+ sky130_fd_sc_hs__dfxtp_4_47/a_544_485# sky130_fd_sc_hs__dfxtp_4_47/a_1178_124# sky130_fd_sc_hs__dfxtp_4_47/a_1034_424#
+ sky130_fd_sc_hs__dfxtp_4
Xsky130_fd_sc_hs__xnor2_1_0 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__xnor2_1_1/A sky130_fd_sc_hs__xnor2_1_7/A
+ sky130_fd_sc_hs__xnor2_1_1/B sky130_fd_sc_hs__xnor2_1_1/a_376_368# sky130_fd_sc_hs__xnor2_1_1/a_112_119#
+ sky130_fd_sc_hs__xnor2_1_1/a_138_385# sky130_fd_sc_hs__xnor2_1_1/a_293_74# sky130_fd_sc_hs__xnor2_1
Xsky130_fd_sc_hs__a22o_1_62 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__a22o_1_63/X sky130_fd_sc_hs__nand2_1_53/B
+ sky130_fd_sc_hs__and2b_2_1/X init_val[28] rst sky130_fd_sc_hs__a22o_1_63/a_222_392#
+ sky130_fd_sc_hs__a22o_1_63/a_230_79# sky130_fd_sc_hs__a22o_1_63/a_52_123# sky130_fd_sc_hs__a22o_1_63/a_132_392#
+ sky130_fd_sc_hs__a22o_1
Xsky130_fd_sc_hs__a22o_1_51 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__a22o_1_51/X sky130_fd_sc_hs__nand2_1_57/B
+ sky130_fd_sc_hs__and2b_2_1/X init_val[31] rst sky130_fd_sc_hs__a22o_1_51/a_222_392#
+ sky130_fd_sc_hs__a22o_1_51/a_230_79# sky130_fd_sc_hs__a22o_1_51/a_52_123# sky130_fd_sc_hs__a22o_1_51/a_132_392#
+ sky130_fd_sc_hs__a22o_1
Xsky130_fd_sc_hs__a22o_1_40 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__a22o_1_41/X sky130_fd_sc_hs__nand2_1_43/B
+ sky130_fd_sc_hs__and2b_2_1/X init_val[19] rst sky130_fd_sc_hs__a22o_1_41/a_222_392#
+ sky130_fd_sc_hs__a22o_1_41/a_230_79# sky130_fd_sc_hs__a22o_1_41/a_52_123# sky130_fd_sc_hs__a22o_1_41/a_132_392#
+ sky130_fd_sc_hs__a22o_1
Xsky130_fd_sc_hs__nand2_1_40 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_1_41/B sky130_fd_sc_hs__xnor2_1_53/A
+ eqn[0] sky130_fd_sc_hs__nand2_1_41/a_117_74# sky130_fd_sc_hs__nand2_1
Xsky130_fd_sc_hs__nand2_1_51 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_1_51/B sky130_fd_sc_hs__xnor2_1_59/B
+ eqn[22] sky130_fd_sc_hs__nand2_1_51/a_117_74# sky130_fd_sc_hs__nand2_1
Xsky130_fd_sc_hs__dfxtp_4_14 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_1_21/B sky130_fd_sc_hs__a22o_1_15/X
+ sky130_fd_sc_hs__dfxtp_4_9/CLK sky130_fd_sc_hs__dfxtp_4_15/a_1226_296# sky130_fd_sc_hs__dfxtp_4_15/a_735_102#
+ sky130_fd_sc_hs__dfxtp_4_15/a_1141_508# sky130_fd_sc_hs__dfxtp_4_15/a_206_368# sky130_fd_sc_hs__dfxtp_4_15/a_437_503#
+ sky130_fd_sc_hs__dfxtp_4_15/a_27_74# sky130_fd_sc_hs__dfxtp_4_15/a_651_503# sky130_fd_sc_hs__dfxtp_4_15/a_696_458#
+ sky130_fd_sc_hs__dfxtp_4_15/a_544_485# sky130_fd_sc_hs__dfxtp_4_15/a_1178_124# sky130_fd_sc_hs__dfxtp_4_15/a_1034_424#
+ sky130_fd_sc_hs__dfxtp_4
Xsky130_fd_sc_hs__dfxtp_4_25 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_1_25/B sky130_fd_sc_hs__a22o_1_19/X
+ sky130_fd_sc_hs__dfxtp_4_9/CLK sky130_fd_sc_hs__dfxtp_4_25/a_1226_296# sky130_fd_sc_hs__dfxtp_4_25/a_735_102#
+ sky130_fd_sc_hs__dfxtp_4_25/a_1141_508# sky130_fd_sc_hs__dfxtp_4_25/a_206_368# sky130_fd_sc_hs__dfxtp_4_25/a_437_503#
+ sky130_fd_sc_hs__dfxtp_4_25/a_27_74# sky130_fd_sc_hs__dfxtp_4_25/a_651_503# sky130_fd_sc_hs__dfxtp_4_25/a_696_458#
+ sky130_fd_sc_hs__dfxtp_4_25/a_544_485# sky130_fd_sc_hs__dfxtp_4_25/a_1178_124# sky130_fd_sc_hs__dfxtp_4_25/a_1034_424#
+ sky130_fd_sc_hs__dfxtp_4
Xsky130_fd_sc_hs__dfxtp_4_36 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_1_33/B sky130_fd_sc_hs__a22o_1_43/X
+ sky130_fd_sc_hs__dfxtp_4_9/CLK sky130_fd_sc_hs__dfxtp_4_37/a_1226_296# sky130_fd_sc_hs__dfxtp_4_37/a_735_102#
+ sky130_fd_sc_hs__dfxtp_4_37/a_1141_508# sky130_fd_sc_hs__dfxtp_4_37/a_206_368# sky130_fd_sc_hs__dfxtp_4_37/a_437_503#
+ sky130_fd_sc_hs__dfxtp_4_37/a_27_74# sky130_fd_sc_hs__dfxtp_4_37/a_651_503# sky130_fd_sc_hs__dfxtp_4_37/a_696_458#
+ sky130_fd_sc_hs__dfxtp_4_37/a_544_485# sky130_fd_sc_hs__dfxtp_4_37/a_1178_124# sky130_fd_sc_hs__dfxtp_4_37/a_1034_424#
+ sky130_fd_sc_hs__dfxtp_4
Xsky130_fd_sc_hs__dfxtp_4_69 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_1_49/B sky130_fd_sc_hs__a22o_1_63/X
+ sky130_fd_sc_hs__dfxtp_4_9/CLK sky130_fd_sc_hs__dfxtp_4_69/a_1226_296# sky130_fd_sc_hs__dfxtp_4_69/a_735_102#
+ sky130_fd_sc_hs__dfxtp_4_69/a_1141_508# sky130_fd_sc_hs__dfxtp_4_69/a_206_368# sky130_fd_sc_hs__dfxtp_4_69/a_437_503#
+ sky130_fd_sc_hs__dfxtp_4_69/a_27_74# sky130_fd_sc_hs__dfxtp_4_69/a_651_503# sky130_fd_sc_hs__dfxtp_4_69/a_696_458#
+ sky130_fd_sc_hs__dfxtp_4_69/a_544_485# sky130_fd_sc_hs__dfxtp_4_69/a_1178_124# sky130_fd_sc_hs__dfxtp_4_69/a_1034_424#
+ sky130_fd_sc_hs__dfxtp_4
Xsky130_fd_sc_hs__dfxtp_4_58 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_1_35/B sky130_fd_sc_hs__a22o_1_55/X
+ sky130_fd_sc_hs__dfxtp_4_9/CLK sky130_fd_sc_hs__dfxtp_4_59/a_1226_296# sky130_fd_sc_hs__dfxtp_4_59/a_735_102#
+ sky130_fd_sc_hs__dfxtp_4_59/a_1141_508# sky130_fd_sc_hs__dfxtp_4_59/a_206_368# sky130_fd_sc_hs__dfxtp_4_59/a_437_503#
+ sky130_fd_sc_hs__dfxtp_4_59/a_27_74# sky130_fd_sc_hs__dfxtp_4_59/a_651_503# sky130_fd_sc_hs__dfxtp_4_59/a_696_458#
+ sky130_fd_sc_hs__dfxtp_4_59/a_544_485# sky130_fd_sc_hs__dfxtp_4_59/a_1178_124# sky130_fd_sc_hs__dfxtp_4_59/a_1034_424#
+ sky130_fd_sc_hs__dfxtp_4
Xsky130_fd_sc_hs__dfxtp_4_47 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_2_5/B sky130_fd_sc_hs__a22o_1_51/X
+ sky130_fd_sc_hs__dfxtp_4_9/CLK sky130_fd_sc_hs__dfxtp_4_47/a_1226_296# sky130_fd_sc_hs__dfxtp_4_47/a_735_102#
+ sky130_fd_sc_hs__dfxtp_4_47/a_1141_508# sky130_fd_sc_hs__dfxtp_4_47/a_206_368# sky130_fd_sc_hs__dfxtp_4_47/a_437_503#
+ sky130_fd_sc_hs__dfxtp_4_47/a_27_74# sky130_fd_sc_hs__dfxtp_4_47/a_651_503# sky130_fd_sc_hs__dfxtp_4_47/a_696_458#
+ sky130_fd_sc_hs__dfxtp_4_47/a_544_485# sky130_fd_sc_hs__dfxtp_4_47/a_1178_124# sky130_fd_sc_hs__dfxtp_4_47/a_1034_424#
+ sky130_fd_sc_hs__dfxtp_4
Xsky130_fd_sc_hs__xnor2_1_1 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__xnor2_1_1/A sky130_fd_sc_hs__xnor2_1_7/A
+ sky130_fd_sc_hs__xnor2_1_1/B sky130_fd_sc_hs__xnor2_1_1/a_376_368# sky130_fd_sc_hs__xnor2_1_1/a_112_119#
+ sky130_fd_sc_hs__xnor2_1_1/a_138_385# sky130_fd_sc_hs__xnor2_1_1/a_293_74# sky130_fd_sc_hs__xnor2_1
Xsky130_fd_sc_hs__or2_1_0 DVSS DVDD DVDD DVSS cke rst sky130_fd_sc_hs__or2_1_1/X sky130_fd_sc_hs__or2_1_1/a_152_368#
+ sky130_fd_sc_hs__or2_1_1/a_63_368# sky130_fd_sc_hs__or2_1
Xsky130_fd_sc_hs__a22o_1_30 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__a22o_1_31/X sky130_fd_sc_hs__nand2_1_31/B
+ sky130_fd_sc_hs__and2b_2_1/X init_val[18] rst sky130_fd_sc_hs__a22o_1_31/a_222_392#
+ sky130_fd_sc_hs__a22o_1_31/a_230_79# sky130_fd_sc_hs__a22o_1_31/a_52_123# sky130_fd_sc_hs__a22o_1_31/a_132_392#
+ sky130_fd_sc_hs__a22o_1
Xsky130_fd_sc_hs__a22o_1_52 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__a22o_1_53/X sky130_fd_sc_hs__nand2_1_35/B
+ sky130_fd_sc_hs__and2b_2_1/X init_val[24] rst sky130_fd_sc_hs__a22o_1_53/a_222_392#
+ sky130_fd_sc_hs__a22o_1_53/a_230_79# sky130_fd_sc_hs__a22o_1_53/a_52_123# sky130_fd_sc_hs__a22o_1_53/a_132_392#
+ sky130_fd_sc_hs__a22o_1
Xsky130_fd_sc_hs__a22o_1_63 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__a22o_1_63/X sky130_fd_sc_hs__nand2_1_53/B
+ sky130_fd_sc_hs__and2b_2_1/X init_val[28] rst sky130_fd_sc_hs__a22o_1_63/a_222_392#
+ sky130_fd_sc_hs__a22o_1_63/a_230_79# sky130_fd_sc_hs__a22o_1_63/a_52_123# sky130_fd_sc_hs__a22o_1_63/a_132_392#
+ sky130_fd_sc_hs__a22o_1
Xsky130_fd_sc_hs__a22o_1_41 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__a22o_1_41/X sky130_fd_sc_hs__nand2_1_43/B
+ sky130_fd_sc_hs__and2b_2_1/X init_val[19] rst sky130_fd_sc_hs__a22o_1_41/a_222_392#
+ sky130_fd_sc_hs__a22o_1_41/a_230_79# sky130_fd_sc_hs__a22o_1_41/a_52_123# sky130_fd_sc_hs__a22o_1_41/a_132_392#
+ sky130_fd_sc_hs__a22o_1
Xsky130_fd_sc_hs__nand2_1_30 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_1_31/B sky130_fd_sc_hs__xnor2_1_21/A
+ eqn[17] sky130_fd_sc_hs__nand2_1_31/a_117_74# sky130_fd_sc_hs__nand2_1
Xsky130_fd_sc_hs__nand2_1_41 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_1_41/B sky130_fd_sc_hs__xnor2_1_53/A
+ eqn[0] sky130_fd_sc_hs__nand2_1_41/a_117_74# sky130_fd_sc_hs__nand2_1
Xsky130_fd_sc_hs__nand2_1_52 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_1_53/B sky130_fd_sc_hs__xnor2_1_61/A
+ eqn[27] sky130_fd_sc_hs__nand2_1_53/a_117_74# sky130_fd_sc_hs__nand2_1
Xsky130_fd_sc_hs__dfxtp_4_15 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_1_21/B sky130_fd_sc_hs__a22o_1_15/X
+ sky130_fd_sc_hs__dfxtp_4_9/CLK sky130_fd_sc_hs__dfxtp_4_15/a_1226_296# sky130_fd_sc_hs__dfxtp_4_15/a_735_102#
+ sky130_fd_sc_hs__dfxtp_4_15/a_1141_508# sky130_fd_sc_hs__dfxtp_4_15/a_206_368# sky130_fd_sc_hs__dfxtp_4_15/a_437_503#
+ sky130_fd_sc_hs__dfxtp_4_15/a_27_74# sky130_fd_sc_hs__dfxtp_4_15/a_651_503# sky130_fd_sc_hs__dfxtp_4_15/a_696_458#
+ sky130_fd_sc_hs__dfxtp_4_15/a_544_485# sky130_fd_sc_hs__dfxtp_4_15/a_1178_124# sky130_fd_sc_hs__dfxtp_4_15/a_1034_424#
+ sky130_fd_sc_hs__dfxtp_4
Xsky130_fd_sc_hs__dfxtp_4_26 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_1_9/B sky130_fd_sc_hs__a22o_1_27/X
+ sky130_fd_sc_hs__dfxtp_4_9/CLK sky130_fd_sc_hs__dfxtp_4_27/a_1226_296# sky130_fd_sc_hs__dfxtp_4_27/a_735_102#
+ sky130_fd_sc_hs__dfxtp_4_27/a_1141_508# sky130_fd_sc_hs__dfxtp_4_27/a_206_368# sky130_fd_sc_hs__dfxtp_4_27/a_437_503#
+ sky130_fd_sc_hs__dfxtp_4_27/a_27_74# sky130_fd_sc_hs__dfxtp_4_27/a_651_503# sky130_fd_sc_hs__dfxtp_4_27/a_696_458#
+ sky130_fd_sc_hs__dfxtp_4_27/a_544_485# sky130_fd_sc_hs__dfxtp_4_27/a_1178_124# sky130_fd_sc_hs__dfxtp_4_27/a_1034_424#
+ sky130_fd_sc_hs__dfxtp_4
Xsky130_fd_sc_hs__dfxtp_4_37 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_1_33/B sky130_fd_sc_hs__a22o_1_43/X
+ sky130_fd_sc_hs__dfxtp_4_9/CLK sky130_fd_sc_hs__dfxtp_4_37/a_1226_296# sky130_fd_sc_hs__dfxtp_4_37/a_735_102#
+ sky130_fd_sc_hs__dfxtp_4_37/a_1141_508# sky130_fd_sc_hs__dfxtp_4_37/a_206_368# sky130_fd_sc_hs__dfxtp_4_37/a_437_503#
+ sky130_fd_sc_hs__dfxtp_4_37/a_27_74# sky130_fd_sc_hs__dfxtp_4_37/a_651_503# sky130_fd_sc_hs__dfxtp_4_37/a_696_458#
+ sky130_fd_sc_hs__dfxtp_4_37/a_544_485# sky130_fd_sc_hs__dfxtp_4_37/a_1178_124# sky130_fd_sc_hs__dfxtp_4_37/a_1034_424#
+ sky130_fd_sc_hs__dfxtp_4
Xsky130_fd_sc_hs__dfxtp_4_59 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_1_35/B sky130_fd_sc_hs__a22o_1_55/X
+ sky130_fd_sc_hs__dfxtp_4_9/CLK sky130_fd_sc_hs__dfxtp_4_59/a_1226_296# sky130_fd_sc_hs__dfxtp_4_59/a_735_102#
+ sky130_fd_sc_hs__dfxtp_4_59/a_1141_508# sky130_fd_sc_hs__dfxtp_4_59/a_206_368# sky130_fd_sc_hs__dfxtp_4_59/a_437_503#
+ sky130_fd_sc_hs__dfxtp_4_59/a_27_74# sky130_fd_sc_hs__dfxtp_4_59/a_651_503# sky130_fd_sc_hs__dfxtp_4_59/a_696_458#
+ sky130_fd_sc_hs__dfxtp_4_59/a_544_485# sky130_fd_sc_hs__dfxtp_4_59/a_1178_124# sky130_fd_sc_hs__dfxtp_4_59/a_1034_424#
+ sky130_fd_sc_hs__dfxtp_4
Xsky130_fd_sc_hs__dfxtp_4_48 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_1_57/B sky130_fd_sc_hs__a22o_1_39/X
+ sky130_fd_sc_hs__dfxtp_4_9/CLK sky130_fd_sc_hs__dfxtp_4_49/a_1226_296# sky130_fd_sc_hs__dfxtp_4_49/a_735_102#
+ sky130_fd_sc_hs__dfxtp_4_49/a_1141_508# sky130_fd_sc_hs__dfxtp_4_49/a_206_368# sky130_fd_sc_hs__dfxtp_4_49/a_437_503#
+ sky130_fd_sc_hs__dfxtp_4_49/a_27_74# sky130_fd_sc_hs__dfxtp_4_49/a_651_503# sky130_fd_sc_hs__dfxtp_4_49/a_696_458#
+ sky130_fd_sc_hs__dfxtp_4_49/a_544_485# sky130_fd_sc_hs__dfxtp_4_49/a_1178_124# sky130_fd_sc_hs__dfxtp_4_49/a_1034_424#
+ sky130_fd_sc_hs__dfxtp_4
Xsky130_fd_sc_hs__nand2_2_0 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__xnor2_1_3/A sky130_fd_sc_hs__nand2_2_1/B
+ eqn[11] sky130_fd_sc_hs__nand2_2_1/a_27_74# sky130_fd_sc_hs__nand2_2
Xsky130_fd_sc_hs__xnor2_1_2 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__xnor2_1_3/A sky130_fd_sc_hs__xnor2_1_5/A
+ sky130_fd_sc_hs__xnor2_1_3/B sky130_fd_sc_hs__xnor2_1_3/a_376_368# sky130_fd_sc_hs__xnor2_1_3/a_112_119#
+ sky130_fd_sc_hs__xnor2_1_3/a_138_385# sky130_fd_sc_hs__xnor2_1_3/a_293_74# sky130_fd_sc_hs__xnor2_1
Xsky130_fd_sc_hs__or2_1_1 DVSS DVDD DVDD DVSS cke rst sky130_fd_sc_hs__or2_1_1/X sky130_fd_sc_hs__or2_1_1/a_152_368#
+ sky130_fd_sc_hs__or2_1_1/a_63_368# sky130_fd_sc_hs__or2_1
Xsky130_fd_sc_hs__a22o_1_20 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__a22o_1_21/X sky130_fd_sc_hs__nand2_1_19/B
+ sky130_fd_sc_hs__and2b_2_1/X init_val[17] rst sky130_fd_sc_hs__a22o_1_21/a_222_392#
+ sky130_fd_sc_hs__a22o_1_21/a_230_79# sky130_fd_sc_hs__a22o_1_21/a_52_123# sky130_fd_sc_hs__a22o_1_21/a_132_392#
+ sky130_fd_sc_hs__a22o_1
Xsky130_fd_sc_hs__a22o_1_31 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__a22o_1_31/X sky130_fd_sc_hs__nand2_1_31/B
+ sky130_fd_sc_hs__and2b_2_1/X init_val[18] rst sky130_fd_sc_hs__a22o_1_31/a_222_392#
+ sky130_fd_sc_hs__a22o_1_31/a_230_79# sky130_fd_sc_hs__a22o_1_31/a_52_123# sky130_fd_sc_hs__a22o_1_31/a_132_392#
+ sky130_fd_sc_hs__a22o_1
Xsky130_fd_sc_hs__a22o_1_53 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__a22o_1_53/X sky130_fd_sc_hs__nand2_1_35/B
+ sky130_fd_sc_hs__and2b_2_1/X init_val[24] rst sky130_fd_sc_hs__a22o_1_53/a_222_392#
+ sky130_fd_sc_hs__a22o_1_53/a_230_79# sky130_fd_sc_hs__a22o_1_53/a_52_123# sky130_fd_sc_hs__a22o_1_53/a_132_392#
+ sky130_fd_sc_hs__a22o_1
Xsky130_fd_sc_hs__a22o_1_42 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__a22o_1_43/X sky130_fd_sc_hs__nand2_1_47/B
+ sky130_fd_sc_hs__and2b_2_1/X init_val[20] rst sky130_fd_sc_hs__a22o_1_43/a_222_392#
+ sky130_fd_sc_hs__a22o_1_43/a_230_79# sky130_fd_sc_hs__a22o_1_43/a_52_123# sky130_fd_sc_hs__a22o_1_43/a_132_392#
+ sky130_fd_sc_hs__a22o_1
Xsky130_fd_sc_hs__nand2_1_20 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_1_21/B sky130_fd_sc_hs__xnor2_1_13/A
+ eqn[7] sky130_fd_sc_hs__nand2_1_21/a_117_74# sky130_fd_sc_hs__nand2_1
Xsky130_fd_sc_hs__nand2_1_31 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_1_31/B sky130_fd_sc_hs__xnor2_1_21/A
+ eqn[17] sky130_fd_sc_hs__nand2_1_31/a_117_74# sky130_fd_sc_hs__nand2_1
Xsky130_fd_sc_hs__nand2_1_42 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_1_43/B sky130_fd_sc_hs__xnor2_1_55/A
+ eqn[18] sky130_fd_sc_hs__nand2_1_43/a_117_74# sky130_fd_sc_hs__nand2_1
Xsky130_fd_sc_hs__nand2_1_53 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_1_53/B sky130_fd_sc_hs__xnor2_1_61/A
+ eqn[27] sky130_fd_sc_hs__nand2_1_53/a_117_74# sky130_fd_sc_hs__nand2_1
Xsky130_fd_sc_hs__dfxtp_4_16 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_1_19/B sky130_fd_sc_hs__a22o_1_13/X
+ sky130_fd_sc_hs__dfxtp_4_9/CLK sky130_fd_sc_hs__dfxtp_4_17/a_1226_296# sky130_fd_sc_hs__dfxtp_4_17/a_735_102#
+ sky130_fd_sc_hs__dfxtp_4_17/a_1141_508# sky130_fd_sc_hs__dfxtp_4_17/a_206_368# sky130_fd_sc_hs__dfxtp_4_17/a_437_503#
+ sky130_fd_sc_hs__dfxtp_4_17/a_27_74# sky130_fd_sc_hs__dfxtp_4_17/a_651_503# sky130_fd_sc_hs__dfxtp_4_17/a_696_458#
+ sky130_fd_sc_hs__dfxtp_4_17/a_544_485# sky130_fd_sc_hs__dfxtp_4_17/a_1178_124# sky130_fd_sc_hs__dfxtp_4_17/a_1034_424#
+ sky130_fd_sc_hs__dfxtp_4
Xsky130_fd_sc_hs__dfxtp_4_27 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_1_9/B sky130_fd_sc_hs__a22o_1_27/X
+ sky130_fd_sc_hs__dfxtp_4_9/CLK sky130_fd_sc_hs__dfxtp_4_27/a_1226_296# sky130_fd_sc_hs__dfxtp_4_27/a_735_102#
+ sky130_fd_sc_hs__dfxtp_4_27/a_1141_508# sky130_fd_sc_hs__dfxtp_4_27/a_206_368# sky130_fd_sc_hs__dfxtp_4_27/a_437_503#
+ sky130_fd_sc_hs__dfxtp_4_27/a_27_74# sky130_fd_sc_hs__dfxtp_4_27/a_651_503# sky130_fd_sc_hs__dfxtp_4_27/a_696_458#
+ sky130_fd_sc_hs__dfxtp_4_27/a_544_485# sky130_fd_sc_hs__dfxtp_4_27/a_1178_124# sky130_fd_sc_hs__dfxtp_4_27/a_1034_424#
+ sky130_fd_sc_hs__dfxtp_4
Xsky130_fd_sc_hs__dfxtp_4_38 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_1_27/B sky130_fd_sc_hs__a22o_1_35/X
+ sky130_fd_sc_hs__dfxtp_4_9/CLK sky130_fd_sc_hs__dfxtp_4_39/a_1226_296# sky130_fd_sc_hs__dfxtp_4_39/a_735_102#
+ sky130_fd_sc_hs__dfxtp_4_39/a_1141_508# sky130_fd_sc_hs__dfxtp_4_39/a_206_368# sky130_fd_sc_hs__dfxtp_4_39/a_437_503#
+ sky130_fd_sc_hs__dfxtp_4_39/a_27_74# sky130_fd_sc_hs__dfxtp_4_39/a_651_503# sky130_fd_sc_hs__dfxtp_4_39/a_696_458#
+ sky130_fd_sc_hs__dfxtp_4_39/a_544_485# sky130_fd_sc_hs__dfxtp_4_39/a_1178_124# sky130_fd_sc_hs__dfxtp_4_39/a_1034_424#
+ sky130_fd_sc_hs__dfxtp_4
Xsky130_fd_sc_hs__dfxtp_4_49 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_1_57/B sky130_fd_sc_hs__a22o_1_39/X
+ sky130_fd_sc_hs__dfxtp_4_9/CLK sky130_fd_sc_hs__dfxtp_4_49/a_1226_296# sky130_fd_sc_hs__dfxtp_4_49/a_735_102#
+ sky130_fd_sc_hs__dfxtp_4_49/a_1141_508# sky130_fd_sc_hs__dfxtp_4_49/a_206_368# sky130_fd_sc_hs__dfxtp_4_49/a_437_503#
+ sky130_fd_sc_hs__dfxtp_4_49/a_27_74# sky130_fd_sc_hs__dfxtp_4_49/a_651_503# sky130_fd_sc_hs__dfxtp_4_49/a_696_458#
+ sky130_fd_sc_hs__dfxtp_4_49/a_544_485# sky130_fd_sc_hs__dfxtp_4_49/a_1178_124# sky130_fd_sc_hs__dfxtp_4_49/a_1034_424#
+ sky130_fd_sc_hs__dfxtp_4
Xsky130_fd_sc_hs__nand2_2_1 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__xnor2_1_3/A sky130_fd_sc_hs__nand2_2_1/B
+ eqn[11] sky130_fd_sc_hs__nand2_2_1/a_27_74# sky130_fd_sc_hs__nand2_2
Xsky130_fd_sc_hs__xnor2_1_3 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__xnor2_1_3/A sky130_fd_sc_hs__xnor2_1_5/A
+ sky130_fd_sc_hs__xnor2_1_3/B sky130_fd_sc_hs__xnor2_1_3/a_376_368# sky130_fd_sc_hs__xnor2_1_3/a_112_119#
+ sky130_fd_sc_hs__xnor2_1_3/a_138_385# sky130_fd_sc_hs__xnor2_1_3/a_293_74# sky130_fd_sc_hs__xnor2_1
Xsky130_fd_sc_hs__a22o_1_10 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__dfxtp_4_8/D sky130_fd_sc_hs__nand2_1_21/B
+ sky130_fd_sc_hs__and2b_2_1/X init_val[8] rst sky130_fd_sc_hs__a22o_1_11/a_222_392#
+ sky130_fd_sc_hs__a22o_1_11/a_230_79# sky130_fd_sc_hs__a22o_1_11/a_52_123# sky130_fd_sc_hs__a22o_1_11/a_132_392#
+ sky130_fd_sc_hs__a22o_1
Xsky130_fd_sc_hs__a22o_1_21 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__a22o_1_21/X sky130_fd_sc_hs__nand2_1_19/B
+ sky130_fd_sc_hs__and2b_2_1/X init_val[17] rst sky130_fd_sc_hs__a22o_1_21/a_222_392#
+ sky130_fd_sc_hs__a22o_1_21/a_230_79# sky130_fd_sc_hs__a22o_1_21/a_52_123# sky130_fd_sc_hs__a22o_1_21/a_132_392#
+ sky130_fd_sc_hs__a22o_1
Xsky130_fd_sc_hs__a22o_1_32 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__a22o_1_33/X sky130_fd_sc_hs__nand2_1_45/B
+ sky130_fd_sc_hs__and2b_2_1/X init_val[2] rst sky130_fd_sc_hs__a22o_1_33/a_222_392#
+ sky130_fd_sc_hs__a22o_1_33/a_230_79# sky130_fd_sc_hs__a22o_1_33/a_52_123# sky130_fd_sc_hs__a22o_1_33/a_132_392#
+ sky130_fd_sc_hs__a22o_1
Xsky130_fd_sc_hs__a22o_1_54 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__a22o_1_55/X sky130_fd_sc_hs__nand2_1_51/B
+ sky130_fd_sc_hs__and2b_2_1/X init_val[23] rst sky130_fd_sc_hs__a22o_1_55/a_222_392#
+ sky130_fd_sc_hs__a22o_1_55/a_230_79# sky130_fd_sc_hs__a22o_1_55/a_52_123# sky130_fd_sc_hs__a22o_1_55/a_132_392#
+ sky130_fd_sc_hs__a22o_1
Xsky130_fd_sc_hs__a22o_1_43 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__a22o_1_43/X sky130_fd_sc_hs__nand2_1_47/B
+ sky130_fd_sc_hs__and2b_2_1/X init_val[20] rst sky130_fd_sc_hs__a22o_1_43/a_222_392#
+ sky130_fd_sc_hs__a22o_1_43/a_230_79# sky130_fd_sc_hs__a22o_1_43/a_52_123# sky130_fd_sc_hs__a22o_1_43/a_132_392#
+ sky130_fd_sc_hs__a22o_1
Xsky130_fd_sc_hs__nand2_1_10 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__dfxtp_4_7/Q sky130_fd_sc_hs__xnor2_1_35/B
+ eqn[10] sky130_fd_sc_hs__nand2_1_11/a_117_74# sky130_fd_sc_hs__nand2_1
Xsky130_fd_sc_hs__nand2_1_21 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_1_21/B sky130_fd_sc_hs__xnor2_1_13/A
+ eqn[7] sky130_fd_sc_hs__nand2_1_21/a_117_74# sky130_fd_sc_hs__nand2_1
Xsky130_fd_sc_hs__nand2_1_32 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_1_33/B sky130_fd_sc_hs__xnor2_1_21/B
+ eqn[20] sky130_fd_sc_hs__nand2_1_33/a_117_74# sky130_fd_sc_hs__nand2_1
Xsky130_fd_sc_hs__nand2_1_43 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_1_43/B sky130_fd_sc_hs__xnor2_1_55/A
+ eqn[18] sky130_fd_sc_hs__nand2_1_43/a_117_74# sky130_fd_sc_hs__nand2_1
Xsky130_fd_sc_hs__nand2_1_54 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_1_55/B sky130_fd_sc_hs__xnor2_1_31/B
+ eqn[29] sky130_fd_sc_hs__nand2_1_55/a_117_74# sky130_fd_sc_hs__nand2_1
Xsky130_fd_sc_hs__dfxtp_4_0 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__dfxtp_4_1/Q sky130_fd_sc_hs__a22o_1_1/X
+ sky130_fd_sc_hs__dfxtp_4_9/CLK sky130_fd_sc_hs__dfxtp_4_1/a_1226_296# sky130_fd_sc_hs__dfxtp_4_1/a_735_102#
+ sky130_fd_sc_hs__dfxtp_4_1/a_1141_508# sky130_fd_sc_hs__dfxtp_4_1/a_206_368# sky130_fd_sc_hs__dfxtp_4_1/a_437_503#
+ sky130_fd_sc_hs__dfxtp_4_1/a_27_74# sky130_fd_sc_hs__dfxtp_4_1/a_651_503# sky130_fd_sc_hs__dfxtp_4_1/a_696_458#
+ sky130_fd_sc_hs__dfxtp_4_1/a_544_485# sky130_fd_sc_hs__dfxtp_4_1/a_1178_124# sky130_fd_sc_hs__dfxtp_4_1/a_1034_424#
+ sky130_fd_sc_hs__dfxtp_4
Xsky130_fd_sc_hs__dfxtp_4_17 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_1_19/B sky130_fd_sc_hs__a22o_1_13/X
+ sky130_fd_sc_hs__dfxtp_4_9/CLK sky130_fd_sc_hs__dfxtp_4_17/a_1226_296# sky130_fd_sc_hs__dfxtp_4_17/a_735_102#
+ sky130_fd_sc_hs__dfxtp_4_17/a_1141_508# sky130_fd_sc_hs__dfxtp_4_17/a_206_368# sky130_fd_sc_hs__dfxtp_4_17/a_437_503#
+ sky130_fd_sc_hs__dfxtp_4_17/a_27_74# sky130_fd_sc_hs__dfxtp_4_17/a_651_503# sky130_fd_sc_hs__dfxtp_4_17/a_696_458#
+ sky130_fd_sc_hs__dfxtp_4_17/a_544_485# sky130_fd_sc_hs__dfxtp_4_17/a_1178_124# sky130_fd_sc_hs__dfxtp_4_17/a_1034_424#
+ sky130_fd_sc_hs__dfxtp_4
Xsky130_fd_sc_hs__dfxtp_4_28 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_1_17/B sky130_fd_sc_hs__a22o_1_29/X
+ sky130_fd_sc_hs__dfxtp_4_9/CLK sky130_fd_sc_hs__dfxtp_4_29/a_1226_296# sky130_fd_sc_hs__dfxtp_4_29/a_735_102#
+ sky130_fd_sc_hs__dfxtp_4_29/a_1141_508# sky130_fd_sc_hs__dfxtp_4_29/a_206_368# sky130_fd_sc_hs__dfxtp_4_29/a_437_503#
+ sky130_fd_sc_hs__dfxtp_4_29/a_27_74# sky130_fd_sc_hs__dfxtp_4_29/a_651_503# sky130_fd_sc_hs__dfxtp_4_29/a_696_458#
+ sky130_fd_sc_hs__dfxtp_4_29/a_544_485# sky130_fd_sc_hs__dfxtp_4_29/a_1178_124# sky130_fd_sc_hs__dfxtp_4_29/a_1034_424#
+ sky130_fd_sc_hs__dfxtp_4
Xsky130_fd_sc_hs__dfxtp_4_39 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_1_27/B sky130_fd_sc_hs__a22o_1_35/X
+ sky130_fd_sc_hs__dfxtp_4_9/CLK sky130_fd_sc_hs__dfxtp_4_39/a_1226_296# sky130_fd_sc_hs__dfxtp_4_39/a_735_102#
+ sky130_fd_sc_hs__dfxtp_4_39/a_1141_508# sky130_fd_sc_hs__dfxtp_4_39/a_206_368# sky130_fd_sc_hs__dfxtp_4_39/a_437_503#
+ sky130_fd_sc_hs__dfxtp_4_39/a_27_74# sky130_fd_sc_hs__dfxtp_4_39/a_651_503# sky130_fd_sc_hs__dfxtp_4_39/a_696_458#
+ sky130_fd_sc_hs__dfxtp_4_39/a_544_485# sky130_fd_sc_hs__dfxtp_4_39/a_1178_124# sky130_fd_sc_hs__dfxtp_4_39/a_1034_424#
+ sky130_fd_sc_hs__dfxtp_4
Xsky130_fd_sc_hs__nand2_2_2 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_2_3/Y sky130_fd_sc_hs__nand2_2_3/B
+ eqn[25] sky130_fd_sc_hs__nand2_2_3/a_27_74# sky130_fd_sc_hs__nand2_2
Xsky130_fd_sc_hs__xnor2_1_4 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__xnor2_1_5/A sky130_fd_sc_hs__xnor2_1_5/Y
+ sky130_fd_sc_hs__xnor2_1_7/Y sky130_fd_sc_hs__xnor2_1_5/a_376_368# sky130_fd_sc_hs__xnor2_1_5/a_112_119#
+ sky130_fd_sc_hs__xnor2_1_5/a_138_385# sky130_fd_sc_hs__xnor2_1_5/a_293_74# sky130_fd_sc_hs__xnor2_1
Xsky130_fd_sc_hs__a22o_1_11 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__dfxtp_4_8/D sky130_fd_sc_hs__nand2_1_21/B
+ sky130_fd_sc_hs__and2b_2_1/X init_val[8] rst sky130_fd_sc_hs__a22o_1_11/a_222_392#
+ sky130_fd_sc_hs__a22o_1_11/a_230_79# sky130_fd_sc_hs__a22o_1_11/a_52_123# sky130_fd_sc_hs__a22o_1_11/a_132_392#
+ sky130_fd_sc_hs__a22o_1
Xsky130_fd_sc_hs__a22o_1_22 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__a22o_1_23/X sky130_fd_sc_hs__nand2_1_5/B
+ sky130_fd_sc_hs__and2b_2_1/X init_val[6] rst sky130_fd_sc_hs__a22o_1_23/a_222_392#
+ sky130_fd_sc_hs__a22o_1_23/a_230_79# sky130_fd_sc_hs__a22o_1_23/a_52_123# sky130_fd_sc_hs__a22o_1_23/a_132_392#
+ sky130_fd_sc_hs__a22o_1
Xsky130_fd_sc_hs__a22o_1_33 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__a22o_1_33/X sky130_fd_sc_hs__nand2_1_45/B
+ sky130_fd_sc_hs__and2b_2_1/X init_val[2] rst sky130_fd_sc_hs__a22o_1_33/a_222_392#
+ sky130_fd_sc_hs__a22o_1_33/a_230_79# sky130_fd_sc_hs__a22o_1_33/a_52_123# sky130_fd_sc_hs__a22o_1_33/a_132_392#
+ sky130_fd_sc_hs__a22o_1
Xsky130_fd_sc_hs__a22o_1_55 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__a22o_1_55/X sky130_fd_sc_hs__nand2_1_51/B
+ sky130_fd_sc_hs__and2b_2_1/X init_val[23] rst sky130_fd_sc_hs__a22o_1_55/a_222_392#
+ sky130_fd_sc_hs__a22o_1_55/a_230_79# sky130_fd_sc_hs__a22o_1_55/a_52_123# sky130_fd_sc_hs__a22o_1_55/a_132_392#
+ sky130_fd_sc_hs__a22o_1
Xsky130_fd_sc_hs__a22o_1_44 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__a22o_1_45/X sky130_fd_sc_hs__nand2_1_41/B
+ sky130_fd_sc_hs__and2b_2_1/X init_val[1] rst sky130_fd_sc_hs__a22o_1_45/a_222_392#
+ sky130_fd_sc_hs__a22o_1_45/a_230_79# sky130_fd_sc_hs__a22o_1_45/a_52_123# sky130_fd_sc_hs__a22o_1_45/a_132_392#
+ sky130_fd_sc_hs__a22o_1
Xsky130_fd_sc_hs__nand2_1_11 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__dfxtp_4_7/Q sky130_fd_sc_hs__xnor2_1_35/B
+ eqn[10] sky130_fd_sc_hs__nand2_1_11/a_117_74# sky130_fd_sc_hs__nand2_1
Xsky130_fd_sc_hs__nand2_1_22 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_1_23/B sky130_fd_sc_hs__xnor2_1_15/B
+ eqn[2] sky130_fd_sc_hs__nand2_1_23/a_117_74# sky130_fd_sc_hs__nand2_1
Xsky130_fd_sc_hs__nand2_1_33 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_1_33/B sky130_fd_sc_hs__xnor2_1_21/B
+ eqn[20] sky130_fd_sc_hs__nand2_1_33/a_117_74# sky130_fd_sc_hs__nand2_1
Xsky130_fd_sc_hs__nand2_1_44 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_1_45/B sky130_fd_sc_hs__xnor2_1_61/B
+ eqn[1] sky130_fd_sc_hs__nand2_1_45/a_117_74# sky130_fd_sc_hs__nand2_1
Xsky130_fd_sc_hs__nand2_1_55 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_1_55/B sky130_fd_sc_hs__xnor2_1_31/B
+ eqn[29] sky130_fd_sc_hs__nand2_1_55/a_117_74# sky130_fd_sc_hs__nand2_1
Xsky130_fd_sc_hs__dfxtp_4_1 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__dfxtp_4_1/Q sky130_fd_sc_hs__a22o_1_1/X
+ sky130_fd_sc_hs__dfxtp_4_9/CLK sky130_fd_sc_hs__dfxtp_4_1/a_1226_296# sky130_fd_sc_hs__dfxtp_4_1/a_735_102#
+ sky130_fd_sc_hs__dfxtp_4_1/a_1141_508# sky130_fd_sc_hs__dfxtp_4_1/a_206_368# sky130_fd_sc_hs__dfxtp_4_1/a_437_503#
+ sky130_fd_sc_hs__dfxtp_4_1/a_27_74# sky130_fd_sc_hs__dfxtp_4_1/a_651_503# sky130_fd_sc_hs__dfxtp_4_1/a_696_458#
+ sky130_fd_sc_hs__dfxtp_4_1/a_544_485# sky130_fd_sc_hs__dfxtp_4_1/a_1178_124# sky130_fd_sc_hs__dfxtp_4_1/a_1034_424#
+ sky130_fd_sc_hs__dfxtp_4
Xsky130_fd_sc_hs__dfxtp_4_18 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_1_29/B sky130_fd_sc_hs__a22o_1_23/X
+ sky130_fd_sc_hs__dfxtp_4_9/CLK sky130_fd_sc_hs__dfxtp_4_19/a_1226_296# sky130_fd_sc_hs__dfxtp_4_19/a_735_102#
+ sky130_fd_sc_hs__dfxtp_4_19/a_1141_508# sky130_fd_sc_hs__dfxtp_4_19/a_206_368# sky130_fd_sc_hs__dfxtp_4_19/a_437_503#
+ sky130_fd_sc_hs__dfxtp_4_19/a_27_74# sky130_fd_sc_hs__dfxtp_4_19/a_651_503# sky130_fd_sc_hs__dfxtp_4_19/a_696_458#
+ sky130_fd_sc_hs__dfxtp_4_19/a_544_485# sky130_fd_sc_hs__dfxtp_4_19/a_1178_124# sky130_fd_sc_hs__dfxtp_4_19/a_1034_424#
+ sky130_fd_sc_hs__dfxtp_4
Xsky130_fd_sc_hs__dfxtp_4_29 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_1_17/B sky130_fd_sc_hs__a22o_1_29/X
+ sky130_fd_sc_hs__dfxtp_4_9/CLK sky130_fd_sc_hs__dfxtp_4_29/a_1226_296# sky130_fd_sc_hs__dfxtp_4_29/a_735_102#
+ sky130_fd_sc_hs__dfxtp_4_29/a_1141_508# sky130_fd_sc_hs__dfxtp_4_29/a_206_368# sky130_fd_sc_hs__dfxtp_4_29/a_437_503#
+ sky130_fd_sc_hs__dfxtp_4_29/a_27_74# sky130_fd_sc_hs__dfxtp_4_29/a_651_503# sky130_fd_sc_hs__dfxtp_4_29/a_696_458#
+ sky130_fd_sc_hs__dfxtp_4_29/a_544_485# sky130_fd_sc_hs__dfxtp_4_29/a_1178_124# sky130_fd_sc_hs__dfxtp_4_29/a_1034_424#
+ sky130_fd_sc_hs__dfxtp_4
Xsky130_fd_sc_hs__nand2_2_3 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_2_3/Y sky130_fd_sc_hs__nand2_2_3/B
+ eqn[25] sky130_fd_sc_hs__nand2_2_3/a_27_74# sky130_fd_sc_hs__nand2_2
Xsky130_fd_sc_hs__xnor2_1_5 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__xnor2_1_5/A sky130_fd_sc_hs__xnor2_1_5/Y
+ sky130_fd_sc_hs__xnor2_1_7/Y sky130_fd_sc_hs__xnor2_1_5/a_376_368# sky130_fd_sc_hs__xnor2_1_5/a_112_119#
+ sky130_fd_sc_hs__xnor2_1_5/a_138_385# sky130_fd_sc_hs__xnor2_1_5/a_293_74# sky130_fd_sc_hs__xnor2_1
Xsky130_fd_sc_hs__a22o_1_12 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__a22o_1_13/X sky130_fd_sc_hs__nand2_1_13/B
+ sky130_fd_sc_hs__and2b_2_1/X init_val[16] rst sky130_fd_sc_hs__a22o_1_13/a_222_392#
+ sky130_fd_sc_hs__a22o_1_13/a_230_79# sky130_fd_sc_hs__a22o_1_13/a_52_123# sky130_fd_sc_hs__a22o_1_13/a_132_392#
+ sky130_fd_sc_hs__a22o_1
Xsky130_fd_sc_hs__a22o_1_23 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__a22o_1_23/X sky130_fd_sc_hs__nand2_1_5/B
+ sky130_fd_sc_hs__and2b_2_1/X init_val[6] rst sky130_fd_sc_hs__a22o_1_23/a_222_392#
+ sky130_fd_sc_hs__a22o_1_23/a_230_79# sky130_fd_sc_hs__a22o_1_23/a_52_123# sky130_fd_sc_hs__a22o_1_23/a_132_392#
+ sky130_fd_sc_hs__a22o_1
Xsky130_fd_sc_hs__a22o_1_34 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__a22o_1_35/X sky130_fd_sc_hs__nand2_1_33/B
+ sky130_fd_sc_hs__and2b_2_1/X init_val[21] rst sky130_fd_sc_hs__a22o_1_35/a_222_392#
+ sky130_fd_sc_hs__a22o_1_35/a_230_79# sky130_fd_sc_hs__a22o_1_35/a_52_123# sky130_fd_sc_hs__a22o_1_35/a_132_392#
+ sky130_fd_sc_hs__a22o_1
Xsky130_fd_sc_hs__a22o_1_56 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__a22o_1_57/X sky130_fd_sc_hs__nand2_1_37/B
+ sky130_fd_sc_hs__and2b_2_1/X init_val[25] rst sky130_fd_sc_hs__a22o_1_57/a_222_392#
+ sky130_fd_sc_hs__a22o_1_57/a_230_79# sky130_fd_sc_hs__a22o_1_57/a_52_123# sky130_fd_sc_hs__a22o_1_57/a_132_392#
+ sky130_fd_sc_hs__a22o_1
Xsky130_fd_sc_hs__a22o_1_45 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__a22o_1_45/X sky130_fd_sc_hs__nand2_1_41/B
+ sky130_fd_sc_hs__and2b_2_1/X init_val[1] rst sky130_fd_sc_hs__a22o_1_45/a_222_392#
+ sky130_fd_sc_hs__a22o_1_45/a_230_79# sky130_fd_sc_hs__a22o_1_45/a_52_123# sky130_fd_sc_hs__a22o_1_45/a_132_392#
+ sky130_fd_sc_hs__a22o_1
Xsky130_fd_sc_hs__nand2_1_12 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_1_13/B sky130_fd_sc_hs__xnor2_1_13/B
+ eqn[15] sky130_fd_sc_hs__nand2_1_13/a_117_74# sky130_fd_sc_hs__nand2_1
Xsky130_fd_sc_hs__nand2_1_23 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_1_23/B sky130_fd_sc_hs__xnor2_1_15/B
+ eqn[2] sky130_fd_sc_hs__nand2_1_23/a_117_74# sky130_fd_sc_hs__nand2_1
Xsky130_fd_sc_hs__nand2_1_34 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_1_35/B sky130_fd_sc_hs__xnor2_1_37/A
+ eqn[23] sky130_fd_sc_hs__nand2_1_35/a_117_74# sky130_fd_sc_hs__nand2_1
Xsky130_fd_sc_hs__nand2_1_45 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_1_45/B sky130_fd_sc_hs__xnor2_1_61/B
+ eqn[1] sky130_fd_sc_hs__nand2_1_45/a_117_74# sky130_fd_sc_hs__nand2_1
Xsky130_fd_sc_hs__nand2_1_56 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_1_57/B sky130_fd_sc_hs__xnor2_1_53/B
+ eqn[30] sky130_fd_sc_hs__nand2_1_57/a_117_74# sky130_fd_sc_hs__nand2_1
Xsky130_fd_sc_hs__dfxtp_4_2 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_2_1/B sky130_fd_sc_hs__a22o_1_5/X
+ sky130_fd_sc_hs__dfxtp_4_9/CLK sky130_fd_sc_hs__dfxtp_4_4/a_1226_296# sky130_fd_sc_hs__dfxtp_4_4/a_735_102#
+ sky130_fd_sc_hs__dfxtp_4_4/a_1141_508# sky130_fd_sc_hs__dfxtp_4_4/a_206_368# sky130_fd_sc_hs__dfxtp_4_4/a_437_503#
+ sky130_fd_sc_hs__dfxtp_4_4/a_27_74# sky130_fd_sc_hs__dfxtp_4_4/a_651_503# sky130_fd_sc_hs__dfxtp_4_4/a_696_458#
+ sky130_fd_sc_hs__dfxtp_4_4/a_544_485# sky130_fd_sc_hs__dfxtp_4_4/a_1178_124# sky130_fd_sc_hs__dfxtp_4_4/a_1034_424#
+ sky130_fd_sc_hs__dfxtp_4
Xsky130_fd_sc_hs__dfxtp_4_19 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_1_29/B sky130_fd_sc_hs__a22o_1_23/X
+ sky130_fd_sc_hs__dfxtp_4_9/CLK sky130_fd_sc_hs__dfxtp_4_19/a_1226_296# sky130_fd_sc_hs__dfxtp_4_19/a_735_102#
+ sky130_fd_sc_hs__dfxtp_4_19/a_1141_508# sky130_fd_sc_hs__dfxtp_4_19/a_206_368# sky130_fd_sc_hs__dfxtp_4_19/a_437_503#
+ sky130_fd_sc_hs__dfxtp_4_19/a_27_74# sky130_fd_sc_hs__dfxtp_4_19/a_651_503# sky130_fd_sc_hs__dfxtp_4_19/a_696_458#
+ sky130_fd_sc_hs__dfxtp_4_19/a_544_485# sky130_fd_sc_hs__dfxtp_4_19/a_1178_124# sky130_fd_sc_hs__dfxtp_4_19/a_1034_424#
+ sky130_fd_sc_hs__dfxtp_4
Xsky130_fd_sc_hs__nand2_2_4 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_2_5/Y sky130_fd_sc_hs__nand2_2_5/B
+ eqn[31] sky130_fd_sc_hs__nand2_2_5/a_27_74# sky130_fd_sc_hs__nand2_2
Xsky130_fd_sc_hs__xnor2_1_6 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__xnor2_1_7/A sky130_fd_sc_hs__xnor2_1_7/Y
+ sky130_fd_sc_hs__xnor2_1_9/Y sky130_fd_sc_hs__xnor2_1_7/a_376_368# sky130_fd_sc_hs__xnor2_1_7/a_112_119#
+ sky130_fd_sc_hs__xnor2_1_7/a_138_385# sky130_fd_sc_hs__xnor2_1_7/a_293_74# sky130_fd_sc_hs__xnor2_1
Xsky130_fd_sc_hs__a22o_1_13 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__a22o_1_13/X sky130_fd_sc_hs__nand2_1_13/B
+ sky130_fd_sc_hs__and2b_2_1/X init_val[16] rst sky130_fd_sc_hs__a22o_1_13/a_222_392#
+ sky130_fd_sc_hs__a22o_1_13/a_230_79# sky130_fd_sc_hs__a22o_1_13/a_52_123# sky130_fd_sc_hs__a22o_1_13/a_132_392#
+ sky130_fd_sc_hs__a22o_1
Xsky130_fd_sc_hs__a22o_1_24 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__a22o_1_25/X sky130_fd_sc_hs__nand2_1_9/B
+ sky130_fd_sc_hs__and2b_2_1/X init_val[5] rst sky130_fd_sc_hs__a22o_1_25/a_222_392#
+ sky130_fd_sc_hs__a22o_1_25/a_230_79# sky130_fd_sc_hs__a22o_1_25/a_52_123# sky130_fd_sc_hs__a22o_1_25/a_132_392#
+ sky130_fd_sc_hs__a22o_1
Xsky130_fd_sc_hs__a22o_1_35 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__a22o_1_35/X sky130_fd_sc_hs__nand2_1_33/B
+ sky130_fd_sc_hs__and2b_2_1/X init_val[21] rst sky130_fd_sc_hs__a22o_1_35/a_222_392#
+ sky130_fd_sc_hs__a22o_1_35/a_230_79# sky130_fd_sc_hs__a22o_1_35/a_52_123# sky130_fd_sc_hs__a22o_1_35/a_132_392#
+ sky130_fd_sc_hs__a22o_1
Xsky130_fd_sc_hs__a22o_1_57 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__a22o_1_57/X sky130_fd_sc_hs__nand2_1_37/B
+ sky130_fd_sc_hs__and2b_2_1/X init_val[25] rst sky130_fd_sc_hs__a22o_1_57/a_222_392#
+ sky130_fd_sc_hs__a22o_1_57/a_230_79# sky130_fd_sc_hs__a22o_1_57/a_52_123# sky130_fd_sc_hs__a22o_1_57/a_132_392#
+ sky130_fd_sc_hs__a22o_1
Xsky130_fd_sc_hs__a22o_1_46 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__a22o_1_47/X sky130_fd_sc_hs__nand2_1_49/B
+ sky130_fd_sc_hs__and2b_2_1/X init_val[29] rst sky130_fd_sc_hs__a22o_1_47/a_222_392#
+ sky130_fd_sc_hs__a22o_1_47/a_230_79# sky130_fd_sc_hs__a22o_1_47/a_52_123# sky130_fd_sc_hs__a22o_1_47/a_132_392#
+ sky130_fd_sc_hs__a22o_1
Xsky130_fd_sc_hs__nand2_1_13 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_1_13/B sky130_fd_sc_hs__xnor2_1_13/B
+ eqn[15] sky130_fd_sc_hs__nand2_1_13/a_117_74# sky130_fd_sc_hs__nand2_1
Xsky130_fd_sc_hs__nand2_1_24 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_1_25/B sky130_fd_sc_hs__xnor2_1_31/A
+ eqn[14] sky130_fd_sc_hs__nand2_1_25/a_117_74# sky130_fd_sc_hs__nand2_1
Xsky130_fd_sc_hs__nand2_1_35 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_1_35/B sky130_fd_sc_hs__xnor2_1_37/A
+ eqn[23] sky130_fd_sc_hs__nand2_1_35/a_117_74# sky130_fd_sc_hs__nand2_1
Xsky130_fd_sc_hs__nand2_1_46 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_1_47/B sky130_fd_sc_hs__xnor2_1_55/B
+ eqn[19] sky130_fd_sc_hs__nand2_1_47/a_117_74# sky130_fd_sc_hs__nand2_1
Xsky130_fd_sc_hs__nand2_1_57 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_1_57/B sky130_fd_sc_hs__xnor2_1_53/B
+ eqn[30] sky130_fd_sc_hs__nand2_1_57/a_117_74# sky130_fd_sc_hs__nand2_1
Xsky130_fd_sc_hs__dfxtp_4_3 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_1_3/B sky130_fd_sc_hs__a22o_1_3/X
+ sky130_fd_sc_hs__dfxtp_4_9/CLK sky130_fd_sc_hs__dfxtp_4_5/a_1226_296# sky130_fd_sc_hs__dfxtp_4_5/a_735_102#
+ sky130_fd_sc_hs__dfxtp_4_5/a_1141_508# sky130_fd_sc_hs__dfxtp_4_5/a_206_368# sky130_fd_sc_hs__dfxtp_4_5/a_437_503#
+ sky130_fd_sc_hs__dfxtp_4_5/a_27_74# sky130_fd_sc_hs__dfxtp_4_5/a_651_503# sky130_fd_sc_hs__dfxtp_4_5/a_696_458#
+ sky130_fd_sc_hs__dfxtp_4_5/a_544_485# sky130_fd_sc_hs__dfxtp_4_5/a_1178_124# sky130_fd_sc_hs__dfxtp_4_5/a_1034_424#
+ sky130_fd_sc_hs__dfxtp_4
Xsky130_fd_sc_hs__nand2_2_5 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_2_5/Y sky130_fd_sc_hs__nand2_2_5/B
+ eqn[31] sky130_fd_sc_hs__nand2_2_5/a_27_74# sky130_fd_sc_hs__nand2_2
.ends

.subckt sky130_fd_sc_hs__or2b_2 VNB VPB VPWR VGND X B_N A a_470_368# a_27_368# a_187_48#
X0 VGND B_N a_27_368# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=550000u l=150000u
X1 VGND a_27_368# a_187_48# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X2 VPWR a_187_48# X VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X3 VGND a_187_48# X VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X4 a_187_48# A VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X5 a_187_48# a_27_368# a_470_368# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 a_470_368# A VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 X a_187_48# VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X8 X a_187_48# VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X9 VPWR B_N a_27_368# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
.ends

.subckt sky130_fd_sc_hs__o21ai_2 VNB VPB VPWR VGND B1 A2 A1 Y a_116_368# a_27_74#
X0 a_27_74# B1 Y VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X1 a_27_74# A1 VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X2 VGND A1 a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X3 a_116_368# A2 Y VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X4 VGND A2 a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X5 Y B1 a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X6 Y A2 a_116_368# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X7 a_27_74# A2 VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X8 VPWR B1 Y VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X9 Y B1 VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X10 a_116_368# A1 VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X11 VPWR A1 a_116_368# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
.ends

.subckt sky130_fd_sc_hs__einvp_8 VNB VPB VPWR VGND Z TE A a_802_323# a_27_74# a_27_368#
X0 a_27_74# TE VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X1 VPWR a_802_323# a_27_368# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X2 a_27_368# A Z VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X3 a_27_74# A Z VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X4 a_27_74# A Z VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X5 Z A a_27_368# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X6 a_27_74# TE VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X7 a_27_368# A Z VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X8 Z A a_27_368# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X9 Z A a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X10 a_27_74# TE VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X11 a_27_368# A Z VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X12 VGND TE a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X13 Z A a_27_368# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X14 VPWR TE a_802_323# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X15 Z A a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X16 a_27_368# A Z VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X17 Z A a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X18 VGND TE a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X19 VGND TE a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X20 a_27_368# a_802_323# VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X21 a_27_74# A Z VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X22 VPWR a_802_323# a_27_368# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X23 a_27_74# A Z VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X24 VGND TE a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X25 a_27_368# a_802_323# VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X26 VPWR a_802_323# a_27_368# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X27 VPWR a_802_323# a_27_368# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X28 a_27_368# a_802_323# VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X29 a_27_368# a_802_323# VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X30 Z A a_27_368# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X31 a_27_74# TE VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X32 VGND TE a_802_323# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X33 Z A a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
.ends

.subckt sky130_fd_sc_hs__diode_2 DIODE VNB VPB VPWR VGND
X0 VNB DIODE sky130_fd_pr__diode_pw2nd_05v5 area=6.417e+11p
.ends

.subckt sky130_fd_sc_hs__einvn_1 VNB VPB VPWR VGND A Z TE_B a_281_100# a_278_368#
+ a_22_46#
X0 Z A a_278_368# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X1 VGND TE_B a_22_46# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 a_278_368# TE_B VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X3 VPWR TE_B a_22_46# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X4 Z A a_281_100# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X5 a_281_100# a_22_46# VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
.ends

.subckt sky130_fd_sc_hs__o22ai_1 VNB VPB VPWR VGND B2 B1 Y A2 A1 a_340_368# a_142_368#
+ a_27_74#
X0 Y B2 a_142_368# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X1 a_27_74# B2 Y VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X2 Y B1 a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X3 a_27_74# A1 VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X4 a_142_368# B1 VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X5 a_340_368# A2 Y VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X6 VPWR A1 a_340_368# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X7 VGND A2 a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
.ends

.subckt sky130_fd_sc_hs__nand2_4 VNB VPB VPWR VGND Y B A a_27_74#
X0 Y B VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X1 VPWR A Y VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X2 Y A VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X3 Y A a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X4 VGND B a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X5 a_27_74# A Y VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X6 VPWR B Y VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X7 a_27_74# B VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X8 a_27_74# A Y VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X9 a_27_74# B VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X10 VGND B a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X11 Y A a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
.ends

.subckt sky130_fd_sc_hs__o21ai_1 VNB VPB VPWR VGND Y B1 A2 A1 a_162_368# a_27_74#
X0 a_27_74# A2 VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X1 VGND A1 a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X2 Y B1 a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X3 Y A2 a_162_368# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X4 a_162_368# A1 VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X5 VPWR B1 Y VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
.ends

.subckt sky130_fd_sc_hs__inv_2 VNB VPB VPWR VGND A Y
X0 Y A VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X1 VPWR A Y VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X2 VGND A Y VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X3 Y A VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
.ends

.subckt sky130_fd_sc_hs__dfxtp_2 VNB VPB VPWR VGND Q CLK D a_431_508# a_1125_508#
+ a_206_368# a_27_74# a_708_101# a_1019_424# a_1172_124# a_644_504# a_1217_314# a_538_429#
+ a_695_459#
X0 VPWR a_1217_314# Q VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X1 a_1019_424# a_27_74# a_695_459# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X2 Q a_1217_314# VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X3 a_206_368# a_27_74# VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X4 a_644_504# a_27_74# a_538_429# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 VPWR a_1019_424# a_1217_314# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 VGND a_1217_314# a_1172_124# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7 a_538_429# a_27_74# a_431_508# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8 VGND CLK a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X9 a_1172_124# a_27_74# a_1019_424# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10 VGND a_695_459# a_708_101# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11 a_1125_508# a_206_368# a_1019_424# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12 VGND a_1217_314# Q VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X13 a_1019_424# a_206_368# a_695_459# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=550000u l=150000u
X14 a_206_368# a_27_74# VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X15 a_708_101# a_206_368# a_538_429# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16 a_695_459# a_538_429# VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X17 a_431_508# D VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18 a_538_429# a_206_368# a_431_508# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19 VPWR a_695_459# a_644_504# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20 VPWR a_1217_314# a_1125_508# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21 Q a_1217_314# VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X22 VGND a_1019_424# a_1217_314# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X23 a_695_459# a_538_429# VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=550000u l=150000u
X24 a_431_508# D VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X25 VPWR CLK a_27_74# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
.ends

.subckt sky130_fd_sc_hs__a21oi_1 VNB VPB VPWR VGND B1 Y A2 A1 a_117_74# a_29_368#
X0 Y A1 a_117_74# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X1 a_117_74# A2 VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X2 Y B1 a_29_368# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X3 a_29_368# A1 VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X4 VPWR A2 a_29_368# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X5 VGND B1 Y VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
.ends

.subckt sky130_fd_sc_hs__maj3_1 VNB VPB VPWR VGND A B X C a_598_384# a_226_384# a_84_74#
+ a_403_136# a_406_384# a_595_136# a_223_120#
X0 a_406_384# B a_84_74# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_598_384# A VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 a_226_384# A VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 VGND C a_403_136# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X4 a_84_74# C a_595_136# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X5 a_403_136# B a_84_74# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X6 a_595_136# A VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X7 VGND a_84_74# X VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X8 VPWR a_84_74# X VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X9 a_84_74# B a_223_120# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X10 a_223_120# A VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X11 VPWR C a_406_384# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 a_84_74# C a_598_384# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13 a_84_74# B a_226_384# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_sc_hs__nor2_2 VNB VPB VPWR VGND B Y A a_35_368#
X0 Y B VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X1 Y B a_35_368# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X2 VGND A Y VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X3 a_35_368# A VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X4 VPWR A a_35_368# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X5 a_35_368# B Y VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
.ends

.subckt sky130_fd_sc_hs__nor2_1 VNB VPB VPWR VGND B Y A a_116_368#
X0 Y A VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X1 Y B a_116_368# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X2 VGND B Y VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X3 a_116_368# A VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
.ends

.subckt sky130_fd_sc_hs__nand3_1 VNB VPB VPWR VGND C Y B A a_155_74# a_233_74#
X0 VPWR B Y VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X1 a_233_74# B a_155_74# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X2 Y C VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X3 Y A VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X4 a_155_74# C VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X5 Y A a_233_74# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
.ends

.subckt sky130_fd_sc_hs__dfrtp_4 VNB VPB RESET_B VPWR VGND D CLK Q a_37_78# a_494_366#
+ a_699_463# a_313_74# a_1627_493# a_1678_395# a_1827_81# a_789_463# a_1350_392# a_834_355#
+ a_812_138# a_124_78# a_1647_81# a_2010_409# a_890_138#
X0 a_37_78# D VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1 a_834_355# a_699_463# VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X2 VPWR a_2010_409# Q VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X3 VPWR a_1678_395# a_1627_493# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4 a_1647_81# a_313_74# a_1350_392# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 VGND CLK a_313_74# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X6 VPWR a_1350_392# a_1678_395# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7 a_699_463# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8 a_1627_493# a_494_366# a_1350_392# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9 a_1678_395# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10 VGND RESET_B a_890_138# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11 a_1827_81# RESET_B VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12 Q a_2010_409# VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X13 a_1350_392# a_313_74# a_834_355# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14 a_890_138# a_834_355# a_812_138# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15 a_834_355# a_699_463# VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16 Q a_2010_409# VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X17 a_812_138# a_494_366# a_699_463# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18 VGND a_2010_409# Q VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X19 VPWR a_1350_392# a_2010_409# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X20 Q a_2010_409# VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X21 VGND a_1678_395# a_1647_81# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22 VGND a_2010_409# Q VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X23 VPWR RESET_B a_37_78# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24 VPWR a_834_355# a_789_463# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X25 a_1678_395# a_1350_392# a_1827_81# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X26 a_699_463# a_313_74# a_37_78# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X27 a_1350_392# a_494_366# a_834_355# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X28 a_124_78# D a_37_78# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X29 a_789_463# a_313_74# a_699_463# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X30 a_2010_409# a_1350_392# VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X31 VPWR a_2010_409# Q VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X32 Q a_2010_409# VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X33 a_699_463# a_494_366# a_37_78# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X34 a_2010_409# a_1350_392# VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X35 a_494_366# a_313_74# VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X36 VPWR CLK a_313_74# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X37 VGND RESET_B a_124_78# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X38 a_494_366# a_313_74# VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
.ends

.subckt sky130_fd_sc_hs__o31ai_1 VNB VPB VPWR VGND A3 A2 B1 A1 Y a_114_74# a_119_368#
+ a_203_368#
X0 VPWR B1 Y VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X1 a_203_368# A2 a_119_368# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X2 Y A3 a_203_368# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X3 a_114_74# A1 VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X4 Y B1 a_114_74# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X5 a_119_368# A1 VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X6 VGND A2 a_114_74# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X7 a_114_74# A3 VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
.ends

.subckt sky130_fd_sc_hs__dfrtn_1 VNB VPB RESET_B VPWR VGND CLK_N Q D a_1266_119# a_1736_119#
+ a_817_508# a_120_74# a_1547_508# a_922_127# a_33_74# a_714_127# a_1934_94# a_1550_119#
+ a_1598_93# a_300_74# a_507_368# a_856_304# a_850_127#
X0 a_1266_119# a_300_74# a_856_304# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X1 a_33_74# D VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 a_856_304# a_714_127# VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 a_1266_119# a_507_368# a_856_304# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 a_714_127# a_507_368# a_33_74# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 VPWR a_1266_119# a_1598_93# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 VGND RESET_B a_120_74# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7 a_507_368# a_300_74# VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X8 a_1736_119# RESET_B VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9 a_300_74# CLK_N VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X10 VPWR a_1598_93# a_1547_508# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11 a_1550_119# a_507_368# a_1266_119# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12 a_850_127# a_300_74# a_714_127# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13 a_856_304# a_714_127# VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X14 a_300_74# CLK_N VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X15 a_1547_508# a_300_74# a_1266_119# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16 a_1598_93# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17 a_120_74# D a_33_74# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18 Q a_1934_94# VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X19 VPWR RESET_B a_33_74# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20 VGND a_1266_119# a_1934_94# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=550000u l=150000u
X21 VGND RESET_B a_922_127# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22 VPWR a_856_304# a_817_508# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23 VPWR a_1266_119# a_1934_94# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X24 a_507_368# a_300_74# VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X25 a_714_127# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X26 Q a_1934_94# VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X27 a_1598_93# a_1266_119# a_1736_119# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X28 a_922_127# a_856_304# a_850_127# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X29 VGND a_1598_93# a_1550_119# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X30 a_817_508# a_507_368# a_714_127# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X31 a_714_127# a_300_74# a_33_74# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
.ends

.subckt sky130_fd_sc_hs__dfstp_2 VNB VPB SET_B VPWR VGND CLK D Q a_1566_92# a_1521_508#
+ a_716_456# a_1266_341# a_1278_74# a_398_74# a_1057_118# a_1489_118# a_27_74# a_1596_118#
+ a_225_74# a_1356_74# a_612_74# a_781_74# a_767_384# a_2022_94#
X0 a_1596_118# a_1566_92# a_1489_118# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1 VPWR a_767_384# a_716_456# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 VGND a_1356_74# a_2022_94# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X3 a_1489_118# a_225_74# a_1356_74# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4 VGND SET_B a_1596_118# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 a_716_456# a_225_74# a_612_74# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 VPWR D a_27_74# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7 VGND D a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8 a_1356_74# a_225_74# a_1266_341# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 a_1566_92# a_1356_74# VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10 a_1356_74# a_398_74# a_1278_74# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X11 a_612_74# a_398_74# a_27_74# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12 a_767_384# a_612_74# VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13 VPWR SET_B a_767_384# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14 VGND CLK a_225_74# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X15 VPWR a_1566_92# a_1521_508# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16 VPWR a_2022_94# Q VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X17 VGND SET_B a_1057_118# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18 Q a_2022_94# VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X19 a_1521_508# a_398_74# a_1356_74# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20 a_1356_74# SET_B VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21 VGND a_2022_94# Q VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X22 a_398_74# a_225_74# VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X23 a_1266_341# a_612_74# VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X24 VPWR a_1356_74# a_2022_94# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X25 VGND a_767_384# a_781_74# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X26 VPWR CLK a_225_74# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X27 a_398_74# a_225_74# VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X28 a_1057_118# a_612_74# a_767_384# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X29 a_1566_92# a_1356_74# VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X30 a_612_74# a_225_74# a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X31 a_781_74# a_398_74# a_612_74# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X32 Q a_2022_94# VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X33 a_1278_74# a_612_74# VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
.ends

.subckt sky130_fd_sc_hs__dfrbp_1 VNB VPB RESET_B VPWR VGND Q CLK D Q_N a_498_360#
+ a_1224_74# a_2026_424# a_1482_48# a_125_78# a_796_463# a_910_118# a_1465_471# a_832_118#
+ a_841_401# a_38_78# a_1434_74# a_706_463# a_319_360# a_1624_74#
X0 a_796_463# a_319_360# a_706_463# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1 a_841_401# a_706_463# VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X2 a_706_463# a_498_360# a_38_78# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3 Q_N a_1224_74# VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X4 a_706_463# a_319_360# a_38_78# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 a_498_360# a_319_360# VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X6 a_38_78# D VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7 a_1624_74# RESET_B VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8 a_1224_74# a_498_360# a_841_401# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X9 a_706_463# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10 VGND RESET_B a_910_118# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11 VGND a_1482_48# a_1434_74# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12 a_910_118# a_841_401# a_832_118# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13 VPWR a_1482_48# a_1465_471# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14 VPWR a_1224_74# a_1482_48# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15 Q a_2026_424# VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X16 a_498_360# a_319_360# VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X17 a_1482_48# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18 a_1224_74# a_319_360# a_841_401# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X19 Q a_2026_424# VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X20 VPWR CLK a_319_360# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X21 a_1465_471# a_498_360# a_1224_74# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22 a_1482_48# a_1224_74# a_1624_74# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23 a_125_78# D a_38_78# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24 Q_N a_1224_74# VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X25 VPWR RESET_B a_38_78# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X26 a_832_118# a_498_360# a_706_463# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X27 VGND CLK a_319_360# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X28 VPWR a_1224_74# a_2026_424# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X29 a_1434_74# a_319_360# a_1224_74# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X30 VGND a_1224_74# a_2026_424# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=550000u l=150000u
X31 VPWR a_841_401# a_796_463# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X32 VGND RESET_B a_125_78# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X33 a_841_401# a_706_463# VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_sc_hs__a222o_1 VNB VPB VPWR VGND C2 X C1 B2 A2 A1 B1 a_27_390# a_386_74#
+ a_119_74# a_651_74# a_32_74# a_337_390#
X0 a_32_74# B1 a_386_74# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1 a_119_74# C1 a_32_74# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X2 a_27_390# B1 a_337_390# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 X a_32_74# VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X4 VGND C2 a_119_74# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X5 a_337_390# B2 a_27_390# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 a_32_74# C1 a_27_390# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 VGND A2 a_651_74# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X8 a_651_74# A1 a_32_74# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X9 a_27_390# C2 a_32_74# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 a_386_74# B2 VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X11 X a_32_74# VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X12 VPWR A2 a_337_390# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13 a_337_390# A1 VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_sc_hs__nor3_1 VNB VPB VPWR VGND Y C B A a_198_368# a_114_368#
X0 a_198_368# B a_114_368# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X1 Y C a_198_368# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X2 Y A VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X3 Y C VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X4 a_114_368# A VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X5 VGND B Y VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
.ends

.subckt sky130_fd_sc_hs__a22oi_1 VNB VPB VPWR VGND B2 Y B1 A2 A1 a_71_368# a_159_74#
+ a_339_74#
X0 Y B1 a_159_74# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X1 a_159_74# B2 VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X2 VGND A2 a_339_74# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X3 a_339_74# A1 Y VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X4 VPWR A1 a_71_368# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X5 a_71_368# B1 Y VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X6 Y B2 a_71_368# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X7 a_71_368# A2 VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
.ends

.subckt sky130_fd_sc_hs__a211oi_1 VNB VPB VPWR VGND C1 Y B1 A2 A1 a_354_368# a_71_368#
+ a_159_74#
X0 Y A1 a_159_74# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X1 a_159_74# A2 VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X2 Y C1 VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X3 VGND B1 Y VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X4 VPWR A2 a_71_368# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X5 Y C1 a_354_368# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X6 a_354_368# B1 a_71_368# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X7 a_71_368# A1 VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
.ends

.subckt sky130_fd_sc_hs__nand4_2 VNB VPB VPWR VGND Y C D B A a_304_74# a_27_74# a_515_74#
X0 a_515_74# A Y VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X1 VPWR D Y VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X2 Y D VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X3 VPWR C Y VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X4 VGND D a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X5 a_304_74# C a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X6 Y A a_515_74# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X7 Y C VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X8 a_27_74# D VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X9 a_304_74# B a_515_74# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X10 VPWR A Y VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X11 Y A VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X12 a_515_74# B a_304_74# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X13 VPWR B Y VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X14 Y B VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X15 a_27_74# C a_304_74# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
.ends

.subckt sky130_fd_sc_hs__sdlclkp_4 VNB VPB VPWR VGND SCE GATE CLK GCLK a_1289_368#
+ a_744_74# a_785_455# a_634_74# a_1292_74# a_792_48# a_324_79# a_116_395# a_354_105#
+ a_119_143#
X0 VPWR a_792_48# a_785_455# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1 a_634_74# a_324_79# a_119_143# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=550000u l=150000u
X2 a_116_395# SCE VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X3 a_354_105# a_324_79# VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X4 a_785_455# a_324_79# a_634_74# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 VPWR a_792_48# a_1289_368# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X6 a_119_143# SCE VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=550000u l=150000u
X7 a_634_74# a_354_105# a_119_143# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X8 a_792_48# a_634_74# VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X9 GCLK a_1289_368# VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X10 a_792_48# a_634_74# VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X11 a_1289_368# CLK VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X12 VGND a_792_48# a_744_74# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13 a_354_105# a_324_79# VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X14 VPWR CLK a_324_79# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X15 a_1292_74# CLK VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X16 a_119_143# GATE a_116_395# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X17 GCLK a_1289_368# VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X18 VPWR a_1289_368# GCLK VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X19 VGND GATE a_119_143# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=550000u l=150000u
X20 VGND CLK a_324_79# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X21 VGND a_1289_368# GCLK VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X22 VPWR a_1289_368# GCLK VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X23 GCLK a_1289_368# VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X24 VGND a_1289_368# GCLK VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X25 a_744_74# a_354_105# a_634_74# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X26 a_1289_368# a_792_48# a_1292_74# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X27 GCLK a_1289_368# VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
.ends

.subckt sky130_fd_sc_hs__xor2_1 VNB VPB VPWR VGND A B X a_194_125# a_355_368# a_455_87#
+ a_158_392#
X0 X B a_455_87# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X1 X a_194_125# a_355_368# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X2 a_194_125# B a_158_392# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 a_158_392# A VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 VPWR A a_355_368# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X5 a_355_368# B VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X6 a_194_125# A VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=550000u l=150000u
X7 a_455_87# A VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X8 VGND B a_194_125# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=550000u l=150000u
X9 VGND a_194_125# X VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
.ends

.subckt sky130_fd_sc_hs__fa_2 VNB VPB A VPWR VGND CIN B COUT SUM a_27_378# a_701_79#
+ a_484_347# a_1094_347# a_1205_79# a_27_79# a_1202_368# a_336_347# a_992_347# a_1119_79#
+ a_487_79# a_683_347#
X0 a_992_347# a_336_347# a_683_347# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 COUT a_336_347# VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X2 a_487_79# B a_336_347# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X3 a_336_347# CIN a_27_378# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 VPWR A a_484_347# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 a_683_347# A VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 a_701_79# CIN VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X7 VGND a_336_347# COUT VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X8 a_27_378# B VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 a_484_347# B a_336_347# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 VGND a_992_347# SUM VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X11 a_1094_347# CIN a_992_347# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 a_992_347# a_336_347# a_701_79# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X13 VGND B a_701_79# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X14 a_336_347# CIN a_27_79# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X15 a_683_347# CIN VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16 VPWR a_336_347# COUT VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X17 COUT a_336_347# VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X18 SUM a_992_347# VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X19 a_701_79# A VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X20 VGND A a_487_79# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X21 a_1205_79# B a_1119_79# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X22 VPWR B a_683_347# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X23 VPWR A a_27_378# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X24 a_1119_79# CIN a_992_347# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X25 VPWR a_992_347# SUM VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X26 VPWR A a_1202_368# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X27 SUM a_992_347# VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X28 a_1202_368# B a_1094_347# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X29 VGND A a_27_79# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X30 a_27_79# B VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X31 VGND A a_1205_79# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
.ends

.subckt sky130_fd_sc_hs__nand2b_1 VNB VPB VPWR VGND A_N B Y a_269_74# a_27_112#
X0 VPWR a_27_112# Y VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X1 a_269_74# B VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X2 Y B VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X3 VGND A_N a_27_112# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=550000u l=150000u
X4 Y a_27_112# a_269_74# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X5 VPWR A_N a_27_112# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
.ends

.subckt sky130_fd_sc_hs__o211ai_1 VNB VPB VPWR VGND B1 Y C1 A2 A1 a_31_74# a_311_74#
+ a_116_368#
X0 VGND A1 a_31_74# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X1 VPWR B1 Y VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X2 Y C1 a_311_74# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X3 Y A2 a_116_368# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X4 a_31_74# A2 VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X5 a_311_74# B1 a_31_74# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X6 Y C1 VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X7 a_116_368# A1 VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
.ends

.subckt sky130_fd_sc_hs__a222oi_1 VNB VPB VPWR VGND C2 C1 B1 A2 A1 Y B2 a_461_74#
+ a_697_74# a_119_74# a_116_392# a_369_392#
X0 a_116_392# C1 Y VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_369_392# B1 a_116_392# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 a_119_74# C1 Y VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X3 Y B1 a_461_74# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X4 a_461_74# B2 VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X5 VGND C2 a_119_74# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X6 Y C2 a_116_392# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 a_116_392# B2 a_369_392# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 VGND A2 a_697_74# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X9 VPWR A1 a_369_392# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 a_369_392# A2 VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 a_697_74# A1 Y VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
.ends

.subckt sky130_fd_sc_hs__a32oi_1 VNB VPB VPWR VGND A3 B2 B1 A2 Y A1 a_391_74# a_27_368#
+ a_119_74# a_469_74#
X0 a_119_74# B2 VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X1 VPWR A1 a_27_368# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X2 VGND A3 a_469_74# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X3 Y B1 a_119_74# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X4 a_27_368# B1 Y VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X5 VPWR A3 a_27_368# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X6 a_469_74# A2 a_391_74# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X7 a_27_368# A2 VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X8 a_391_74# A1 Y VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X9 Y B2 a_27_368# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
.ends

.subckt sky130_fd_sc_hs__a31oi_1 VNB VPB VPWR VGND Y A3 B1 A2 A1 a_136_368# a_223_74#
+ a_145_74#
X0 VPWR A2 a_136_368# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X1 a_136_368# A3 VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X2 a_145_74# A3 VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X3 Y B1 a_136_368# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X4 Y A1 a_223_74# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X5 a_136_368# A1 VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X6 a_223_74# A2 a_145_74# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X7 VGND B1 Y VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
.ends

.subckt sky130_fd_sc_hs__o21a_1 VNB VPB VPWR VGND X A2 B1 A1 a_320_74# a_376_387#
+ a_83_244#
X0 VGND a_83_244# X VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X1 a_320_74# A1 VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X2 a_320_74# B1 a_83_244# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X3 a_376_387# A2 a_83_244# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 a_83_244# B1 VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X5 VPWR A1 a_376_387# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 VGND A2 a_320_74# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X7 VPWR a_83_244# X VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
.ends

.subckt sky130_fd_sc_hs__nand3b_2 VNB VPB VPWR VGND Y A_N C B a_27_94# a_403_54# a_206_74#
X0 VGND C a_206_74# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X1 Y a_27_94# a_403_54# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X2 Y C VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X3 a_206_74# B a_403_54# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X4 a_206_74# C VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X5 VPWR A_N a_27_94# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 VPWR a_27_94# Y VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X7 a_403_54# a_27_94# Y VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X8 Y a_27_94# VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X9 a_403_54# B a_206_74# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X10 VGND A_N a_27_94# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X11 Y B VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X12 VPWR C Y VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X13 VPWR B Y VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
.ends

.subckt sky130_fd_sc_hs__o2bb2ai_1 VNB VPB VPWR VGND Y B2 A1_N B1 A2_N a_114_74# a_490_368#
+ a_397_74# a_131_383#
X0 a_131_383# A1_N VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X1 a_397_74# B1 VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X2 a_114_74# A1_N VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X3 a_131_383# A2_N a_114_74# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X4 VGND B2 a_397_74# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X5 a_397_74# a_131_383# Y VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X6 VPWR A2_N a_131_383# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X7 a_490_368# B2 Y VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X8 VPWR B1 a_490_368# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X9 Y a_131_383# VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
.ends

.subckt sky130_fd_sc_hs__a211oi_4 VNB VPB VPWR VGND Y C1 B1 A2 A1 a_901_368# a_77_368#
+ a_92_74#
X0 VGND B1 Y VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X1 Y A1 a_92_74# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X2 a_901_368# C1 Y VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X3 Y C1 a_901_368# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X4 a_77_368# A1 VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X5 a_92_74# A1 Y VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X6 VPWR A1 a_77_368# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X7 a_77_368# A1 VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X8 VPWR A1 a_77_368# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X9 a_92_74# A1 Y VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X10 a_92_74# A2 VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X11 a_901_368# C1 Y VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X12 Y C1 a_901_368# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X13 a_901_368# B1 a_77_368# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X14 a_92_74# A2 VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X15 Y C1 VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X16 a_77_368# B1 a_901_368# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X17 a_77_368# B1 a_901_368# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X18 a_901_368# B1 a_77_368# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X19 a_77_368# A2 VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X20 Y A1 a_92_74# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X21 Y B1 VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X22 VPWR A2 a_77_368# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X23 a_77_368# A2 VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X24 VGND A2 a_92_74# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X25 VPWR A2 a_77_368# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X26 VGND C1 Y VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X27 VGND A2 a_92_74# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
.ends

.subckt sky130_fd_sc_hs__a2bb2oi_1 VNB VPB VPWR VGND Y A2_N A1_N B2 B1 a_399_368#
+ a_126_112# a_117_392# a_488_74#
X0 Y a_126_112# VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X1 a_117_392# A1_N VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 VGND B1 a_488_74# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X3 a_488_74# B2 Y VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X4 a_126_112# A2_N a_117_392# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 VPWR B2 a_399_368# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X6 a_399_368# B1 VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X7 a_399_368# a_126_112# Y VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X8 VGND A2_N a_126_112# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=550000u l=150000u
X9 a_126_112# A1_N VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=550000u l=150000u
.ends

.subckt sky130_fd_sc_hs__dfsbp_2 VNB VPB SET_B VPWR VGND CLK D Q_N Q a_595_97# a_731_97#
+ a_1521_508# a_2221_74# a_1339_74# a_1531_118# a_1453_118# a_398_74# a_27_74# a_225_74#
+ a_1501_92# a_757_401# a_1258_341# a_1001_74# a_706_463# a_1261_74#
X0 a_1261_74# a_595_97# VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1 a_706_463# a_225_74# a_595_97# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 VPWR SET_B a_757_401# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3 a_595_97# a_398_74# a_27_74# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4 VGND a_1339_74# Q_N VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X5 Q_N a_1339_74# VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X6 VGND a_1339_74# a_2221_74# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X7 VPWR D a_27_74# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8 VGND D a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9 a_1258_341# a_595_97# VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 a_731_97# a_398_74# a_595_97# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11 VPWR a_1339_74# Q_N VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X12 VGND SET_B a_1531_118# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13 VGND a_757_401# a_731_97# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14 a_1339_74# SET_B VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15 Q a_2221_74# VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X16 VGND CLK a_225_74# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X17 VPWR a_1501_92# a_1521_508# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18 VPWR a_2221_74# Q VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X19 Q_N a_1339_74# VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X20 Q a_2221_74# VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X21 a_1521_508# a_398_74# a_1339_74# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22 VPWR a_1339_74# a_1501_92# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23 a_1001_74# a_595_97# a_757_401# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24 a_398_74# a_225_74# VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X25 VGND SET_B a_1001_74# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X26 a_1531_118# a_1501_92# a_1453_118# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X27 VGND a_2221_74# Q VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X28 VPWR CLK a_225_74# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X29 a_398_74# a_225_74# VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X30 a_595_97# a_225_74# a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X31 a_757_401# a_595_97# VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X32 VPWR a_1339_74# a_2221_74# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X33 a_1453_118# a_225_74# a_1339_74# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X34 a_1501_92# a_1339_74# VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X35 a_1339_74# a_398_74# a_1261_74# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X36 a_1339_74# a_225_74# a_1258_341# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X37 VPWR a_757_401# a_706_463# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
.ends

.subckt sky130_fd_sc_hs__nand2b_4 VNB VPB VPWR VGND A_N Y B a_31_74# a_243_74#
X0 VGND A_N a_31_74# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X1 a_243_74# B VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X2 a_243_74# a_31_74# Y VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X3 Y a_31_74# VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X4 VPWR B Y VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X5 a_243_74# B VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X6 VGND B a_243_74# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X7 VPWR A_N a_31_74# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X8 a_31_74# A_N VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X9 VGND B a_243_74# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X10 VPWR a_31_74# Y VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X11 Y B VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X12 a_243_74# a_31_74# Y VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X13 Y a_31_74# a_243_74# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X14 Y a_31_74# a_243_74# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
.ends

.subckt sky130_fd_sc_hs__or3b_2 VNB VPB VPWR VGND X A B C_N a_542_368# a_27_368# a_190_260#
+ a_458_368#
X0 a_190_260# a_27_368# VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1 X a_190_260# VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X2 a_542_368# B a_458_368# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 a_190_260# a_27_368# a_542_368# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 VGND B a_190_260# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X5 a_458_368# A VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 VGND C_N a_27_368# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=550000u l=150000u
X7 VGND a_190_260# X VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X8 VPWR a_190_260# X VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X9 X a_190_260# VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X10 a_190_260# A VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X11 VPWR C_N a_27_368# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
.ends

.subckt sky130_fd_sc_hs__nand4_1 VNB VPB VPWR VGND C Y D B A a_259_74# a_373_74# a_181_74#
X0 Y B VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X1 a_259_74# C a_181_74# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X2 a_181_74# D VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X3 Y A a_373_74# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X4 a_373_74# B a_259_74# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X5 VPWR C Y VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X6 Y D VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X7 VPWR A Y VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
.ends

.subckt sky130_fd_sc_hs__a31oi_2 VNB VPB VPWR VGND A2 A1 A3 Y B1 a_114_74# a_27_368#
+ a_200_74#
X0 VGND A3 a_114_74# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X1 Y A1 a_200_74# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X2 a_27_368# B1 Y VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X3 a_114_74# A3 VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X4 VPWR A2 a_27_368# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X5 Y B1 a_27_368# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X6 a_114_74# A2 a_200_74# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X7 a_200_74# A1 Y VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X8 a_200_74# A2 a_114_74# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X9 a_27_368# A1 VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X10 a_27_368# A2 VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X11 VPWR A1 a_27_368# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X12 Y B1 VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X13 VPWR A3 a_27_368# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X14 a_27_368# A3 VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
.ends

.subckt sky130_fd_sc_hs__nor2_4 VNB VPB VPWR VGND Y A B a_27_368#
X0 Y A VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X1 Y B a_27_368# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X2 Y B VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X3 VGND A Y VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X4 a_27_368# B Y VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X5 Y B a_27_368# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X6 a_27_368# A VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X7 VPWR A a_27_368# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X8 a_27_368# A VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X9 a_27_368# B Y VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X10 VGND B Y VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X11 VPWR A a_27_368# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
.ends

.subckt sky130_fd_sc_hs__nor4_1 VNB VPB VPWR VGND Y D C B A a_144_368# a_342_368#
+ a_228_368#
X0 VGND B Y VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X1 Y C VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X2 Y A VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X3 a_228_368# B a_144_368# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X4 a_144_368# A VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X5 a_342_368# C a_228_368# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X6 VGND D Y VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X7 Y D a_342_368# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
.ends

.subckt sky130_fd_sc_hs__nor2b_2 VNB VPB VPWR VGND A B_N Y a_27_392# a_228_368#
X0 a_228_368# A VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X1 VPWR A a_228_368# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X2 a_228_368# a_27_392# Y VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X3 VGND A Y VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X4 Y a_27_392# a_228_368# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X5 Y A VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X6 Y a_27_392# VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X7 VGND B_N a_27_392# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X8 VGND a_27_392# Y VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X9 VPWR B_N a_27_392# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_sc_hs__sdlclkp_1 VNB VPB VPWR VGND GCLK CLK GATE SCE a_114_112#
+ a_667_80# a_1166_94# a_288_48# a_722_492# a_1238_94# a_116_424# a_709_54# a_566_74#
+ a_318_74#
X0 a_114_112# GATE a_116_424# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X1 a_1238_94# CLK VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X2 GCLK a_1238_94# VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X3 a_709_54# a_566_74# VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X4 a_318_74# a_288_48# VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X5 VPWR CLK a_288_48# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X6 GCLK a_1238_94# VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X7 a_318_74# a_288_48# VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X8 VPWR a_709_54# a_722_492# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9 a_1166_94# CLK VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X10 a_116_424# SCE VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X11 a_722_492# a_288_48# a_566_74# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12 a_1238_94# a_709_54# a_1166_94# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X13 VGND CLK a_288_48# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X14 VGND GATE a_114_112# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=550000u l=150000u
X15 a_566_74# a_288_48# a_114_112# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=550000u l=150000u
X16 a_667_80# a_318_74# a_566_74# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17 a_114_112# SCE VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=550000u l=150000u
X18 a_709_54# a_566_74# VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X19 VGND a_709_54# a_667_80# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20 a_566_74# a_318_74# a_114_112# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X21 VPWR a_709_54# a_1238_94# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
.ends

.subckt fine_freq_track clk_out div_ratio_half[5] div_ratio_half[4] div_ratio_half[3]
+ div_ratio_half[2] div_ratio_half[1] div_ratio_half[0] ref_clk rst aux_osc_en fftl_en
+ fine_control_avg_window_select[4] fine_control_avg_window_select[3] fine_control_avg_window_select[2]
+ fine_control_avg_window_select[1] fine_control_avg_window_select[0] fine_con_step_size[3]
+ fine_con_step_size[2] fine_con_step_size[1] fine_con_step_size[0] manual_control_osc[12]
+ manual_control_osc[11] manual_control_osc[10] manual_control_osc[9] manual_control_osc[8]
+ manual_control_osc[7] manual_control_osc[6] manual_control_osc[5] manual_control_osc[4]
+ manual_control_osc[3] manual_control_osc[2] manual_control_osc[1] manual_control_osc[0]
+ aux_clk_out out_star osc_fine_con_final[12] osc_fine_con_final[11] osc_fine_con_final[10]
+ osc_fine_con_final[9] osc_fine_con_final[8] osc_fine_con_final[7] osc_fine_con_final[6]
+ osc_fine_con_final[5] osc_fine_con_final[4] osc_fine_con_final[3] osc_fine_con_final[2]
+ osc_fine_con_final[1] osc_fine_con_final[0] DVSS DVDD sky130_fd_sc_hs__dfrtp_4_9/a_1827_81#
+ sky130_fd_sc_hs__nor2b_1_23/Y sky130_fd_sc_hs__o21a_1_51/B1 sky130_fd_sc_hs__dfrbp_1_19/a_498_360#
+ sky130_fd_sc_hs__inv_4_65/Y sky130_fd_sc_hs__dfrtp_4_79/a_1350_392# sky130_fd_sc_hs__dfrtp_4_63/a_789_463#
+ sky130_fd_sc_hs__dfstp_2_4/a_2022_94# sky130_fd_sc_hs__nor2_1_35/B sky130_fd_sc_hs__dfstp_2_7/a_1278_74#
+ sky130_fd_sc_hs__nor2_1_3/a_116_368# sky130_fd_sc_hs__dfrbp_1_15/a_706_463# sky130_fd_sc_hs__inv_2_7/Y
+ sky130_fd_sc_hs__a22o_1_27/a_222_392# sky130_fd_sc_hs__a32oi_1_3/Y sky130_fd_sc_hs__a22o_1_21/a_52_123#
+ sky130_fd_sc_hs__dfrtp_4_3/a_37_78# sky130_fd_sc_hs__dfrtp_4_75/a_1678_395# sky130_fd_sc_hs__inv_4_45/A
+ sky130_fd_sc_hs__dfrtp_4_45/a_834_355# sky130_fd_sc_hs__dfrtp_4_37/a_1627_493# sky130_fd_sc_hs__dfrbp_1_45/a_319_360#
+ sky130_fd_sc_hs__fa_2_11/a_1205_79# sky130_fd_sc_hs__fa_2_1/CIN sky130_fd_sc_hs__nor2_1_31/Y
+ sky130_fd_sc_hs__a32oi_1_3/B1 sky130_fd_sc_hs__nand2_4_13/Y sky130_fd_sc_hs__nand3_1_1/a_155_74#
+ sky130_fd_sc_hs__nor2_1_37/B sky130_fd_sc_hs__dfrtp_4_59/a_313_74# sky130_fd_sc_hs__sdlclkp_1_1/a_114_112#
+ sky130_fd_sc_hs__nor2b_1_25/Y sky130_fd_sc_hs__o21a_1_7/A1 sky130_fd_sc_hs__sdlclkp_4_1/a_634_74#
+ sky130_fd_sc_hs__nor4_1_1/D sky130_fd_sc_hs__inv_4_63/Y sky130_fd_sc_hs__inv_4_125/A
+ sky130_fd_sc_hs__inv_4_59/A sky130_fd_sc_hs__dfxtp_2_3/a_1217_314# sky130_fd_sc_hs__dfrtp_4_25/a_313_74#
+ sky130_fd_sc_hs__clkbuf_8_1/X sky130_fd_sc_hs__inv_4_47/A sky130_fd_sc_hs__o21a_1_5/X
+ sky130_fd_sc_hs__o21a_1_37/a_376_387# sky130_fd_sc_hs__inv_4_55/Y sky130_fd_sc_hs__dfrtp_4_39/a_890_138#
+ sky130_fd_sc_hs__clkbuf_2_1/X sky130_fd_sc_hs__dfxtp_2_9/a_206_368# sky130_fd_sc_hs__xnor2_1_3/B
+ sky130_fd_sc_hs__nor2_1_61/B sky130_fd_sc_hs__dfrbp_1_25/a_125_78# sky130_fd_sc_hs__o21a_1_77/a_376_387#
+ sky130_fd_sc_hs__dfsbp_2_1/a_225_74# sky130_fd_sc_hs__nor2b_1_7/a_27_112# sky130_fd_sc_hs__dfrtn_1_7/a_714_127#
+ sky130_fd_sc_hs__o21a_1_77/a_83_244# sky130_fd_sc_hs__nand2_1_9/A sky130_fd_sc_hs__nand2_1_113/a_117_74#
+ sky130_fd_sc_hs__dfrbp_1_15/a_38_78# sky130_fd_sc_hs__inv_4_135/Y sky130_fd_sc_hs__nand4_2_1/B
+ sky130_fd_sc_hs__inv_4_73/A sky130_fd_sc_hs__nand2_1_47/B sky130_fd_sc_hs__nor2_1_43/a_116_368#
+ sky130_fd_sc_hs__a22oi_1_19/a_339_74# sky130_fd_sc_hs__dfrbp_1_5/a_1224_74# sky130_fd_sc_hs__xnor2_1_15/Y
+ sky130_fd_sc_hs__dfrbp_1_43/D sky130_fd_sc_hs__inv_4_137/A sky130_fd_sc_hs__dfstp_2_1/CLK
+ sky130_fd_sc_hs__nor2_1_41/Y sky130_fd_sc_hs__dfxtp_4_2/a_1141_508# sky130_fd_sc_hs__dfrtp_4_5/a_124_78#
+ sky130_fd_sc_hs__inv_4_103/A sky130_fd_sc_hs__dfrtn_1_23/D sky130_fd_sc_hs__nor2_1_45/B
+ sky130_fd_sc_hs__nor2b_1_45/a_27_112# sky130_fd_sc_hs__dfstp_2_7/Q sky130_fd_sc_hs__a31oi_2_1/Y
+ sky130_fd_sc_hs__dfrtp_4_81/a_699_463# sky130_fd_sc_hs__o22ai_1_9/B1 sky130_fd_sc_hs__xnor2_1_1/B
+ sky130_fd_sc_hs__nor2b_1_19/a_278_368# sky130_fd_sc_hs__nor3_1_5/Y sky130_fd_sc_hs__inv_4_87/Y
+ sky130_fd_sc_hs__nand2_1_77/a_117_74# sky130_fd_sc_hs__dfrbp_1_43/a_841_401# sky130_fd_sc_hs__o22ai_1_9/a_27_74#
+ sky130_fd_sc_hs__inv_4_133/Y sky130_fd_sc_hs__nor3_1_1/a_198_368# sky130_fd_sc_hs__o21a_1_71/A1
+ sky130_fd_sc_hs__a22o_1_3/a_222_392# sky130_fd_sc_hs__a21oi_1_97/Y sky130_fd_sc_hs__nor3_1_13/A
+ sky130_fd_sc_hs__inv_4_17/Y sky130_fd_sc_hs__nand2_1_43/a_117_74# sky130_fd_sc_hs__dfrtp_4_45/a_812_138#
+ sky130_fd_sc_hs__dfrtn_1_23/a_856_304# sky130_fd_sc_hs__o31ai_1_1/a_119_368# sky130_fd_sc_hs__fa_2_21/a_27_79#
+ sky130_fd_sc_hs__o211ai_1_7/a_311_74# sky130_fd_sc_hs__dfrtn_1_23/a_850_127# sky130_fd_sc_hs__nor3_1_13/C
+ sky130_fd_sc_hs__nand2_1_11/a_117_74# sky130_fd_sc_hs__dfrtn_1_17/a_33_74# sky130_fd_sc_hs__nand4_1_5/C
+ sky130_fd_sc_hs__dfrtp_4_29/a_1647_81# sky130_fd_sc_hs__fa_2_21/a_484_347# sky130_fd_sc_hs__dfxtp_2_3/a_695_459#
+ sky130_fd_sc_hs__dfrtp_4_81/a_124_78# sky130_fd_sc_hs__dfrbp_1_31/a_38_78# sky130_fd_sc_hs__dfrtp_4_67/a_1647_81#
+ sky130_fd_sc_hs__dfrbp_1_29/a_1224_74# sky130_fd_sc_hs__inv_4_75/A sky130_fd_sc_hs__dfrbp_1_5/a_38_78#
+ sky130_fd_sc_hs__nand2_1_5/a_117_74# sky130_fd_sc_hs__nor2_1_51/Y sky130_fd_sc_hs__dfrtn_1_41/a_507_368#
+ sky130_fd_sc_hs__or3b_2_1/a_458_368# sky130_fd_sc_hs__o21a_1_71/a_320_74# sky130_fd_sc_hs__a21oi_1_27/a_29_368#
+ sky130_fd_sc_hs__dfrbp_1_43/Q_N sky130_fd_sc_hs__nor2_1_37/Y sky130_fd_sc_hs__dfrtp_4_53/a_789_463#
+ sky130_fd_sc_hs__dfrbp_1_47/a_498_360# sky130_fd_sc_hs__dfstp_2_1/a_767_384# sky130_fd_sc_hs__dfrtn_1_49/a_1547_508#
+ sky130_fd_sc_hs__a22o_1_17/a_222_392# sky130_fd_sc_hs__dfrbp_1_35/Q_N sky130_fd_sc_hs__dfrtp_4_73/a_1678_395#
+ sky130_fd_sc_hs__dfrtp_4_35/a_834_355# sky130_fd_sc_hs__dfrtp_4_91/a_37_78# sky130_fd_sc_hs__fa_2_7/a_27_79#
+ sky130_fd_sc_hs__xnor2_1_7/Y sky130_fd_sc_hs__a21oi_1_9/a_29_368# sky130_fd_sc_hs__a21oi_1_71/a_29_368#
+ sky130_fd_sc_hs__xor2_1_5/a_455_87# sky130_fd_sc_hs__dfrbp_1_25/Q_N sky130_fd_sc_hs__dfrtp_4_43/D
+ sky130_fd_sc_hs__inv_4_85/Y sky130_fd_sc_hs__dfrtp_4_73/a_834_355# sky130_fd_sc_hs__dfrtn_1_39/a_922_127#
+ sky130_fd_sc_hs__dfrtp_4_27/a_1350_392# sky130_fd_sc_hs__dfrbp_1_21/D sky130_fd_sc_hs__maj3_1_3/a_598_384#
+ sky130_fd_sc_hs__nor2_1_47/B sky130_fd_sc_hs__o21a_1_15/A1 sky130_fd_sc_hs__inv_4_65/A
+ sky130_fd_sc_hs__dfrtn_1_33/a_33_74# sky130_fd_sc_hs__a22oi_1_15/Y sky130_fd_sc_hs__o21a_1_9/a_83_244#
+ sky130_fd_sc_hs__dfrtp_4_23/a_1678_395# sky130_fd_sc_hs__o21a_1_27/a_376_387# sky130_fd_sc_hs__dfrbp_1_41/a_2026_424#
+ sky130_fd_sc_hs__inv_4_37/A sky130_fd_sc_hs__dfrbp_1_23/a_832_118# sky130_fd_sc_hs__dfrtp_4_29/a_890_138#
+ sky130_fd_sc_hs__a22oi_1_21/Y sky130_fd_sc_hs__o21a_1_67/a_376_387# sky130_fd_sc_hs__maj3_1_1/a_595_136#
+ sky130_fd_sc_hs__or2_1_3/A sky130_fd_sc_hs__dfrbp_1_25/a_1465_471# sky130_fd_sc_hs__a21oi_1_17/Y
+ sky130_fd_sc_hs__inv_4_45/Y sky130_fd_sc_hs__nor3_1_5/A sky130_fd_sc_hs__dfrtp_4_67/a_890_138#
+ sky130_fd_sc_hs__dfrtn_1_13/D sky130_fd_sc_hs__xor2_1_11/B sky130_fd_sc_hs__o21a_1_35/X
+ sky130_fd_sc_hs__dfrtp_4_57/a_2010_409# sky130_fd_sc_hs__nor4_1_1/C sky130_fd_sc_hs__a21oi_1_57/a_117_74#
+ sky130_fd_sc_hs__or3b_2_1/B sky130_fd_sc_hs__dfrtn_1_37/a_817_508# sky130_fd_sc_hs__a211oi_1_1/Y
+ sky130_fd_sc_hs__nor2_1_97/A sky130_fd_sc_hs__inv_4_79/Y sky130_fd_sc_hs__dfxtp_4_9/a_27_74#
+ sky130_fd_sc_hs__dfrbp_1_41/a_910_118# sky130_fd_sc_hs__nor2_1_33/a_116_368# sky130_fd_sc_hs__inv_4_43/Y
+ sky130_fd_sc_hs__nor2_1_71/a_116_368# sky130_fd_sc_hs__nand2_2_3/A sky130_fd_sc_hs__dfrtp_4_7/a_699_463#
+ sky130_fd_sc_hs__nand2_2_3/a_27_74# sky130_fd_sc_hs__inv_4_41/Y sky130_fd_sc_hs__o21ai_2_1/B1
+ sky130_fd_sc_hs__a31oi_2_1/A1 sky130_fd_sc_hs__dfrtp_4_71/a_699_463# sky130_fd_sc_hs__dfrtn_1_31/a_300_74#
+ sky130_fd_sc_hs__dfrtp_4_59/D sky130_fd_sc_hs__a21oi_1_105/a_29_368# sky130_fd_sc_hs__dfrtp_4_73/a_313_74#
+ sky130_fd_sc_hs__nor2_1_87/Y sky130_fd_sc_hs__nand2_1_117/a_117_74# sky130_fd_sc_hs__dfrbp_1_37/a_1624_74#
+ sky130_fd_sc_hs__dfrbp_1_1/a_319_360# sky130_fd_sc_hs__nor3_1_9/Y sky130_fd_sc_hs__inv_4_129/A
+ sky130_fd_sc_hs__dfstp_2_5/a_27_74# sky130_fd_sc_hs__dfrtn_1_3/a_1736_119# sky130_fd_sc_hs__dfrtp_4_35/a_812_138#
+ sky130_fd_sc_hs__dfrtp_4_41/a_313_74# sky130_fd_sc_hs__inv_4_69/A sky130_fd_sc_hs__dfrbp_1_37/D
+ sky130_fd_sc_hs__inv_4_129/Y sky130_fd_sc_hs__dfrtn_1_3/a_1266_119# sky130_fd_sc_hs__dfrtp_4_73/a_812_138#
+ sky130_fd_sc_hs__nor2_1_35/Y sky130_fd_sc_hs__fa_2_3/a_27_378# sky130_fd_sc_hs__o21a_1_15/a_83_244#
+ sky130_fd_sc_hs__or2_1_1/A sky130_fd_sc_hs__dfrtp_4_9/a_124_78# sky130_fd_sc_hs__xor2_1_9/A
+ sky130_fd_sc_hs__inv_4_77/Y sky130_fd_sc_hs__dfrtp_4_19/a_1647_81# sky130_fd_sc_hs__maj3_1_1/A
+ sky130_fd_sc_hs__dfrtp_4_87/a_1627_493# sky130_fd_sc_hs__o21a_1_23/A1 sky130_fd_sc_hs__nor4_1_3/Y
+ sky130_fd_sc_hs__nor2_2_1/Y sky130_fd_sc_hs__inv_4_55/A sky130_fd_sc_hs__dfrtp_4_45/a_37_78#
+ sky130_fd_sc_hs__inv_4_113/Y sky130_fd_sc_hs__maj3_1_3/A sky130_fd_sc_hs__dfrbp_1_19/a_1224_74#
+ sky130_fd_sc_hs__fa_2_3/CIN sky130_fd_sc_hs__dfrtn_1_31/a_507_368# sky130_fd_sc_hs__dfrtp_4_77/a_1350_392#
+ sky130_fd_sc_hs__nor4_1_1/a_342_368# sky130_fd_sc_hs__o21a_1_65/B1 sky130_fd_sc_hs__xor2_1_11/a_455_87#
+ sky130_fd_sc_hs__xor2_1_9/a_158_392# sky130_fd_sc_hs__dfrtn_1_47/a_1547_508# sky130_fd_sc_hs__dfrtp_4_83/a_789_463#
+ sky130_fd_sc_hs__a22oi_1_5/Y sky130_fd_sc_hs__inv_4_11/A sky130_fd_sc_hs__nand2_1_15/a_117_74#
+ sky130_fd_sc_hs__dfrbp_1_35/a_706_463# sky130_fd_sc_hs__dfrbp_1_25/a_319_360# sky130_fd_sc_hs__inv_4_49/Y
+ sky130_fd_sc_hs__dfrtp_4_63/a_834_355# sky130_fd_sc_hs__dfrtp_4_49/a_494_366# sky130_fd_sc_hs__dfrtp_4_85/a_124_78#
+ sky130_fd_sc_hs__and2_2_5/a_31_74# sky130_fd_sc_hs__dfrtn_1_7/a_1934_94# sky130_fd_sc_hs__nand2_4_9/Y
+ sky130_fd_sc_hs__fa_2_3/a_701_79# sky130_fd_sc_hs__dfrtn_1_29/a_922_127# sky130_fd_sc_hs__dfrtn_1_9/a_1598_93#
+ sky130_fd_sc_hs__dfrtp_4_25/a_1350_392# sky130_fd_sc_hs__dfrtp_4_89/a_494_366# sky130_fd_sc_hs__dfrtn_1_7/D
+ sky130_fd_sc_hs__o211ai_1_9/a_116_368# sky130_fd_sc_hs__o21a_1_75/a_320_74# sky130_fd_sc_hs__nor2_1_31/B
+ sky130_fd_sc_hs__fa_2_11/SUM sky130_fd_sc_hs__dfxtp_2_1/a_1217_314# sky130_fd_sc_hs__dfrbp_1_43/a_1434_74#
+ sky130_fd_sc_hs__xnor2_1_3/A sky130_fd_sc_hs__dfrbp_1_3/a_1624_74# sky130_fd_sc_hs__dfxtp_4_3/a_206_368#
+ sky130_fd_sc_hs__nor2_1_27/B sky130_fd_sc_hs__a22o_1_29/X sky130_fd_sc_hs__dfrtp_4_21/a_1678_395#
+ sky130_fd_sc_hs__xnor2_1_3/a_112_119# sky130_fd_sc_hs__dfrbp_1_13/a_832_118# sky130_fd_sc_hs__dfrtp_4_19/a_890_138#
+ sky130_fd_sc_hs__a21oi_1_75/a_29_368# sky130_fd_sc_hs__xor2_1_9/a_455_87# sky130_fd_sc_hs__o21a_1_57/a_376_387#
+ sky130_fd_sc_hs__a31oi_2_1/a_200_74# sky130_fd_sc_hs__inv_4_63/A sky130_fd_sc_hs__xor2_1_9/X
+ sky130_fd_sc_hs__o21a_1_65/X sky130_fd_sc_hs__a32oi_1_7/B1 sky130_fd_sc_hs__fa_2_5/a_992_347#
+ sky130_fd_sc_hs__or2_1_3/X sky130_fd_sc_hs__dfxtp_4_5/a_696_458# sky130_fd_sc_hs__nor2_1_7/Y
+ sky130_fd_sc_hs__o21ai_1_3/B1 sky130_fd_sc_hs__inv_2_1/A sky130_fd_sc_hs__nor2_1_23/a_116_368#
+ sky130_fd_sc_hs__o21a_1_3/a_376_387# sky130_fd_sc_hs__dfrtp_4_21/a_699_463# sky130_fd_sc_hs__nor2b_1_5/a_278_368#
+ sky130_fd_sc_hs__dfrtp_4_7/D sky130_fd_sc_hs__nand2_4_9/a_27_74# sky130_fd_sc_hs__o21a_1_73/A2
+ sky130_fd_sc_hs__dfrtp_4_61/a_699_463# sky130_fd_sc_hs__dfrtn_1_37/a_1550_119# sky130_fd_sc_hs__nor2_1_107/a_116_368#
+ sky130_fd_sc_hs__nor2_1_65/Y sky130_fd_sc_hs__dfrbp_1_23/a_841_401# sky130_fd_sc_hs__nand2_1_59/Y
+ sky130_fd_sc_hs__fa_2_15/a_336_347# sky130_fd_sc_hs__nor2_1_63/B sky130_fd_sc_hs__dfrtn_1_1/a_1736_119#
+ sky130_fd_sc_hs__inv_4_3/A sky130_fd_sc_hs__inv_4_105/A sky130_fd_sc_hs__dfxtp_2_9/a_708_101#
+ sky130_fd_sc_hs__dfrtn_1_1/a_1266_119# sky130_fd_sc_hs__dfrtp_4_63/a_812_138# sky130_fd_sc_hs__nor2_1_25/B
+ sky130_fd_sc_hs__dfrtn_1_41/a_856_304# sky130_fd_sc_hs__a32oi_1_9/Y sky130_fd_sc_hs__o21a_1_25/A1
+ sky130_fd_sc_hs__fa_2_15/a_27_79# sky130_fd_sc_hs__o21a_1_27/X sky130_fd_sc_hs__dfrtn_1_41/a_850_127#
+ sky130_fd_sc_hs__o31ai_1_1/B1 sky130_fd_sc_hs__a21oi_1_109/a_29_368# sky130_fd_sc_hs__dfrbp_1_7/a_125_78#
+ sky130_fd_sc_hs__inv_4_81/Y sky130_fd_sc_hs__o22ai_1_11/a_340_368# sky130_fd_sc_hs__fa_2_7/a_683_347#
+ sky130_fd_sc_hs__dfrtp_4_47/a_1647_81# sky130_fd_sc_hs__o22ai_1_1/a_340_368# sky130_fd_sc_hs__fa_2_19/CIN
+ sky130_fd_sc_hs__dfrtp_4_43/a_1827_81# sky130_fd_sc_hs__dfrtn_1_21/a_507_368# sky130_fd_sc_hs__dfrtp_4_87/a_1647_81#
+ sky130_fd_sc_hs__dfrbp_1_47/a_1224_74# sky130_fd_sc_hs__dfxtp_4_7/D sky130_fd_sc_hs__dfrtp_4_45/a_313_74#
+ sky130_fd_sc_hs__dfrtp_4_9/a_789_463# sky130_fd_sc_hs__dfrbp_1_27/a_498_360# sky130_fd_sc_hs__nor3_1_11/a_114_368#
+ sky130_fd_sc_hs__nor2_1_27/Y sky130_fd_sc_hs__xnor2_1_11/a_112_119# sky130_fd_sc_hs__a222oi_1_3/a_116_392#
+ sky130_fd_sc_hs__xnor2_1_1/A sky130_fd_sc_hs__fa_2_7/a_27_378# sky130_fd_sc_hs__o21a_1_19/a_83_244#
+ sky130_fd_sc_hs__dfrtp_4_35/a_1627_493# sky130_fd_sc_hs__dfrbp_1_15/a_319_360# sky130_fd_sc_hs__maj3_1_1/C
+ sky130_fd_sc_hs__clkbuf_8_1/A sky130_fd_sc_hs__nor2_1_17/Y sky130_fd_sc_hs__a21oi_1_121/a_29_368#
+ sky130_fd_sc_hs__fa_2_17/a_683_347# sky130_fd_sc_hs__dfrtp_4_53/a_834_355# sky130_fd_sc_hs__maj3_1_3/B
+ sky130_fd_sc_hs__dfrtp_4_85/a_37_78# sky130_fd_sc_hs__nor3_1_3/A sky130_fd_sc_hs__nor4_1_1/a_144_368#
+ sky130_fd_sc_hs__fa_2_21/a_1205_79# sky130_fd_sc_hs__o21a_1_59/A1 sky130_fd_sc_hs__o21ai_1_7/a_162_368#
+ sky130_fd_sc_hs__dfrtn_1_19/a_922_127# sky130_fd_sc_hs__o21a_1_63/a_83_244# sky130_fd_sc_hs__dfrtp_4_79/a_494_366#
+ sky130_fd_sc_hs__maj3_1_1/a_223_120# sky130_fd_sc_hs__inv_4_79/A sky130_fd_sc_hs__inv_4_21/Y
+ sky130_fd_sc_hs__nand4_1_3/a_373_74# sky130_fd_sc_hs__fa_2_21/a_487_79# sky130_fd_sc_hs__nor2_1_9/Y
+ sky130_fd_sc_hs__inv_4_13/A sky130_fd_sc_hs__nand2_1_19/a_117_74# sky130_fd_sc_hs__dfstp_2_1/a_612_74#
+ sky130_fd_sc_hs__nor3_1_1/Y sky130_fd_sc_hs__o21a_1_47/a_376_387# sky130_fd_sc_hs__o21ai_1_3/a_27_74#
+ sky130_fd_sc_hs__inv_4_125/Y sky130_fd_sc_hs__dfxtp_4_3/a_437_503# sky130_fd_sc_hs__dfrbp_1_23/a_1465_471#
+ sky130_fd_sc_hs__dfrtp_4_47/a_890_138# sky130_fd_sc_hs__dfrtp_4_89/a_124_78# sky130_fd_sc_hs__nor2b_1_31/a_27_112#
+ sky130_fd_sc_hs__nor2_4_1/B sky130_fd_sc_hs__dfrtp_4_55/a_2010_409# sky130_fd_sc_hs__fa_2_7/a_701_79#
+ sky130_fd_sc_hs__dfrtp_4_87/a_890_138# sky130_fd_sc_hs__nor3_1_9/B sky130_fd_sc_hs__o21a_1_73/B1
+ sky130_fd_sc_hs__dfrtn_1_37/D sky130_fd_sc_hs__nor2_1_13/a_116_368# sky130_fd_sc_hs__nor4_1_3/B
+ sky130_fd_sc_hs__or3b_2_1/X sky130_fd_sc_hs__nor3_1_11/B sky130_fd_sc_hs__inv_4_39/A
+ sky130_fd_sc_hs__nor2_1_83/B sky130_fd_sc_hs__dfrtp_4_23/a_124_78# sky130_fd_sc_hs__dfsbp_2_1/a_2221_74#
+ sky130_fd_sc_hs__fa_2_19/SUM sky130_fd_sc_hs__nor2b_1_7/Y sky130_fd_sc_hs__dfrtp_4_51/a_699_463#
+ sky130_fd_sc_hs__nor2_1_91/a_116_368# sky130_fd_sc_hs__inv_4_67/Y sky130_fd_sc_hs__nand2_4_7/Y
+ sky130_fd_sc_hs__dfrbp_1_13/a_841_401# sky130_fd_sc_hs__a32oi_1_7/A1 sky130_fd_sc_hs__a22o_1_13/a_132_392#
+ sky130_fd_sc_hs__o31ai_1_1/a_203_368# sky130_fd_sc_hs__o21a_1_75/B1 sky130_fd_sc_hs__dfrbp_1_3/D
+ sky130_fd_sc_hs__nor2_1_45/Y sky130_fd_sc_hs__a21oi_1_13/a_29_368# sky130_fd_sc_hs__dfrtn_1_41/a_33_74#
+ sky130_fd_sc_hs__dfrtp_4_53/a_812_138# sky130_fd_sc_hs__dfrtn_1_31/a_856_304# sky130_fd_sc_hs__nor2_1_5/Y
+ sky130_fd_sc_hs__nor4_1_1/a_228_368# sky130_fd_sc_hs__dfrtn_1_31/a_850_127# sky130_fd_sc_hs__nor3_1_1/B
+ sky130_fd_sc_hs__dfrtp_4_85/a_1627_493# sky130_fd_sc_hs__or3b_2_1/a_542_368# sky130_fd_sc_hs__o21a_1_53/B1
+ sky130_fd_sc_hs__dfrtp_4_37/a_1647_81# sky130_fd_sc_hs__dfrtp_4_3/a_1647_81# sky130_fd_sc_hs__dfrtp_4_33/a_1827_81#
+ sky130_fd_sc_hs__dfrtn_1_39/a_714_127# sky130_fd_sc_hs__dfrtn_1_11/a_507_368# sky130_fd_sc_hs__dfrtp_4_77/a_1647_81#
+ sky130_fd_sc_hs__dfrtp_4_39/a_37_78# sky130_fd_sc_hs__inv_2_5/Y sky130_fd_sc_hs__dfrtp_4_75/a_1350_392#
+ sky130_fd_sc_hs__a32oi_1_1/Y sky130_fd_sc_hs__dfrbp_1_17/a_498_360# sky130_fd_sc_hs__fa_2_11/B
+ sky130_fd_sc_hs__dfrbp_1_31/a_796_463# sky130_fd_sc_hs__o211ai_1_3/Y sky130_fd_sc_hs__nor2_1_25/Y
+ sky130_fd_sc_hs__dfstp_2_1/a_2022_94# sky130_fd_sc_hs__o22ai_1_11/a_142_368# sky130_fd_sc_hs__o22ai_1_1/a_142_368#
+ sky130_fd_sc_hs__nor2_1_1/a_116_368# sky130_fd_sc_hs__dfrtp_4_71/a_1678_395# sky130_fd_sc_hs__dfrtn_1_39/a_300_74#
+ sky130_fd_sc_hs__nor2_1_87/B sky130_fd_sc_hs__fa_2_13/B sky130_fd_sc_hs__dfrtp_4_83/a_834_355#
+ sky130_fd_sc_hs__dfrtp_4_69/a_494_366# sky130_fd_sc_hs__a21oi_1_1/Y sky130_fd_sc_hs__inv_4_53/Y
+ sky130_fd_sc_hs__dfrtn_1_49/a_922_127# sky130_fd_sc_hs__dfrbp_1_23/a_1434_74# sky130_fd_sc_hs__a21oi_1_43/a_117_74#
+ sky130_fd_sc_hs__o22ai_1_1/Y sky130_fd_sc_hs__a32oi_1_3/a_469_74# sky130_fd_sc_hs__dfrtp_4_15/a_313_74#
+ sky130_fd_sc_hs__dfxtp_4_9/CLK sky130_fd_sc_hs__dfrtp_4_39/a_1678_395# sky130_fd_sc_hs__dfrbp_1_33/a_832_118#
+ sky130_fd_sc_hs__dfrtp_4_37/a_890_138# sky130_fd_sc_hs__dfxtp_2_7/a_206_368# sky130_fd_sc_hs__dfrtp_4_53/a_37_78#
+ sky130_fd_sc_hs__dfrbp_1_15/a_125_78# sky130_fd_sc_hs__dfrtp_4_3/a_890_138# sky130_fd_sc_hs__inv_4_87/A
+ sky130_fd_sc_hs__dfrtp_4_53/a_2010_409# sky130_fd_sc_hs__dfrtp_4_77/a_890_138# sky130_fd_sc_hs__o21a_1_67/a_83_244#
+ sky130_fd_sc_hs__nand4_2_1/C sky130_fd_sc_hs__inv_4_59/Y sky130_fd_sc_hs__dfrbp_1_41/D
+ sky130_fd_sc_hs__nand2_2_1/Y sky130_fd_sc_hs__nand2_1_103/a_117_74# sky130_fd_sc_hs__o21a_1_63/A1
+ sky130_fd_sc_hs__maj3_1_1/B sky130_fd_sc_hs__fa_2_3/B sky130_fd_sc_hs__nor2_1_41/a_116_368#
+ sky130_fd_sc_hs__dfrbp_1_7/a_796_463# sky130_fd_sc_hs__dfsbp_2_1/a_1339_74# sky130_fd_sc_hs__o21a_1_67/B1
+ sky130_fd_sc_hs__dfrtp_4_41/a_699_463# sky130_fd_sc_hs__nand2_1_99/a_117_74# sky130_fd_sc_hs__nor2_1_81/a_116_368#
+ sky130_fd_sc_hs__dfrtn_1_35/a_1550_119# sky130_fd_sc_hs__dfrtp_4_5/a_37_78# sky130_fd_sc_hs__nor2_4_3/a_27_368#
+ sky130_fd_sc_hs__dfrbp_1_29/Q_N sky130_fd_sc_hs__nand2_1_67/a_117_74# sky130_fd_sc_hs__o21a_1_59/X
+ sky130_fd_sc_hs__dfrbp_1_45/a_1624_74# sky130_fd_sc_hs__nor2_1_29/Y sky130_fd_sc_hs__or2_1_3/B
+ sky130_fd_sc_hs__xnor2_1_5/B sky130_fd_sc_hs__dfrtp_4_27/a_124_78# sky130_fd_sc_hs__dfrtn_1_21/a_856_304#
+ sky130_fd_sc_hs__fa_2_15/B sky130_fd_sc_hs__dfxtp_2_5/a_431_508# sky130_fd_sc_hs__dfrtp_4_83/a_812_138#
+ sky130_fd_sc_hs__dfrtn_1_21/a_850_127# sky130_fd_sc_hs__a22oi_1_3/a_159_74# sky130_fd_sc_hs__o21a_1_17/a_320_74#
+ sky130_fd_sc_hs__inv_4_33/Y sky130_fd_sc_hs__xnor2_1_3/a_138_385# sky130_fd_sc_hs__nand3_1_1/A
+ sky130_fd_sc_hs__dfrtp_4_23/a_1827_81# sky130_fd_sc_hs__a21oi_1_49/a_29_368# sky130_fd_sc_hs__dfrtn_1_29/a_714_127#
+ sky130_fd_sc_hs__dfrtn_1_3/D sky130_fd_sc_hs__dfrtp_4_71/a_124_78# sky130_fd_sc_hs__dfrbp_1_9/a_832_118#
+ sky130_fd_sc_hs__dfrbp_1_27/a_1224_74# sky130_fd_sc_hs__dfrtp_4_73/a_1350_392# sky130_fd_sc_hs__nor2_1_99/Y
+ sky130_fd_sc_hs__o21a_1_61/a_320_74# sky130_fd_sc_hs__a21oi_1_17/a_29_368# sky130_fd_sc_hs__dfrbp_1_21/a_796_463#
+ sky130_fd_sc_hs__dfrbp_1_19/a_38_78# sky130_fd_sc_hs__dfrtn_1_45/a_1547_508# sky130_fd_sc_hs__o21a_1_17/X
+ sky130_fd_sc_hs__inv_4_83/Y sky130_fd_sc_hs__dfrtp_4_33/a_1627_493# sky130_fd_sc_hs__inv_4_61/A
+ sky130_fd_sc_hs__dfrtp_4_31/D sky130_fd_sc_hs__xnor2_1_13/A sky130_fd_sc_hs__dfrbp_1_43/a_706_463#
+ sky130_fd_sc_hs__dfrbp_1_35/a_319_360# sky130_fd_sc_hs__dfrtp_4_9/a_834_355# sky130_fd_sc_hs__dfrtp_4_89/a_1678_395#
+ sky130_fd_sc_hs__fa_2_11/a_27_378# sky130_fd_sc_hs__a21oi_1_61/a_29_368# sky130_fd_sc_hs__dfrtp_4_23/a_1350_392#
+ sky130_fd_sc_hs__dfrtp_4_59/a_494_366# sky130_fd_sc_hs__dfrtp_4_79/a_37_78# sky130_fd_sc_hs__dfrbp_1_13/a_1434_74#
+ sky130_fd_sc_hs__maj3_1_1/a_598_384# sky130_fd_sc_hs__and2_2_5/X sky130_fd_sc_hs__o21a_1_17/A1
+ sky130_fd_sc_hs__dfrbp_1_39/a_1482_48# sky130_fd_sc_hs__fa_2_3/A sky130_fd_sc_hs__dfrtp_4_37/a_1678_395#
+ sky130_fd_sc_hs__o22ai_1_7/A1 sky130_fd_sc_hs__nor3_1_15/A sky130_fd_sc_hs__fa_2_21/CIN
+ sky130_fd_sc_hs__a21oi_1_79/a_117_74# sky130_fd_sc_hs__fa_2_19/B sky130_fd_sc_hs__dfxtp_4_5/a_544_485#
+ sky130_fd_sc_hs__dfrbp_1_7/a_38_78# sky130_fd_sc_hs__dfrtn_1_27/a_120_74# sky130_fd_sc_hs__nand2_2_1/B
+ sky130_fd_sc_hs__a21oi_1_47/a_117_74# sky130_fd_sc_hs__o21a_1_33/X sky130_fd_sc_hs__inv_4_25/A
+ sky130_fd_sc_hs__fa_2_11/a_701_79# sky130_fd_sc_hs__a32oi_1_7/a_469_74# sky130_fd_sc_hs__dfrtp_4_31/a_699_463#
+ sky130_fd_sc_hs__xnor2_1_11/a_138_385# sky130_fd_sc_hs__a21oi_1_91/a_117_74# sky130_fd_sc_hs__dfrtp_4_23/a_37_78#
+ sky130_fd_sc_hs__dfrtn_1_21/a_300_74# sky130_fd_sc_hs__nor2_1_117/a_116_368# sky130_fd_sc_hs__dfrbp_1_7/Q
+ sky130_fd_sc_hs__a211oi_1_1/a_159_74# sky130_fd_sc_hs__dfxtp_4_3/a_27_74# sky130_fd_sc_hs__dfrtp_4_63/a_313_74#
+ sky130_fd_sc_hs__dfrbp_1_33/a_841_401# sky130_fd_sc_hs__o21a_1_63/X sky130_fd_sc_hs__o21a_1_63/A2
+ sky130_fd_sc_hs__nand2_1_107/a_117_74# sky130_fd_sc_hs__nor2_1_33/Y sky130_fd_sc_hs__dfrtn_1_39/a_1934_94#
+ sky130_fd_sc_hs__xnor2_1_1/a_376_368# sky130_fd_sc_hs__nor2b_1_47/a_278_368# sky130_fd_sc_hs__dfrtn_1_1/a_120_74#
+ sky130_fd_sc_hs__inv_2_3/A sky130_fd_sc_hs__nand4_1_5/A sky130_fd_sc_hs__o21a_1_37/a_83_244#
+ sky130_fd_sc_hs__dfrtp_4_31/a_313_74# sky130_fd_sc_hs__dfrtp_4_9/a_812_138# sky130_fd_sc_hs__nor2_1_7/B
+ sky130_fd_sc_hs__nand4_1_1/C sky130_fd_sc_hs__dfrtn_1_11/a_856_304# sky130_fd_sc_hs__inv_4_123/Y
+ sky130_fd_sc_hs__o21a_1_71/B1 sky130_fd_sc_hs__dfrtn_1_11/a_850_127# sky130_fd_sc_hs__dfrtp_4_83/a_1627_493#
+ sky130_fd_sc_hs__dfrbp_1_31/a_125_78# sky130_fd_sc_hs__nor2b_1_19/Y sky130_fd_sc_hs__dfrtp_4_17/a_1647_81#
+ sky130_fd_sc_hs__fa_2_5/a_1119_79# sky130_fd_sc_hs__dfrtp_4_13/a_1827_81# sky130_fd_sc_hs__dfrtn_1_9/a_1547_508#
+ sky130_fd_sc_hs__dfrtn_1_19/a_714_127# sky130_fd_sc_hs__dfrtp_4_57/a_1647_81# sky130_fd_sc_hs__dfrbp_1_17/a_1224_74#
+ sky130_fd_sc_hs__inv_4_19/A sky130_fd_sc_hs__dfrbp_1_1/Q_N sky130_fd_sc_hs__dfrtp_4_9/a_2010_409#
+ sky130_fd_sc_hs__nor2_1_57/Y sky130_fd_sc_hs__dfrtn_1_3/a_817_508# sky130_fd_sc_hs__dfrbp_1_11/a_796_463#
+ sky130_fd_sc_hs__fa_2_9/SUM sky130_fd_sc_hs__dfrtp_4_43/a_789_463# sky130_fd_sc_hs__o22ai_1_9/Y
+ sky130_fd_sc_hs__dfrtp_4_91/a_1827_81# sky130_fd_sc_hs__dfrbp_1_37/a_498_360# sky130_fd_sc_hs__nor2b_2_1/Y
+ sky130_fd_sc_hs__nor3_1_3/Y sky130_fd_sc_hs__xor2_1_7/a_158_392# sky130_fd_sc_hs__a22oi_1_7/a_159_74#
+ sky130_fd_sc_hs__nand2_2_5/a_27_74# sky130_fd_sc_hs__nor2_1_69/B sky130_fd_sc_hs__o21ai_1_3/Y
+ sky130_fd_sc_hs__nor2_1_5/B sky130_fd_sc_hs__nand3_1_1/B sky130_fd_sc_hs__dfrtn_1_41/D
+ sky130_fd_sc_hs__dfrtp_4_21/a_1350_392# sky130_fd_sc_hs__dfrtp_4_75/a_124_78# sky130_fd_sc_hs__inv_4_41/A
+ sky130_fd_sc_hs__fa_2_5/SUM sky130_fd_sc_hs__o21a_1_27/A1 sky130_fd_sc_hs__nor2_1_99/A
+ sky130_fd_sc_hs__dfrtn_1_7/a_1598_93# sky130_fd_sc_hs__o21a_1_65/a_320_74# sky130_fd_sc_hs__dfrbp_1_9/a_841_401#
+ sky130_fd_sc_hs__a22oi_1_1/a_339_74# sky130_fd_sc_hs__fa_2_23/B sky130_fd_sc_hs__dfrbp_1_1/a_1624_74#
+ sky130_fd_sc_hs__dfxtp_4_2/a_206_368# sky130_fd_sc_hs__sdlclkp_4_1/a_1292_74# sky130_fd_sc_hs__o21a_1_17/a_376_387#
+ sky130_fd_sc_hs__dfrbp_1_21/a_1465_471# sky130_fd_sc_hs__dfrtp_4_17/a_890_138# sky130_fd_sc_hs__a21oi_1_65/a_29_368#
+ sky130_fd_sc_hs__or2_1_1/X sky130_fd_sc_hs__dfrbp_1_39/a_1465_471# sky130_fd_sc_hs__dfrtp_4_57/a_890_138#
+ sky130_fd_sc_hs__dfrtp_4_47/a_37_78# sky130_fd_sc_hs__dfrtn_1_9/a_507_368# sky130_fd_sc_hs__fa_2_3/a_336_347#
+ sky130_fd_sc_hs__inv_4_29/A sky130_fd_sc_hs__nand2_2_5/B sky130_fd_sc_hs__o21a_1_3/A1
+ sky130_fd_sc_hs__dfstp_2_5/a_1566_92# sky130_fd_sc_hs__nor4_1_1/A sky130_fd_sc_hs__nand4_2_1/a_304_74#
+ sky130_fd_sc_hs__nor2_1_21/Y sky130_fd_sc_hs__dfrbp_1_31/a_910_118# sky130_fd_sc_hs__a32oi_1_1/a_391_74#
+ sky130_fd_sc_hs__maj3_1_3/C sky130_fd_sc_hs__nor2_1_63/Y sky130_fd_sc_hs__inv_4_91/A
+ sky130_fd_sc_hs__nor2_1_61/a_116_368# sky130_fd_sc_hs__dfrtn_1_33/a_1550_119# sky130_fd_sc_hs__nor2b_1_3/a_278_368#
+ sky130_fd_sc_hs__fa_2_9/B sky130_fd_sc_hs__dfrbp_1_3/a_498_360# sky130_fd_sc_hs__nor3_1_9/C
+ sky130_fd_sc_hs__nor2_1_73/Y sky130_fd_sc_hs__o31ai_1_3/a_114_74# sky130_fd_sc_hs__inv_4_109/A
+ sky130_fd_sc_hs__a22o_1_23/a_132_392# sky130_fd_sc_hs__fa_2_5/CIN sky130_fd_sc_hs__inv_4_39/Y
+ sky130_fd_sc_hs__dfrtn_1_29/a_1934_94# sky130_fd_sc_hs__dfrbp_1_25/a_1624_74# sky130_fd_sc_hs__fa_2_15/a_992_347#
+ sky130_fd_sc_hs__nor2b_1_37/a_278_368# sky130_fd_sc_hs__dfxtp_2_7/a_708_101# sky130_fd_sc_hs__a21oi_1_95/a_117_74#
+ sky130_fd_sc_hs__dfxtp_4_5/D sky130_fd_sc_hs__dfrtn_1_7/a_1547_508# sky130_fd_sc_hs__dfrtp_4_67/a_313_74#
+ sky130_fd_sc_hs__xnor2_1_5/Y sky130_fd_sc_hs__nand2_1_89/Y sky130_fd_sc_hs__dfrtn_1_43/a_120_74#
+ sky130_fd_sc_hs__dfrtn_1_49/a_714_127# sky130_fd_sc_hs__o31ai_1_3/Y sky130_fd_sc_hs__dfrtn_1_43/a_1547_508#
+ sky130_fd_sc_hs__dfrtp_4_35/a_313_74# sky130_fd_sc_hs__dfrbp_1_9/a_2026_424# sky130_fd_sc_hs__dfrtp_4_33/a_789_463#
+ sky130_fd_sc_hs__o21a_1_1/A1 sky130_fd_sc_hs__nand4_1_1/D sky130_fd_sc_hs__dfrtp_4_81/a_1827_81#
+ sky130_fd_sc_hs__xor2_1_5/a_355_368# sky130_fd_sc_hs__inv_2_5/A sky130_fd_sc_hs__dfrtp_4_31/a_1627_493#
+ sky130_fd_sc_hs__inv_4_99/A sky130_fd_sc_hs__dfrbp_1_7/a_910_118# sky130_fd_sc_hs__dfrbp_1_35/a_125_78#
+ sky130_fd_sc_hs__o21a_1_25/X sky130_fd_sc_hs__dfrbp_1_23/a_706_463# sky130_fd_sc_hs__dfrtp_4_87/a_1678_395#
+ sky130_fd_sc_hs__dfrtp_4_49/a_1627_493# sky130_fd_sc_hs__a21oi_1_111/a_29_368# sky130_fd_sc_hs__inv_4_89/Y
+ sky130_fd_sc_hs__dfrtn_1_19/a_1736_119# sky130_fd_sc_hs__dfrtp_4_39/a_494_366# sky130_fd_sc_hs__dfrtn_1_19/a_1266_119#
+ sky130_fd_sc_hs__o21a_1_53/a_83_244# sky130_fd_sc_hs__inv_4_23/A sky130_fd_sc_hs__o21a_1_61/A2
+ sky130_fd_sc_hs__o21a_1_59/A2 sky130_fd_sc_hs__inv_4_117/Y sky130_fd_sc_hs__o21ai_1_11/Y
+ sky130_fd_sc_hs__dfrbp_1_33/a_1434_74# sky130_fd_sc_hs__nor2_1_49/Y sky130_fd_sc_hs__fa_2_17/a_27_79#
+ sky130_fd_sc_hs__nor3_1_13/B sky130_fd_sc_hs__nand3_1_1/C sky130_fd_sc_hs__xnor2_1_9/Y
+ sky130_fd_sc_hs__dfxtp_4_2/a_437_503# sky130_fd_sc_hs__dfrtp_4_51/a_2010_409# sky130_fd_sc_hs__dfrbp_1_41/a_832_118#
+ sky130_fd_sc_hs__dfrtp_4_79/a_124_78# sky130_fd_sc_hs__nor2b_1_21/a_27_112# sky130_fd_sc_hs__nor2_1_99/B
+ sky130_fd_sc_hs__o21a_1_75/A2 sky130_fd_sc_hs__nand2_1_53/a_117_74# sky130_fd_sc_hs__o21a_1_69/a_320_74#
+ sky130_fd_sc_hs__dfrbp_1_27/a_38_78# sky130_fd_sc_hs__o21a_1_9/X sky130_fd_sc_hs__dfrbp_1_21/a_910_118#
+ sky130_fd_sc_hs__inv_4_69/Y sky130_fd_sc_hs__nor3_1_5/a_114_368# sky130_fd_sc_hs__o21a_1_35/a_320_74#
+ sky130_fd_sc_hs__dfrtp_4_11/a_699_463# sky130_fd_sc_hs__nor2_1_51/a_116_368# sky130_fd_sc_hs__dfrtn_1_31/a_1550_119#
+ sky130_fd_sc_hs__dfrtp_4_13/a_124_78# sky130_fd_sc_hs__fa_2_19/a_27_378# sky130_fd_sc_hs__a21oi_1_69/a_29_368#
+ sky130_fd_sc_hs__inv_4_133/A sky130_fd_sc_hs__a22oi_1_21/a_71_368# sky130_fd_sc_hs__nand2b_1_3/a_27_112#
+ sky130_fd_sc_hs__o21a_1_7/X sky130_fd_sc_hs__dfrtp_4_19/a_2010_409# sky130_fd_sc_hs__dfrtn_1_19/a_1934_94#
+ sky130_fd_sc_hs__dfrbp_1_15/a_1624_74# sky130_fd_sc_hs__a21oi_1_35/a_29_368# sky130_fd_sc_hs__nor2b_1_27/a_278_368#
+ sky130_fd_sc_hs__nor2_1_1/Y sky130_fd_sc_hs__nor4_1_1/B sky130_fd_sc_hs__a32oi_1_5/a_391_74#
+ sky130_fd_sc_hs__fa_2_15/SUM sky130_fd_sc_hs__nand2_1_71/Y sky130_fd_sc_hs__o21a_1_71/X
+ sky130_fd_sc_hs__dfrtp_4_81/a_1627_493# sky130_fd_sc_hs__dfrbp_1_9/a_1434_74# sky130_fd_sc_hs__dfrtn_1_29/a_33_74#
+ sky130_fd_sc_hs__inv_4_71/A sky130_fd_sc_hs__nor2_1_101/Y sky130_fd_sc_hs__o21a_1_9/B1
+ sky130_fd_sc_hs__sdlclkp_1_1/a_1166_94# sky130_fd_sc_hs__inv_2_3/Y sky130_fd_sc_hs__o31ai_1_7/a_114_74#
+ sky130_fd_sc_hs__a32oi_1_1/a_27_368# sky130_fd_sc_hs__dfrtp_4_71/a_1350_392# sky130_fd_sc_hs__o31ai_1_1/Y
+ sky130_fd_sc_hs__dfrtp_4_7/a_1827_81# sky130_fd_sc_hs__dfrtp_4_7/a_2010_409# sky130_fd_sc_hs__o21a_1_19/X
+ sky130_fd_sc_hs__dfrbp_1_37/a_1224_74# sky130_fd_sc_hs__dfrtn_1_41/a_1547_508# sky130_fd_sc_hs__dfrtp_4_23/a_789_463#
+ sky130_fd_sc_hs__fa_2_19/a_701_79# sky130_fd_sc_hs__dfrtp_4_71/a_1827_81# sky130_fd_sc_hs__o31ai_1_7/Y
+ sky130_fd_sc_hs__a22oi_1_23/Y sky130_fd_sc_hs__dfrtp_4_7/a_313_74# sky130_fd_sc_hs__dfrbp_1_13/a_706_463#
+ sky130_fd_sc_hs__a22o_1_25/a_222_392# sky130_fd_sc_hs__a21oi_1_99/a_117_74# sky130_fd_sc_hs__inv_4_89/A
+ sky130_fd_sc_hs__dfrtn_1_29/a_300_74# sky130_fd_sc_hs__inv_4_7/Y sky130_fd_sc_hs__inv_4_51/Y
+ sky130_fd_sc_hs__nand2_1_91/A sky130_fd_sc_hs__dfrbp_1_43/a_319_360# sky130_fd_sc_hs__dfrtp_4_29/a_494_366#
+ sky130_fd_sc_hs__dfrtp_4_43/a_834_355# sky130_fd_sc_hs__o21a_1_7/A2 sky130_fd_sc_hs__xor2_1_9/a_194_125#
+ sky130_fd_sc_hs__nor3_1_15/a_198_368# sky130_fd_sc_hs__dfrtp_4_67/a_494_366# sky130_fd_sc_hs__dfrtp_4_39/a_1350_392#
+ sky130_fd_sc_hs__dfrtp_4_39/a_313_74# sky130_fd_sc_hs__dfstp_2_1/a_781_74# sky130_fd_sc_hs__dfrtn_1_13/a_120_74#
+ sky130_fd_sc_hs__dfrtn_1_47/a_922_127# sky130_fd_sc_hs__o21a_1_75/A1 sky130_fd_sc_hs__dfrtn_1_45/a_33_74#
+ sky130_fd_sc_hs__inv_4_97/A sky130_fd_sc_hs__dfrtn_1_9/a_856_304# sky130_fd_sc_hs__fa_2_5/B
+ sky130_fd_sc_hs__dfrtp_4_35/a_1678_395# sky130_fd_sc_hs__dfrtn_1_9/a_850_127# sky130_fd_sc_hs__inv_4_99/Y
+ sky130_fd_sc_hs__inv_4_1/A sky130_fd_sc_hs__xnor2_1_11/Y sky130_fd_sc_hs__o21a_1_35/a_376_387#
+ sky130_fd_sc_hs__a21oi_1_115/a_29_368# sky130_fd_sc_hs__inv_4_75/Y sky130_fd_sc_hs__dfrtp_4_83/a_313_74#
+ sky130_fd_sc_hs__inv_4_15/Y sky130_fd_sc_hs__o31ai_1_1/A3 sky130_fd_sc_hs__dfrbp_1_19/D
+ sky130_fd_sc_hs__o21a_1_75/a_376_387# sky130_fd_sc_hs__o21a_1_57/a_83_244# sky130_fd_sc_hs__dfrtp_4_69/a_2010_409#
+ sky130_fd_sc_hs__nand2_2_7/Y sky130_fd_sc_hs__xnor2_1_7/B sky130_fd_sc_hs__dfrbp_1_11/a_910_118#
+ sky130_fd_sc_hs__dfrtn_1_45/a_817_508# sky130_fd_sc_hs__fa_2_15/a_487_79# sky130_fd_sc_hs__inv_4_13/Y
+ sky130_fd_sc_hs__dfrbp_1_3/a_1224_74# sky130_fd_sc_hs__o21a_1_57/X sky130_fd_sc_hs__dfstp_2_7/a_1356_74#
+ sky130_fd_sc_hs__nor2b_1_25/a_27_112# sky130_fd_sc_hs__dfrtp_4_17/a_2010_409# sky130_fd_sc_hs__inv_4_107/Y
+ sky130_fd_sc_hs__nor2b_1_17/a_278_368# sky130_fd_sc_hs__nand2_1_57/a_117_74# sky130_fd_sc_hs__dfrbp_1_41/a_841_401#
+ sky130_fd_sc_hs__nand2_2_13/Y sky130_fd_sc_hs__dfrtp_4_49/a_124_78# sky130_fd_sc_hs__a22o_1_1/a_222_392#
+ sky130_fd_sc_hs__a22oi_1_9/a_339_74# sky130_fd_sc_hs__dfrtn_1_49/a_1934_94# sky130_fd_sc_hs__o21a_1_1/X
+ sky130_fd_sc_hs__fa_2_1/SUM sky130_fd_sc_hs__nand3_1_1/a_233_74# sky130_fd_sc_hs__o21a_1_49/X
+ sky130_fd_sc_hs__dfrtp_4_43/a_812_138# sky130_fd_sc_hs__dfxtp_2_3/a_431_508# sky130_fd_sc_hs__o21a_1_67/A2
+ sky130_fd_sc_hs__o211ai_1_9/C1 sky130_fd_sc_hs__a22oi_1_25/a_71_368# sky130_fd_sc_hs__dfrtp_4_27/a_1647_81#
+ sky130_fd_sc_hs__nand2b_1_7/a_27_112# sky130_fd_sc_hs__dfrtp_4_57/a_37_78# sky130_fd_sc_hs__dfrtp_4_21/a_1827_81#
+ sky130_fd_sc_hs__dfrtp_4_61/a_124_78# sky130_fd_sc_hs__dfxtp_2_1/a_695_459# sky130_fd_sc_hs__xor2_1_1/X
+ sky130_fd_sc_hs__dfrtp_4_13/a_789_463# sky130_fd_sc_hs__dfrbp_1_7/a_2026_424# sky130_fd_sc_hs__dfrtp_4_61/a_1827_81#
+ sky130_fd_sc_hs__a32oi_1_9/a_391_74# sky130_fd_sc_hs__dfrtp_4_89/a_1350_392# sky130_fd_sc_hs__o21a_1_51/a_320_74#
+ sky130_fd_sc_hs__dfrbp_1_45/a_498_360# sky130_fd_sc_hs__a22o_1_15/a_222_392# sky130_fd_sc_hs__dfrtp_4_91/a_789_463#
+ sky130_fd_sc_hs__dfrtp_4_85/a_1678_395# sky130_fd_sc_hs__dfrtp_4_47/a_1627_493#
+ sky130_fd_sc_hs__conb_1_1/HI sky130_fd_sc_hs__dfrtn_1_3/a_33_74# sky130_fd_sc_hs__dfrtn_1_17/a_1736_119#
+ sky130_fd_sc_hs__dfrtp_4_33/a_834_355# sky130_fd_sc_hs__dfrtp_4_19/a_494_366# sky130_fd_sc_hs__o21a_1_31/X
+ sky130_fd_sc_hs__a32oi_1_5/a_27_368# sky130_fd_sc_hs__dfrtn_1_17/a_1266_119# sky130_fd_sc_hs__dfrtp_4_37/a_1350_392#
+ sky130_fd_sc_hs__o21a_1_57/B1 sky130_fd_sc_hs__inv_4_135/A sky130_fd_sc_hs__inv_4_113/A
+ sky130_fd_sc_hs__o22ai_1_5/a_27_74# sky130_fd_sc_hs__dfrtp_4_27/a_890_138# sky130_fd_sc_hs__dfrbp_1_37/a_1465_471#
+ sky130_fd_sc_hs__inv_4_31/Y sky130_fd_sc_hs__o211ai_1_1/a_31_74# sky130_fd_sc_hs__o22ai_1_1/A2
+ sky130_fd_sc_hs__dfxtp_4_3/a_651_503# sky130_fd_sc_hs__o21a_1_65/a_376_387# sky130_fd_sc_hs__o21a_1_77/B1
+ sky130_fd_sc_hs__dfrtp_4_67/a_2010_409# sky130_fd_sc_hs__o21a_1_9/A1 sky130_fd_sc_hs__dfrbp_1_5/Q_N
+ sky130_fd_sc_hs__dfrtn_1_17/a_120_74# sky130_fd_sc_hs__dfrtn_1_35/a_817_508# sky130_fd_sc_hs__nor2b_1_33/Y
+ sky130_fd_sc_hs__dfrtn_1_13/a_33_74# sky130_fd_sc_hs__dfxtp_2_9/a_27_74# sky130_fd_sc_hs__nor2_1_31/a_116_368#
+ sky130_fd_sc_hs__o21a_1_1/a_83_244# sky130_fd_sc_hs__o21a_1_21/X sky130_fd_sc_hs__dfrtn_1_45/a_300_74#
+ sky130_fd_sc_hs__nor2_1_75/B sky130_fd_sc_hs__nand2_1_91/B sky130_fd_sc_hs__o21a_1_61/X
+ sky130_fd_sc_hs__nor2_2_1/a_35_368# sky130_fd_sc_hs__a21oi_1_119/a_29_368# sky130_fd_sc_hs__dfrtp_4_5/a_699_463#
+ sky130_fd_sc_hs__dfrtn_1_7/a_300_74# sky130_fd_sc_hs__dfrtp_4_87/a_313_74# sky130_fd_sc_hs__dfrtn_1_49/a_1550_119#
+ sky130_fd_sc_hs__nor2b_1_41/A sky130_fd_sc_hs__inv_4_5/Y sky130_fd_sc_hs__fa_2_9/a_484_347#
+ sky130_fd_sc_hs__a21oi_1_82/a_117_74# sky130_fd_sc_hs__dfrtn_1_11/a_300_74# sky130_fd_sc_hs__dfrtp_4_53/a_313_74#
+ sky130_fd_sc_hs__fa_2_23/a_336_347# sky130_fd_sc_hs__dfrbp_1_35/a_1624_74# sky130_fd_sc_hs__dfrtn_1_5/a_922_127#
+ sky130_fd_sc_hs__dfrtn_1_39/a_1598_93# sky130_fd_sc_hs__o21a_1_27/a_83_244# sky130_fd_sc_hs__dfrtp_4_33/a_812_138#
+ sky130_fd_sc_hs__fa_2_3/a_27_79# sky130_fd_sc_hs__dfrbp_1_21/a_125_78# sky130_fd_sc_hs__fa_2_19/a_484_347#
+ sky130_fd_sc_hs__dfrtn_1_5/a_1547_508# sky130_fd_sc_hs__nor2b_1_29/a_27_112# sky130_fd_sc_hs__nor2b_1_1/a_27_112#
+ sky130_fd_sc_hs__a22o_1_25/a_230_79# sky130_fd_sc_hs__nor4_1_3/C sky130_fd_sc_hs__nor2_2_3/Y
+ sky130_fd_sc_hs__dfrbp_1_5/a_1482_48# sky130_fd_sc_hs__dfrtp_4_5/a_2010_409# sky130_fd_sc_hs__o2bb2ai_1_1/a_114_74#
+ sky130_fd_sc_hs__fa_2_7/CIN sky130_fd_sc_hs__o21ai_1_1/Y sky130_fd_sc_hs__dfrbp_1_37/a_38_78#
+ sky130_fd_sc_hs__dfrtp_4_51/a_1827_81# sky130_fd_sc_hs__nand2_4_5/Y sky130_fd_sc_hs__inv_4_37/Y
+ sky130_fd_sc_hs__inv_4_17/A sky130_fd_sc_hs__o21ai_1_5/B1 sky130_fd_sc_hs__dfrtn_1_1/a_817_508#
+ sky130_fd_sc_hs__inv_4_35/A sky130_fd_sc_hs__dfrtp_4_1/a_124_78# sky130_fd_sc_hs__dfrtn_1_31/D
+ sky130_fd_sc_hs__dfrtp_4_81/a_789_463# sky130_fd_sc_hs__fa_2_13/SUM sky130_fd_sc_hs__a222oi_1_1/Y
+ sky130_fd_sc_hs__dfrbp_1_33/a_706_463# sky130_fd_sc_hs__dfrbp_1_23/a_319_360# sky130_fd_sc_hs__dfrtp_4_23/a_834_355#
+ sky130_fd_sc_hs__fa_2_15/a_1119_79# sky130_fd_sc_hs__dfrtp_4_25/a_37_78# sky130_fd_sc_hs__dfrtp_4_65/a_124_78#
+ sky130_fd_sc_hs__dfrtp_4_47/a_494_366# sky130_fd_sc_hs__dfxtp_4_5/a_27_74# sky130_fd_sc_hs__dfxtp_4_9/a_1178_124#
+ sky130_fd_sc_hs__dfrtn_1_27/a_922_127# sky130_fd_sc_hs__dfrtp_4_87/a_494_366# sky130_fd_sc_hs__o211ai_1_7/a_116_368#
+ sky130_fd_sc_hs__o21a_1_55/a_320_74# sky130_fd_sc_hs__a222o_1_1/X sky130_fd_sc_hs__a32oi_1_1/a_119_74#
+ sky130_fd_sc_hs__dfrbp_1_41/a_1434_74# sky130_fd_sc_hs__dfrtp_4_33/a_1678_395# sky130_fd_sc_hs__o21a_1_21/A1
+ sky130_fd_sc_hs__dfrbp_1_29/a_1482_48# sky130_fd_sc_hs__inv_4_127/A sky130_fd_sc_hs__xnor2_1_1/a_112_119#
+ sky130_fd_sc_hs__nor2b_1_21/Y sky130_fd_sc_hs__a22oi_1_5/a_71_368# sky130_fd_sc_hs__o21a_1_55/a_376_387#
+ sky130_fd_sc_hs__a21oi_1_55/a_29_368# sky130_fd_sc_hs__a32oi_1_9/a_27_368# sky130_fd_sc_hs__nor2_1_61/Y
+ sky130_fd_sc_hs__dfrtn_1_7/a_507_368# sky130_fd_sc_hs__fa_2_3/a_992_347# sky130_fd_sc_hs__dfrtn_1_25/a_817_508#
+ sky130_fd_sc_hs__dfstp_2_4/a_1566_92# sky130_fd_sc_hs__nor2_1_95/A sky130_fd_sc_hs__nor2_1_65/A
+ sky130_fd_sc_hs__nor2_1_21/a_116_368# sky130_fd_sc_hs__o21a_1_1/a_376_387# sky130_fd_sc_hs__nor2_1_3/Y
+ sky130_fd_sc_hs__dfrtp_4_41/a_37_78# sky130_fd_sc_hs__nor2_1_21/B sky130_fd_sc_hs__dfrbp_1_1/a_498_360#
+ sky130_fd_sc_hs__nand2_2_9/a_27_74# sky130_fd_sc_hs__dfrtn_1_47/a_1550_119# sky130_fd_sc_hs__sdlclkp_4_1/a_116_395#
+ sky130_fd_sc_hs__a22oi_1_1/Y sky130_fd_sc_hs__dfrtp_4_15/a_2010_409# sky130_fd_sc_hs__dfrbp_1_9/a_706_463#
+ sky130_fd_sc_hs__a22o_1_21/a_132_392# sky130_fd_sc_hs__fa_2_13/a_336_347# sky130_fd_sc_hs__dfrtn_1_29/a_1598_93#
+ sky130_fd_sc_hs__nor2b_1_35/a_278_368# sky130_fd_sc_hs__inv_2_7/A sky130_fd_sc_hs__xnor2_1_1/a_293_74#
+ sky130_fd_sc_hs__dfrtp_4_23/a_812_138# sky130_fd_sc_hs__o21a_1_5/a_83_244# sky130_fd_sc_hs__dfstp_2_5/a_716_456#
+ sky130_fd_sc_hs__dfrtn_1_49/a_300_74# sky130_fd_sc_hs__o21a_1_53/X sky130_fd_sc_hs__nor2_1_49/B
+ sky130_fd_sc_hs__and2_2_1/a_31_74# sky130_fd_sc_hs__inv_4_1/Y sky130_fd_sc_hs__nand2_1_67/Y
+ sky130_fd_sc_hs__a21oi_1_85/a_117_74# sky130_fd_sc_hs__fa_2_15/CIN sky130_fd_sc_hs__inv_2_9/A
+ sky130_fd_sc_hs__fa_2_5/a_683_347# sky130_fd_sc_hs__fa_2_23/CIN sky130_fd_sc_hs__dfrtn_1_33/a_120_74#
+ sky130_fd_sc_hs__inv_4_51/A sky130_fd_sc_hs__a21oi_1_51/a_117_74# sky130_fd_sc_hs__dfrtp_4_41/a_1827_81#
+ sky130_fd_sc_hs__dfrtn_1_47/a_714_127# sky130_fd_sc_hs__dfrtp_4_87/a_1350_392# sky130_fd_sc_hs__dfrtp_4_85/a_1647_81#
+ sky130_fd_sc_hs__dfrbp_1_45/a_1224_74# sky130_fd_sc_hs__dfrtp_4_7/a_789_463# sky130_fd_sc_hs__dfrbp_1_25/a_498_360#
+ sky130_fd_sc_hs__fa_2_13/CIN sky130_fd_sc_hs__dfrtp_4_71/a_789_463# sky130_fd_sc_hs__dfrtp_4_83/a_1678_395#
+ sky130_fd_sc_hs__a222oi_1_1/a_116_392# sky130_fd_sc_hs__dfrbp_1_31/Q_N sky130_fd_sc_hs__dfxtp_2_9/a_644_504#
+ sky130_fd_sc_hs__a22o_1_27/X sky130_fd_sc_hs__dfrbp_1_13/a_319_360# sky130_fd_sc_hs__dfrtp_4_13/a_834_355#
+ sky130_fd_sc_hs__a21oi_1_101/a_29_368# sky130_fd_sc_hs__a22o_1_29/a_230_79# sky130_fd_sc_hs__dfrtp_4_37/a_494_366#
+ sky130_fd_sc_hs__nand2_1_111/a_117_74# sky130_fd_sc_hs__a21oi_1_1/a_117_74# sky130_fd_sc_hs__sdlclkp_4_1/a_792_48#
+ sky130_fd_sc_hs__dfrtp_4_3/a_494_366# sky130_fd_sc_hs__inv_4_53/A sky130_fd_sc_hs__o21ai_1_5/a_162_368#
+ sky130_fd_sc_hs__dfrtn_1_17/a_922_127# sky130_fd_sc_hs__o21a_1_43/a_83_244# sky130_fd_sc_hs__dfrtp_4_77/a_494_366#
+ sky130_fd_sc_hs__dfrtp_4_91/a_834_355# sky130_fd_sc_hs__dfxtp_2_11/a_206_368# sky130_fd_sc_hs__nor2_1_91/Y
+ sky130_fd_sc_hs__dfrtn_1_33/D sky130_fd_sc_hs__a21oi_1_19/Y sky130_fd_sc_hs__nand2_4_5/a_27_74#
+ sky130_fd_sc_hs__a22o_1_9/a_132_392# sky130_fd_sc_hs__dfxtp_2_11/a_1125_508# sky130_fd_sc_hs__dfrbp_1_19/a_1482_48#
+ sky130_fd_sc_hs__dfrbp_1_35/a_1465_471# sky130_fd_sc_hs__o21a_1_45/a_376_387# sky130_fd_sc_hs__dfrtp_4_69/a_124_78#
+ sky130_fd_sc_hs__nor2b_1_11/a_27_112# sky130_fd_sc_hs__nor2b_1_29/Y sky130_fd_sc_hs__nor2_1_51/B
+ sky130_fd_sc_hs__nand2_4_7/A sky130_fd_sc_hs__dfrtp_4_85/a_890_138# sky130_fd_sc_hs__o21a_1_59/a_320_74#
+ sky130_fd_sc_hs__dfrtn_1_15/a_817_508# sky130_fd_sc_hs__a32oi_1_5/a_119_74# sky130_fd_sc_hs__dfxtp_4_9/a_735_102#
+ sky130_fd_sc_hs__nor2_1_11/a_116_368# sky130_fd_sc_hs__o21a_1_71/A2 sky130_fd_sc_hs__o211ai_1_5/a_311_74#
+ sky130_fd_sc_hs__conb_1_1/LO sky130_fd_sc_hs__fa_2_21/SUM sky130_fd_sc_hs__nor2b_1_13/Y
+ sky130_fd_sc_hs__dfrbp_1_19/a_2026_424# sky130_fd_sc_hs__a21oi_1_59/a_29_368# sky130_fd_sc_hs__nor2_1_23/Y
+ sky130_fd_sc_hs__dfrbp_1_21/a_38_78# sky130_fd_sc_hs__a22oi_1_11/a_71_368# sky130_fd_sc_hs__dfrtn_1_19/a_1598_93#
+ sky130_fd_sc_hs__inv_4_67/A sky130_fd_sc_hs__dfrtp_4_13/a_812_138# sky130_fd_sc_hs__inv_4_3/Y
+ sky130_fd_sc_hs__dfrbp_1_29/D sky130_fd_sc_hs__dfrtp_4_81/a_37_78# sky130_fd_sc_hs__fa_2_21/a_27_378#
+ sky130_fd_sc_hs__dfrtn_1_3/a_1547_508# sky130_fd_sc_hs__xnor2_1_9/B sky130_fd_sc_hs__dfrtp_4_91/a_812_138#
+ sky130_fd_sc_hs__fa_2_9/a_1205_79# sky130_fd_sc_hs__dfrtp_4_1/a_1647_81# sky130_fd_sc_hs__dfrbp_1_5/a_2026_424#
+ sky130_fd_sc_hs__dfrtp_4_31/a_1827_81# sky130_fd_sc_hs__xnor2_1_5/a_293_74# sky130_fd_sc_hs__dfrtp_4_75/a_1647_81#
+ sky130_fd_sc_hs__dfrtp_4_21/a_789_463# sky130_fd_sc_hs__dfrtn_1_23/a_33_74# sky130_fd_sc_hs__dfrbp_1_15/a_498_360#
+ sky130_fd_sc_hs__dfrbp_1_39/a_796_463# sky130_fd_sc_hs__fa_2_1/A sky130_fd_sc_hs__a22o_1_25/a_52_123#
+ sky130_fd_sc_hs__dfrtp_4_61/a_789_463# sky130_fd_sc_hs__dfrtp_4_45/a_1627_493# sky130_fd_sc_hs__dfrtn_1_15/a_1736_119#
+ sky130_fd_sc_hs__maj3_1_1/X sky130_fd_sc_hs__a21oi_1_89/a_117_74# sky130_fd_sc_hs__xor2_1_11/a_355_368#
+ sky130_fd_sc_hs__a222oi_1_3/a_461_74# sky130_fd_sc_hs__dfrtn_1_19/a_300_74# sky130_fd_sc_hs__dfrtn_1_15/a_1266_119#
+ sky130_fd_sc_hs__fa_2_19/a_1205_79# sky130_fd_sc_hs__dfrbp_1_1/Q sky130_fd_sc_hs__dfrtp_4_35/a_1350_392#
+ sky130_fd_sc_hs__dfrtn_1_37/a_120_74# sky130_fd_sc_hs__inv_4_81/A sky130_fd_sc_hs__xor2_1_7/a_194_125#
+ sky130_fd_sc_hs__dfxtp_4_7/a_1178_124# sky130_fd_sc_hs__nor2_1_15/Y sky130_fd_sc_hs__dfrtp_4_81/a_834_355#
+ sky130_fd_sc_hs__o21a_1_23/X sky130_fd_sc_hs__fa_2_21/a_701_79# sky130_fd_sc_hs__inv_4_97/Y
+ sky130_fd_sc_hs__dfrtp_4_29/a_313_74# sky130_fd_sc_hs__xnor2_1_7/A sky130_fd_sc_hs__dfrtp_4_31/a_1678_395#
+ sky130_fd_sc_hs__a21oi_1_23/a_117_74# sky130_fd_sc_hs__dfrtn_1_7/a_856_304# sky130_fd_sc_hs__dfrbp_1_29/a_125_78#
+ sky130_fd_sc_hs__dfrtn_1_7/a_850_127# sky130_fd_sc_hs__dfrtp_4_49/a_1678_395# sky130_fd_sc_hs__dfrbp_1_47/a_1482_48#
+ sky130_fd_sc_hs__dfrbp_1_3/a_125_78# sky130_fd_sc_hs__o21ai_1_9/a_27_74# sky130_fd_sc_hs__dfrbp_1_31/a_832_118#
+ sky130_fd_sc_hs__dfrtp_4_65/a_2010_409# sky130_fd_sc_hs__a21oi_1_5/a_117_74# sky130_fd_sc_hs__dfrtp_4_1/a_890_138#
+ sky130_fd_sc_hs__dfrbp_1_45/a_38_78# sky130_fd_sc_hs__sdlclkp_4_1/a_324_79# sky130_fd_sc_hs__dfrtn_1_5/a_714_127#
+ sky130_fd_sc_hs__dfrtp_4_75/a_890_138# sky130_fd_sc_hs__fa_2_17/CIN sky130_fd_sc_hs__o21a_1_47/a_83_244#
+ sky130_fd_sc_hs__a22o_1_1/a_230_79# sky130_fd_sc_hs__o21a_1_13/a_83_244# sky130_fd_sc_hs__dfrbp_1_1/a_1224_74#
+ sky130_fd_sc_hs__o21a_1_3/a_320_74# sky130_fd_sc_hs__nor2_1_43/B sky130_fd_sc_hs__dfrbp_1_17/a_2026_424#
+ sky130_fd_sc_hs__dfrtp_4_49/a_699_463# sky130_fd_sc_hs__or3b_2_1/C_N sky130_fd_sc_hs__dfrtp_4_35/a_37_78#
+ sky130_fd_sc_hs__and2_2_1/a_118_74# sky130_fd_sc_hs__dfrtp_4_89/a_699_463# sky130_fd_sc_hs__nor2b_1_15/a_27_112#
+ sky130_fd_sc_hs__inv_4_35/Y sky130_fd_sc_hs__o21a_1_47/X sky130_fd_sc_hs__a22o_1_11/a_230_79#
+ sky130_fd_sc_hs__nor3_1_9/a_198_368# sky130_fd_sc_hs__nand2_1_47/a_117_74# sky130_fd_sc_hs__inv_4_47/Y
+ sky130_fd_sc_hs__inv_4_9/A sky130_fd_sc_hs__nand2_4_11/a_27_74# sky130_fd_sc_hs__a32oi_1_9/a_119_74#
+ sky130_fd_sc_hs__dfrtn_1_47/a_1934_94# sky130_fd_sc_hs__dfrbp_1_43/a_1624_74# sky130_fd_sc_hs__dfrtn_1_49/a_1598_93#
+ sky130_fd_sc_hs__dfrtn_1_47/a_33_74# sky130_fd_sc_hs__sdlclkp_4_1/a_354_105# sky130_fd_sc_hs__dfrtn_1_1/a_1547_508#
+ sky130_fd_sc_hs__nand2_1_91/a_117_74# sky130_fd_sc_hs__dfrtp_4_81/a_812_138# sky130_fd_sc_hs__a32oi_1_7/Y
+ sky130_fd_sc_hs__a21oi_1_9/Y sky130_fd_sc_hs__nand2_1_99/A sky130_fd_sc_hs__dfrtp_4_3/a_2010_409#
+ sky130_fd_sc_hs__a22oi_1_15/a_71_368# sky130_fd_sc_hs__xnor2_1_1/a_138_385# sky130_fd_sc_hs__dfrtp_4_25/a_1647_81#
+ sky130_fd_sc_hs__dfrtn_1_27/a_714_127# sky130_fd_sc_hs__dfrtp_4_85/a_1350_392# sky130_fd_sc_hs__dfrbp_1_7/a_832_118#
+ sky130_fd_sc_hs__dfrtp_4_51/a_124_78# sky130_fd_sc_hs__dfrtp_4_65/a_1647_81# sky130_fd_sc_hs__dfrbp_1_25/a_1224_74#
+ sky130_fd_sc_hs__dfrbp_1_7/Q_N sky130_fd_sc_hs__nor2_1_3/B sky130_fd_sc_hs__maj3_1_1/a_84_74#
+ sky130_fd_sc_hs__o21a_1_41/a_320_74# sky130_fd_sc_hs__inv_4_31/A sky130_fd_sc_hs__dfrtp_4_81/a_1678_395#
+ sky130_fd_sc_hs__dfrtp_4_85/D sky130_fd_sc_hs__dfrtp_4_51/a_789_463# sky130_fd_sc_hs__dfrtn_1_13/a_1736_119#
+ sky130_fd_sc_hs__xor2_1_7/a_455_87# sky130_fd_sc_hs__a22o_1_13/a_222_392# sky130_fd_sc_hs__dfrtn_1_13/a_1266_119#
+ sky130_fd_sc_hs__dfrbp_1_41/a_706_463# sky130_fd_sc_hs__dfrtp_4_7/a_834_355# sky130_fd_sc_hs__o21a_1_19/A1
+ sky130_fd_sc_hs__o21a_1_5/A1 sky130_fd_sc_hs__dfrbp_1_33/a_319_360# sky130_fd_sc_hs__dfrtp_4_17/a_494_366#
+ sky130_fd_sc_hs__a21oi_1_41/a_29_368# sky130_fd_sc_hs__inv_4_111/A sky130_fd_sc_hs__inv_4_9/Y
+ sky130_fd_sc_hs__dfrtp_4_57/a_494_366# sky130_fd_sc_hs__dfrtp_4_71/a_834_355# sky130_fd_sc_hs__xnor2_1_9/a_293_74#
+ sky130_fd_sc_hs__dfrtn_1_37/a_922_127# sky130_fd_sc_hs__nand2_2_1/A sky130_fd_sc_hs__a22o_1_29/a_52_123#
+ sky130_fd_sc_hs__dfrbp_1_33/a_1465_471# sky130_fd_sc_hs__o21a_1_25/a_376_387# sky130_fd_sc_hs__dfrtp_4_25/a_890_138#
+ sky130_fd_sc_hs__dfrbp_1_21/a_832_118# sky130_fd_sc_hs__dfrtp_4_63/a_2010_409# sky130_fd_sc_hs__dfxtp_4_2/a_651_503#
+ sky130_fd_sc_hs__nor2_1_7/A sky130_fd_sc_hs__inv_4_121/Y sky130_fd_sc_hs__o31ai_1_3/B1
+ sky130_fd_sc_hs__dfrtp_4_65/a_890_138# sky130_fd_sc_hs__nor2b_1_11/Y sky130_fd_sc_hs__nor2_1_73/B
+ sky130_fd_sc_hs__dfrbp_1_31/D sky130_fd_sc_hs__o21a_1_77/X sky130_fd_sc_hs__a21oi_1_27/a_117_74#
+ sky130_fd_sc_hs__fa_2_19/a_1094_347# sky130_fd_sc_hs__nor2_1_89/A sky130_fd_sc_hs__inv_4_61/Y
+ sky130_fd_sc_hs__nor2_1_75/Y sky130_fd_sc_hs__dfrtn_1_45/a_1550_119# sky130_fd_sc_hs__nand4_2_1/D
+ sky130_fd_sc_hs__dfrtn_1_35/a_300_74# sky130_fd_sc_hs__dfxtp_2_9/a_538_429# sky130_fd_sc_hs__dfrtp_4_13/a_2010_409#
+ sky130_fd_sc_hs__dfrtp_4_77/a_313_74# sky130_fd_sc_hs__dfrtp_4_79/a_699_463# sky130_fd_sc_hs__a21oi_1_71/a_117_74#
+ sky130_fd_sc_hs__a21oi_1_9/a_117_74# sky130_fd_sc_hs__dfxtp_2_11/a_708_101# sky130_fd_sc_hs__nor2_1_115/a_116_368#
+ sky130_fd_sc_hs__dfxtp_2_1/a_27_74# sky130_fd_sc_hs__dfrbp_1_9/a_319_360# sky130_fd_sc_hs__dfrbp_1_31/a_841_401#
+ sky130_fd_sc_hs__nor2_1_77/Y sky130_fd_sc_hs__fa_2_23/a_992_347# sky130_fd_sc_hs__a22o_1_5/a_230_79#
+ sky130_fd_sc_hs__nor2b_1_45/a_278_368# sky130_fd_sc_hs__inv_4_137/Y sky130_fd_sc_hs__dfrtp_4_11/a_313_74#
+ sky130_fd_sc_hs__dfrtp_4_7/a_812_138# sky130_fd_sc_hs__dfrbp_1_43/a_125_78# sky130_fd_sc_hs__nor4_1_3/A
+ sky130_fd_sc_hs__o21a_1_7/a_320_74# sky130_fd_sc_hs__dfrtp_4_71/a_812_138# sky130_fd_sc_hs__dfrtp_4_75/a_37_78#
+ sky130_fd_sc_hs__o21a_1_75/X sky130_fd_sc_hs__dfrbp_1_11/a_125_78# sky130_fd_sc_hs__and2_2_5/a_118_74#
+ sky130_fd_sc_hs__nor2b_1_19/a_27_112# sky130_fd_sc_hs__dfrtp_4_15/a_1647_81# sky130_fd_sc_hs__o21a_1_29/X
+ sky130_fd_sc_hs__a22o_1_15/a_230_79# sky130_fd_sc_hs__fa_2_3/a_1119_79# sky130_fd_sc_hs__dfrbp_1_3/a_2026_424#
+ sky130_fd_sc_hs__dfrtp_4_11/a_1827_81# sky130_fd_sc_hs__dfrtn_1_17/a_714_127# sky130_fd_sc_hs__o22ai_1_1/A1
+ sky130_fd_sc_hs__and2_2_1/X sky130_fd_sc_hs__dfrtp_4_55/a_1647_81# sky130_fd_sc_hs__dfrbp_1_15/a_1224_74#
+ sky130_fd_sc_hs__fa_2_17/B sky130_fd_sc_hs__dfrtn_1_39/a_507_368# sky130_fd_sc_hs__dfxtp_2_5/D
+ sky130_fd_sc_hs__nand2b_4_1/a_243_74# sky130_fd_sc_hs__dfrtp_4_41/a_789_463# sky130_fd_sc_hs__dfrtp_4_43/a_1627_493#
+ sky130_fd_sc_hs__dfrbp_1_35/a_498_360# sky130_fd_sc_hs__a22oi_1_21/a_159_74# sky130_fd_sc_hs__nand2_1_95/a_117_74#
+ sky130_fd_sc_hs__a32oi_1_5/Y sky130_fd_sc_hs__fa_2_5/A sky130_fd_sc_hs__a22oi_1_19/a_71_368#
+ sky130_fd_sc_hs__dfrtp_4_21/a_834_355# sky130_fd_sc_hs__dfrtp_4_33/a_1350_392# sky130_fd_sc_hs__inv_4_71/Y
+ sky130_fd_sc_hs__dfxtp_4_5/a_1178_124# sky130_fd_sc_hs__a21oi_1_105/a_117_74# sky130_fd_sc_hs__dfrtp_4_55/a_124_78#
+ sky130_fd_sc_hs__dfrtp_4_61/a_834_355# sky130_fd_sc_hs__sdlclkp_1_1/a_722_492# sky130_fd_sc_hs__a222oi_1_3/a_369_392#
+ sky130_fd_sc_hs__dfrtn_1_5/a_1934_94# sky130_fd_sc_hs__o211ai_1_5/a_116_368# sky130_fd_sc_hs__o21a_1_45/a_320_74#
+ sky130_fd_sc_hs__dfrbp_1_7/a_841_401# sky130_fd_sc_hs__dfrtp_4_21/a_124_78# sky130_fd_sc_hs__inv_4_101/A
+ sky130_fd_sc_hs__a21oi_1_77/a_29_368# sky130_fd_sc_hs__dfrtp_4_47/a_1678_395# sky130_fd_sc_hs__o21a_1_11/a_320_74#
+ sky130_fd_sc_hs__o21a_1_15/a_376_387# sky130_fd_sc_hs__dfrbp_1_27/a_1482_48# sky130_fd_sc_hs__dfrtp_4_15/a_890_138#
+ sky130_fd_sc_hs__dfrbp_1_11/a_832_118# sky130_fd_sc_hs__a21oi_1_45/a_29_368# sky130_fd_sc_hs__inv_4_85/A
+ sky130_fd_sc_hs__dfrtp_4_55/a_890_138# sky130_fd_sc_hs__a21oi_1_11/a_29_368# sky130_fd_sc_hs__dfrbp_1_39/a_38_78#
+ sky130_fd_sc_hs__dfrtn_1_9/a_1550_119# sky130_fd_sc_hs__dfrtn_1_31/a_33_74# sky130_fd_sc_hs__fa_2_1/a_336_347#
+ sky130_fd_sc_hs__dfxtp_4_3/a_696_458# sky130_fd_sc_hs__dfstp_2_1/a_1566_92# sky130_fd_sc_hs__dfrbp_1_39/a_910_118#
+ sky130_fd_sc_hs__dfrtp_4_35/D sky130_fd_sc_hs__dfrbp_1_15/a_2026_424# sky130_fd_sc_hs__nor2b_1_1/a_278_368#
+ sky130_fd_sc_hs__dfrtp_4_69/a_699_463# sky130_fd_sc_hs__a22o_1_1/a_52_123# sky130_fd_sc_hs__dfrtp_4_29/a_37_78#
+ sky130_fd_sc_hs__nor2_1_105/a_116_368# sky130_fd_sc_hs__dfxtp_4_2/D sky130_fd_sc_hs__fa_2_1/a_487_79#
+ sky130_fd_sc_hs__dfrbp_1_21/a_841_401# sky130_fd_sc_hs__o21a_1_51/X sky130_fd_sc_hs__dfrbp_1_23/a_1624_74#
+ sky130_fd_sc_hs__fa_2_11/a_336_347# sky130_fd_sc_hs__dfrtn_1_27/a_1934_94# sky130_fd_sc_hs__fa_2_13/a_992_347#
+ sky130_fd_sc_hs__dfrbp_1_15/Q_N sky130_fd_sc_hs__dfrbp_1_11/D sky130_fd_sc_hs__dfrtp_4_21/a_812_138#
+ sky130_fd_sc_hs__a22o_1_11/a_52_123# sky130_fd_sc_hs__dfstp_2_4/a_716_456# sky130_fd_sc_hs__dfrtp_4_61/a_812_138#
+ sky130_fd_sc_hs__dfrtp_4_1/a_2010_409# sky130_fd_sc_hs__a21oi_1_75/a_117_74# sky130_fd_sc_hs__o22ai_1_9/a_340_368#
+ sky130_fd_sc_hs__dfrbp_1_1/a_2026_424# sky130_fd_sc_hs__dfstp_2_4/a_27_74# sky130_fd_sc_hs__dfrtp_4_83/a_1350_392#
+ sky130_fd_sc_hs__dfrtp_4_47/a_313_74# sky130_fd_sc_hs__nand2_1_85/Y sky130_fd_sc_hs__dfrtp_4_45/a_1647_81#
+ sky130_fd_sc_hs__a222o_1_1/a_27_390# sky130_fd_sc_hs__dfrtn_1_23/a_120_74# sky130_fd_sc_hs__dfrtn_1_29/a_507_368#
+ sky130_fd_sc_hs__nor2b_1_3/Y sky130_fd_sc_hs__a22o_1_9/a_230_79# sky130_fd_sc_hs__dfrtp_4_31/a_789_463#
+ sky130_fd_sc_hs__dfrbp_1_47/a_125_78# sky130_fd_sc_hs__xor2_1_3/a_355_368# sky130_fd_sc_hs__inv_4_109/Y
+ sky130_fd_sc_hs__dfrtn_1_11/a_1736_119# sky130_fd_sc_hs__a21oi_1_123/a_29_368# sky130_fd_sc_hs__dfrtn_1_11/a_1266_119#
+ sky130_fd_sc_hs__dfxtp_2_7/a_644_504# sky130_fd_sc_hs__or2_1_3/a_63_368# sky130_fd_sc_hs__a22o_1_19/a_230_79#
+ sky130_fd_sc_hs__fa_2_15/a_683_347# sky130_fd_sc_hs__a31oi_1_1/a_145_74# sky130_fd_sc_hs__dfrtp_4_51/a_834_355#
+ sky130_fd_sc_hs__maj3_1_3/X sky130_fd_sc_hs__o21a_1_33/a_83_244# sky130_fd_sc_hs__dfstp_2_7/D
+ sky130_fd_sc_hs__dfrbp_1_31/a_1434_74# sky130_fd_sc_hs__o21a_1_3/X sky130_fd_sc_hs__dfrbp_1_31/a_1465_471#
+ sky130_fd_sc_hs__a22oi_1_25/a_159_74# sky130_fd_sc_hs__nand2b_1_3/Y sky130_fd_sc_hs__dfrbp_1_17/a_1482_48#
+ sky130_fd_sc_hs__nand3b_2_1/a_403_54# sky130_fd_sc_hs__o22ai_1_3/Y sky130_fd_sc_hs__a21oi_1_109/a_117_74#
+ sky130_fd_sc_hs__dfrtp_4_45/a_890_138# sky130_fd_sc_hs__dfrtp_4_59/a_124_78# sky130_fd_sc_hs__dfrtn_1_7/a_1550_119#
+ sky130_fd_sc_hs__nand2_1_33/a_117_74# sky130_fd_sc_hs__o21a_1_49/a_320_74# sky130_fd_sc_hs__dfrtn_1_13/a_817_508#
+ sky130_fd_sc_hs__fa_2_17/a_1094_347# sky130_fd_sc_hs__dfrtp_4_25/a_124_78# sky130_fd_sc_hs__dfrtn_1_43/a_1550_119#
+ sky130_fd_sc_hs__nor3_1_3/a_114_368# sky130_fd_sc_hs__xnor2_1_11/a_293_74# sky130_fd_sc_hs__o22ai_1_9/A1
+ sky130_fd_sc_hs__dfrtp_4_11/a_2010_409# sky130_fd_sc_hs__dfrtp_4_59/a_699_463# sky130_fd_sc_hs__nor2_1_99/a_116_368#
+ sky130_fd_sc_hs__nor2_1_59/A sky130_fd_sc_hs__a21oi_1_121/a_117_74# sky130_fd_sc_hs__dfrbp_1_11/a_841_401#
+ sky130_fd_sc_hs__a22o_1_11/a_132_392# sky130_fd_sc_hs__dfrtn_1_17/a_1934_94# sky130_fd_sc_hs__dfrbp_1_13/a_1624_74#
+ sky130_fd_sc_hs__clkbuf_2_1/a_43_192# sky130_fd_sc_hs__nor2b_1_25/a_278_368# sky130_fd_sc_hs__o21a_1_15/X
+ sky130_fd_sc_hs__a21oi_1_93/a_29_368# sky130_fd_sc_hs__nand2_4_7/a_27_74# sky130_fd_sc_hs__dfrtp_4_51/a_812_138#
+ sky130_fd_sc_hs__dfrtn_1_39/a_856_304# sky130_fd_sc_hs__nor3_1_1/C sky130_fd_sc_hs__nor2_1_9/B
+ sky130_fd_sc_hs__maj3_1_3/a_226_384# sky130_fd_sc_hs__dfrbp_1_7/a_1434_74# sky130_fd_sc_hs__dfrtn_1_39/a_850_127#
+ sky130_fd_sc_hs__a22o_1_5/a_52_123# sky130_fd_sc_hs__dfrtp_4_69/a_37_78# sky130_fd_sc_hs__fa_2_5/a_487_79#
+ sky130_fd_sc_hs__dfrtp_4_35/a_1647_81# sky130_fd_sc_hs__nor2_1_83/Y sky130_fd_sc_hs__dfrtn_1_19/a_507_368#
+ sky130_fd_sc_hs__dfrtp_4_5/a_1827_81# sky130_fd_sc_hs__nand4_1_1/Y sky130_fd_sc_hs__dfrtn_1_37/a_714_127#
+ sky130_fd_sc_hs__dfrtp_4_73/a_1647_81# sky130_fd_sc_hs__dfrbp_1_35/a_1224_74# sky130_fd_sc_hs__dfrtp_4_41/a_1627_493#
+ sky130_fd_sc_hs__a22o_1_15/a_52_123# sky130_fd_sc_hs__o22ai_1_9/a_142_368# sky130_fd_sc_hs__dfstp_2_5/a_1278_74#
+ sky130_fd_sc_hs__a22o_1_23/a_222_392# sky130_fd_sc_hs__dfrtn_1_29/a_1736_119# sky130_fd_sc_hs__inv_4_95/Y
+ sky130_fd_sc_hs__dfrtp_4_31/a_1350_392# sky130_fd_sc_hs__dfrbp_1_23/a_38_78# sky130_fd_sc_hs__dfrbp_1_41/a_319_360#
+ sky130_fd_sc_hs__dfrtp_4_27/a_494_366# sky130_fd_sc_hs__dfrtp_4_41/a_834_355# sky130_fd_sc_hs__dfrtn_1_29/a_1266_119#
+ sky130_fd_sc_hs__dfrtp_4_49/a_1350_392# sky130_fd_sc_hs__a21oi_1_82/Y sky130_fd_sc_hs__nor3_1_13/a_198_368#
+ sky130_fd_sc_hs__dfrtp_4_19/a_313_74# sky130_fd_sc_hs__dfrbp_1_21/a_1434_74# sky130_fd_sc_hs__a21oi_1_13/a_117_74#
+ sky130_fd_sc_hs__o2bb2ai_1_1/a_131_383# sky130_fd_sc_hs__dfrbp_1_19/a_125_78# sky130_fd_sc_hs__dfrtp_4_13/a_37_78#
+ sky130_fd_sc_hs__dfrtp_4_61/a_2010_409# sky130_fd_sc_hs__nand4_1_1/a_259_74# sky130_fd_sc_hs__dfxtp_2_5/a_206_368#
+ sky130_fd_sc_hs__dfrtp_4_35/a_890_138# sky130_fd_sc_hs__a31oi_1_1/A2 sky130_fd_sc_hs__o21a_1_73/a_376_387#
+ sky130_fd_sc_hs__nor4_1_3/D sky130_fd_sc_hs__dfrtp_4_73/a_890_138# sky130_fd_sc_hs__nor3_1_9/A
+ sky130_fd_sc_hs__nor2b_1_1/Y sky130_fd_sc_hs__dfsbp_2_1/Q sky130_fd_sc_hs__dfrtn_1_43/a_817_508#
+ sky130_fd_sc_hs__dfrtn_1_41/a_1550_119# sky130_fd_sc_hs__dfrbp_1_13/a_2026_424#
+ sky130_fd_sc_hs__nor2_1_41/B sky130_fd_sc_hs__o21a_1_45/X sky130_fd_sc_hs__dfrbp_1_5/a_796_463#
+ sky130_fd_sc_hs__nor2_1_89/a_116_368# sky130_fd_sc_hs__dfrtp_4_29/a_2010_409# sky130_fd_sc_hs__nor2b_1_15/a_278_368#
+ sky130_fd_sc_hs__nand2_1_37/a_117_74# sky130_fd_sc_hs__a22oi_1_23/a_339_74# sky130_fd_sc_hs__dfsbp_2_1/a_1501_92#
+ sky130_fd_sc_hs__dfrtn_1_47/a_1598_93# sky130_fd_sc_hs__dfsbp_2_1/a_1521_508# sky130_fd_sc_hs__dfrtp_4_91/a_1627_493#
+ sky130_fd_sc_hs__a22oi_1_5/a_159_74# sky130_fd_sc_hs__xnor2_1_15/a_293_74# sky130_fd_sc_hs__dfrtp_4_41/a_812_138#
+ sky130_fd_sc_hs__dfrtn_1_29/a_856_304# sky130_fd_sc_hs__dfrtn_1_29/a_850_127# sky130_fd_sc_hs__dfxtp_2_1/a_431_508#
+ sky130_fd_sc_hs__nand2_1_81/a_117_74# sky130_fd_sc_hs__dfrtp_4_73/a_124_78# sky130_fd_sc_hs__dfrtp_4_81/a_1350_392#
+ sky130_fd_sc_hs__dfrtp_4_83/D sky130_fd_sc_hs__dfrtp_4_41/a_124_78# sky130_fd_sc_hs__o21a_1_13/A1
+ sky130_fd_sc_hs__dfrtp_4_63/a_1647_81# sky130_fd_sc_hs__dfrtp_4_11/a_789_463# sky130_fd_sc_hs__dfrtn_1_49/a_507_368#
+ sky130_fd_sc_hs__a21oi_1_97/a_29_368# sky130_fd_sc_hs__dfrbp_1_29/a_796_463# sky130_fd_sc_hs__o21a_1_31/a_320_74#
+ sky130_fd_sc_hs__dfrbp_1_43/a_498_360# sky130_fd_sc_hs__dfstp_2_5/a_398_74# sky130_fd_sc_hs__a2bb2oi_1_1/Y
+ sky130_fd_sc_hs__fa_2_15/a_27_378# sky130_fd_sc_hs__dfrtp_4_59/a_1627_493# sky130_fd_sc_hs__a22o_1_9/a_52_123#
+ sky130_fd_sc_hs__dfxtp_4_3/a_1178_124# sky130_fd_sc_hs__dfrtp_4_37/a_37_78# sky130_fd_sc_hs__dfrtp_4_31/a_834_355#
+ sky130_fd_sc_hs__fa_2_9/a_487_79# sky130_fd_sc_hs__a21oi_1_31/a_29_368# sky130_fd_sc_hs__fa_2_23/a_1119_79#
+ sky130_fd_sc_hs__o211ai_1_5/Y sky130_fd_sc_hs__nand2_1_23/Y sky130_fd_sc_hs__nand2_4_15/a_27_74#
+ sky130_fd_sc_hs__dfrtn_1_19/a_1547_508# sky130_fd_sc_hs__nor2_1_13/Y sky130_fd_sc_hs__dfrbp_1_11/a_1434_74#
+ sky130_fd_sc_hs__a22o_1_19/a_52_123# sky130_fd_sc_hs__dfrtp_4_45/a_1678_395# sky130_fd_sc_hs__o21ai_1_9/Y
+ sky130_fd_sc_hs__dfrbp_1_37/a_1482_48# sky130_fd_sc_hs__dfrbp_1_47/a_1465_471# sky130_fd_sc_hs__o21a_1_63/a_376_387#
+ sky130_fd_sc_hs__nor2_2_1/A sky130_fd_sc_hs__dfrtp_4_79/a_2010_409# sky130_fd_sc_hs__a21oi_1_49/a_117_74#
+ sky130_fd_sc_hs__dfrtp_4_63/a_890_138# sky130_fd_sc_hs__dfxtp_4_3/a_544_485# sky130_fd_sc_hs__fa_2_15/a_701_79#
+ sky130_fd_sc_hs__a21oi_1_17/a_117_74# sky130_fd_sc_hs__dfrtp_4_3/a_313_74# sky130_fd_sc_hs__dfrtn_1_33/a_817_508#
+ sky130_fd_sc_hs__nor2_1_79/a_116_368# sky130_fd_sc_hs__dfrtp_4_39/a_699_463# sky130_fd_sc_hs__dfrtn_1_25/a_300_74#
+ sky130_fd_sc_hs__dfxtp_2_7/a_538_429# sky130_fd_sc_hs__nand4_1_5/a_259_74# sky130_fd_sc_hs__dfrtn_1_41/a_120_74#
+ sky130_fd_sc_hs__fa_2_7/a_484_347# sky130_fd_sc_hs__dfrbp_1_5/D sky130_fd_sc_hs__a21oi_1_61/a_117_74#
+ sky130_fd_sc_hs__dfrtn_1_5/a_120_74# sky130_fd_sc_hs__xnor2_1_9/a_376_368# sky130_fd_sc_hs__dfrtn_1_37/a_1934_94#
+ sky130_fd_sc_hs__dfrbp_1_33/a_1624_74# sky130_fd_sc_hs__inv_2_1/Y sky130_fd_sc_hs__fa_2_21/a_336_347#
+ sky130_fd_sc_hs__dfrtn_1_3/a_922_127# sky130_fd_sc_hs__dfrtn_1_19/a_856_304# sky130_fd_sc_hs__dfrtp_4_31/a_812_138#
+ sky130_fd_sc_hs__a32oi_1_5/A1 sky130_fd_sc_hs__o21a_1_37/X sky130_fd_sc_hs__dfrtn_1_19/a_850_127#
+ sky130_fd_sc_hs__nand2_1_121/a_117_74# sky130_fd_sc_hs__fa_2_17/a_484_347# sky130_fd_sc_hs__dfrbp_1_3/a_1482_48#
+ sky130_fd_sc_hs__dfrtp_4_53/a_1647_81# sky130_fd_sc_hs__dfrbp_1_19/a_796_463# sky130_fd_sc_hs__dfrbp_1_45/Q_N
+ sky130_fd_sc_hs__o22ai_1_1/a_27_74# sky130_fd_sc_hs__a22oi_1_11/a_159_74# sky130_fd_sc_hs__dfxtp_2_9/a_1125_508#
+ sky130_fd_sc_hs__xor2_1_5/a_158_392# sky130_fd_sc_hs__dfrtn_1_27/a_1736_119# sky130_fd_sc_hs__nand2_1_85/a_117_74#
+ sky130_fd_sc_hs__dfrbp_1_37/Q_N sky130_fd_sc_hs__nand3b_2_1/a_206_74# sky130_fd_sc_hs__dfxtp_4_2/a_1178_124#
+ sky130_fd_sc_hs__conb_1_1/a_21_290# sky130_fd_sc_hs__dfrtn_1_9/a_33_74# sky130_fd_sc_hs__dfrbp_1_31/a_706_463#
+ sky130_fd_sc_hs__dfrtn_1_27/a_1266_119# sky130_fd_sc_hs__fa_2_13/a_1119_79# sky130_fd_sc_hs__dfrbp_1_27/Q_N
+ sky130_fd_sc_hs__dfrtp_4_47/a_1350_392# sky130_fd_sc_hs__sdlclkp_4_1/a_119_143#
+ sky130_fd_sc_hs__dfrbp_1_17/a_38_78# sky130_fd_sc_hs__nor2_1_11/Y sky130_fd_sc_hs__dfrtp_4_45/a_124_78#
+ sky130_fd_sc_hs__dfxtp_2_5/a_27_74# sky130_fd_sc_hs__dfrtn_1_5/a_1598_93# sky130_fd_sc_hs__dfrbp_1_19/Q_N
+ sky130_fd_sc_hs__dfrtp_4_85/a_494_366# sky130_fd_sc_hs__o31ai_1_5/Y sky130_fd_sc_hs__dfrbp_1_9/a_1624_74#
+ sky130_fd_sc_hs__dfstp_2_7/a_398_74# sky130_fd_sc_hs__dfxtp_4_9/a_206_368# sky130_fd_sc_hs__o21a_1_13/a_376_387#
+ sky130_fd_sc_hs__sdlclkp_4_1/a_1289_368# sky130_fd_sc_hs__nand2_2_3/Y sky130_fd_sc_hs__o21a_1_53/a_376_387#
+ sky130_fd_sc_hs__o211ai_1_7/a_31_74# sky130_fd_sc_hs__dfrtn_1_5/a_1550_119# sky130_fd_sc_hs__dfrtp_4_53/a_890_138#
+ sky130_fd_sc_hs__fa_2_15/a_1094_347# sky130_fd_sc_hs__fa_2_23/a_27_79# sky130_fd_sc_hs__fa_2_1/a_992_347#
+ sky130_fd_sc_hs__dfxtp_4_2/a_696_458# sky130_fd_sc_hs__dfrtn_1_23/a_817_508# sky130_fd_sc_hs__o21a_1_9/a_376_387#
+ sky130_fd_sc_hs__dfrtn_1_19/a_33_74# sky130_fd_sc_hs__o31ai_1_5/a_114_74# sky130_fd_sc_hs__dfrtp_4_29/a_699_463#
+ sky130_fd_sc_hs__nor2_1_69/a_116_368# sky130_fd_sc_hs__inv_4_73/Y sky130_fd_sc_hs__dfrtp_4_27/a_2010_409#
+ sky130_fd_sc_hs__dfrbp_1_33/a_38_78# sky130_fd_sc_hs__dfrtp_4_67/a_699_463# sky130_fd_sc_hs__dfrtn_1_15/D
+ sky130_fd_sc_hs__dfrbp_1_7/a_706_463# sky130_fd_sc_hs__fa_2_11/a_992_347# sky130_fd_sc_hs__dfrtn_1_27/a_1598_93#
+ sky130_fd_sc_hs__o21ai_1_1/B1 sky130_fd_sc_hs__dfxtp_2_5/a_708_101# sky130_fd_sc_hs__fa_2_9/a_27_79#
+ sky130_fd_sc_hs__dfrtp_4_21/a_37_78# sky130_fd_sc_hs__dfstp_2_1/a_716_456# sky130_fd_sc_hs__dfrtn_1_49/a_856_304#
+ sky130_fd_sc_hs__dfxtp_4_2/a_27_74# sky130_fd_sc_hs__dfxtp_4_7/Q sky130_fd_sc_hs__dfrtn_1_49/a_850_127#
+ sky130_fd_sc_hs__a21oi_1_65/a_117_74# sky130_fd_sc_hs__dfrtn_1_9/a_120_74# sky130_fd_sc_hs__dfrtp_4_37/a_313_74#
+ sky130_fd_sc_hs__fa_2_3/a_683_347# sky130_fd_sc_hs__dfrtp_4_49/a_1827_81# sky130_fd_sc_hs__dfrtn_1_35/a_33_74#
+ sky130_fd_sc_hs__dfrtp_4_83/a_1647_81# sky130_fd_sc_hs__dfrbp_1_43/a_1224_74# sky130_fd_sc_hs__dfrtp_4_89/a_1827_81#
+ sky130_fd_sc_hs__dfrtp_4_5/a_789_463# sky130_fd_sc_hs__dfrbp_1_23/a_498_360# sky130_fd_sc_hs__dfrbp_1_47/a_796_463#
+ sky130_fd_sc_hs__dfrtp_4_57/a_1627_493# sky130_fd_sc_hs__a21oi_1_113/a_29_368# sky130_fd_sc_hs__dfxtp_2_7/a_1125_508#
+ sky130_fd_sc_hs__dfrtn_1_3/a_300_74# sky130_fd_sc_hs__dfrbp_1_5/a_910_118# sky130_fd_sc_hs__dfrbp_1_21/a_706_463#
+ sky130_fd_sc_hs__dfrtp_4_11/a_834_355# sky130_fd_sc_hs__dfrtn_1_17/a_1547_508# sky130_fd_sc_hs__dfrtp_4_1/a_494_366#
+ sky130_fd_sc_hs__nand2_2_15/a_27_74# sky130_fd_sc_hs__o21ai_1_3/a_162_368# sky130_fd_sc_hs__o21a_1_23/a_83_244#
+ sky130_fd_sc_hs__dfrtp_4_75/a_494_366# sky130_fd_sc_hs__dfrtp_4_43/a_1678_395# sky130_fd_sc_hs__fa_2_9/A
+ sky130_fd_sc_hs__a222oi_1_3/a_697_74# sky130_fd_sc_hs__a22oi_1_15/a_159_74# sky130_fd_sc_hs__a22o_1_7/a_132_392#
+ sky130_fd_sc_hs__nand2_1_89/a_117_74# sky130_fd_sc_hs__dfrbp_1_45/a_1465_471# sky130_fd_sc_hs__dfxtp_4_9/a_437_503#
+ sky130_fd_sc_hs__o21a_1_43/a_376_387# sky130_fd_sc_hs__dfrtp_4_77/a_2010_409# sky130_fd_sc_hs__xnor2_1_1/Y
+ sky130_fd_sc_hs__nor2_1_95/B sky130_fd_sc_hs__nand2b_1_3/a_269_74# sky130_fd_sc_hs__dfrtp_4_83/a_890_138#
+ sky130_fd_sc_hs__nand2_1_23/a_117_74# sky130_fd_sc_hs__o21a_1_39/a_320_74# sky130_fd_sc_hs__fa_2_7/B
+ sky130_fd_sc_hs__nor2_1_47/Y sky130_fd_sc_hs__dfrbp_1_11/a_2026_424# sky130_fd_sc_hs__dfsbp_2_1/a_1531_118#
+ sky130_fd_sc_hs__dfrbp_1_29/a_910_118# sky130_fd_sc_hs__dfrtp_4_15/a_124_78# sky130_fd_sc_hs__nor3_1_3/B
+ sky130_fd_sc_hs__dfxtp_4_7/a_735_102# sky130_fd_sc_hs__nor2_1_91/B sky130_fd_sc_hs__dfrtp_4_19/a_699_463#
+ sky130_fd_sc_hs__nor2_1_59/a_116_368# sky130_fd_sc_hs__fa_2_9/a_1094_347# sky130_fd_sc_hs__dfrtp_4_25/a_2010_409#
+ sky130_fd_sc_hs__a21oi_1_39/a_29_368# sky130_fd_sc_hs__a21oi_1_111/a_117_74# sky130_fd_sc_hs__dfrtp_4_25/D
+ sky130_fd_sc_hs__dfrtn_1_17/a_1598_93# sky130_fd_sc_hs__fa_2_1/B sky130_fd_sc_hs__dfxtp_4_9/a_1034_424#
+ sky130_fd_sc_hs__dfrtp_4_11/a_812_138# sky130_fd_sc_hs__a22oi_1_13/Y sky130_fd_sc_hs__inv_4_83/A
+ sky130_fd_sc_hs__nand4_1_3/a_181_74# sky130_fd_sc_hs__maj3_1_1/a_226_384# sky130_fd_sc_hs__a22oi_1_1/a_71_368#
+ sky130_fd_sc_hs__fa_2_7/a_1205_79# sky130_fd_sc_hs__dfrtp_4_9/a_1647_81# sky130_fd_sc_hs__nand2_4_1/a_27_74#
+ sky130_fd_sc_hs__dfrtp_4_79/a_1827_81# sky130_fd_sc_hs__o21a_1_13/X sky130_fd_sc_hs__dfrbp_1_13/a_498_360#
+ sky130_fd_sc_hs__sdlclkp_1_1/a_1238_94# sky130_fd_sc_hs__nor2_1_9/a_116_368# sky130_fd_sc_hs__dfstp_2_4/a_1278_74#
+ sky130_fd_sc_hs__inv_4_5/A sky130_fd_sc_hs__dfrbp_1_11/a_706_463# sky130_fd_sc_hs__a22o_1_21/a_222_392#
+ sky130_fd_sc_hs__a21oi_1_69/a_117_74# sky130_fd_sc_hs__nor2_1_43/Y sky130_fd_sc_hs__fa_2_17/a_1205_79#
+ sky130_fd_sc_hs__dfrtp_4_25/a_494_366# sky130_fd_sc_hs__a211oi_4_1/a_901_368# sky130_fd_sc_hs__a21oi_1_35/a_117_74#
+ sky130_fd_sc_hs__dfrtp_4_65/a_494_366# sky130_fd_sc_hs__dfrtn_1_45/a_922_127# sky130_fd_sc_hs__nand4_2_1/a_515_74#
+ sky130_fd_sc_hs__nor3_1_7/A sky130_fd_sc_hs__o21a_1_33/a_376_387# sky130_fd_sc_hs__dfrbp_1_45/a_1482_48#
+ sky130_fd_sc_hs__dfrbp_1_39/a_832_118# sky130_fd_sc_hs__fa_2_21/B sky130_fd_sc_hs__dfrtn_1_3/a_1550_119#
+ sky130_fd_sc_hs__dfxtp_2_3/a_206_368# sky130_fd_sc_hs__dfrtp_4_9/a_890_138# sky130_fd_sc_hs__fa_2_13/a_1094_347#
+ sky130_fd_sc_hs__dfrtn_1_3/a_714_127# sky130_fd_sc_hs__o21a_1_43/X sky130_fd_sc_hs__fa_2_17/a_487_79#
+ sky130_fd_sc_hs__dfrbp_1_19/a_910_118# sky130_fd_sc_hs__dfrtn_1_41/a_817_508# sky130_fd_sc_hs__a22oi_1_19/a_159_74#
+ sky130_fd_sc_hs__nor2_1_49/a_116_368# sky130_fd_sc_hs__dfrbp_1_29/a_2026_424# sky130_fd_sc_hs__dfrtp_4_47/a_699_463#
+ sky130_fd_sc_hs__o21a_1_71/a_83_244# sky130_fd_sc_hs__dfrtp_4_5/D sky130_fd_sc_hs__nand2b_1_7/a_269_74#
+ sky130_fd_sc_hs__dfrtp_4_87/a_699_463# sky130_fd_sc_hs__nor2_1_123/a_116_368# sky130_fd_sc_hs__a222oi_1_3/a_119_74#
+ sky130_fd_sc_hs__nor2b_1_13/a_278_368# sky130_fd_sc_hs__nand2_1_27/a_117_74# sky130_fd_sc_hs__a22oi_1_13/a_339_74#
+ sky130_fd_sc_hs__nor3_1_7/a_198_368# sky130_fd_sc_hs__a22o_1_9/a_222_392# sky130_fd_sc_hs__dfrbp_1_41/a_1624_74#
+ sky130_fd_sc_hs__dfstp_2_7/a_1521_508# sky130_fd_sc_hs__o31ai_1_7/a_119_368# sky130_fd_sc_hs__inv_4_19/Y
+ sky130_fd_sc_hs__dfrtp_4_87/a_37_78# sky130_fd_sc_hs__nand2_1_71/a_117_74# sky130_fd_sc_hs__dfrtp_4_15/a_37_78#
+ sky130_fd_sc_hs__a21oi_1_115/a_117_74# sky130_fd_sc_hs__dfrtp_4_63/a_124_78# sky130_fd_sc_hs__dfrtp_4_31/a_124_78#
+ sky130_fd_sc_hs__dfrbp_1_23/a_1224_74# sky130_fd_sc_hs__dfrtp_4_69/a_1827_81# sky130_fd_sc_hs__o211ai_1_1/a_311_74#
+ sky130_fd_sc_hs__dfrtn_1_47/a_507_368# sky130_fd_sc_hs__a21oi_1_87/a_29_368# sky130_fd_sc_hs__dfrbp_1_27/a_796_463#
+ sky130_fd_sc_hs__dfrtp_4_55/a_1627_493# sky130_fd_sc_hs__o21a_1_21/a_320_74# sky130_fd_sc_hs__dfrtn_1_25/a_1736_119#
+ sky130_fd_sc_hs__o21ai_1_5/a_27_74# sky130_fd_sc_hs__dfstp_2_7/a_767_384# sky130_fd_sc_hs__a21oi_1_53/a_29_368#
+ sky130_fd_sc_hs__dfrtn_1_25/a_1266_119# sky130_fd_sc_hs__dfrbp_1_41/a_38_78# sky130_fd_sc_hs__dfrtp_4_45/a_1350_392#
+ sky130_fd_sc_hs__dfrbp_1_31/a_319_360# sky130_fd_sc_hs__dfrtp_4_15/a_494_366# sky130_fd_sc_hs__dfrtp_4_5/a_834_355#
+ sky130_fd_sc_hs__a21oi_1_21/a_29_368# sky130_fd_sc_hs__inv_4_93/A sky130_fd_sc_hs__o21ai_1_7/Y
+ sky130_fd_sc_hs__dfrtp_4_55/a_494_366# sky130_fd_sc_hs__dfrtp_4_41/a_1678_395# sky130_fd_sc_hs__dfrtn_1_35/a_922_127#
+ sky130_fd_sc_hs__o21a_1_73/X sky130_fd_sc_hs__dfrtp_4_31/a_37_78# sky130_fd_sc_hs__dfrbp_1_43/a_1465_471#
+ sky130_fd_sc_hs__a21oi_1_3/a_29_368# sky130_fd_sc_hs__o21a_1_23/a_376_387# sky130_fd_sc_hs__dfrtp_4_75/a_2010_409#
+ sky130_fd_sc_hs__fa_2_19/a_1202_368# sky130_fd_sc_hs__dfrtn_1_1/a_1550_119# sky130_fd_sc_hs__fa_2_11/a_1094_347#
+ sky130_fd_sc_hs__dfxtp_4_2/a_544_485# sky130_fd_sc_hs__dfrtn_1_47/a_300_74# sky130_fd_sc_hs__nor2_2_3/a_35_368#
+ sky130_fd_sc_hs__dfrtn_1_31/a_817_508# sky130_fd_sc_hs__dfrbp_1_47/a_910_118# sky130_fd_sc_hs__nor2_1_39/a_116_368#
+ sky130_fd_sc_hs__dfrbp_1_27/a_2026_424# sky130_fd_sc_hs__o21a_1_5/B1 sky130_fd_sc_hs__fa_2_7/a_1094_347#
+ sky130_fd_sc_hs__dfrbp_1_39/Q_N sky130_fd_sc_hs__dfrtp_4_37/a_699_463# sky130_fd_sc_hs__dfrtn_1_15/a_300_74#
+ sky130_fd_sc_hs__dfrtp_4_3/a_699_463# sky130_fd_sc_hs__dfrtp_4_57/a_313_74# sky130_fd_sc_hs__dfrtp_4_77/a_699_463#
+ sky130_fd_sc_hs__dfrtn_1_31/a_120_74# sky130_fd_sc_hs__nor2_1_113/a_116_368# sky130_fd_sc_hs__dfrbp_1_39/a_841_401#
+ sky130_fd_sc_hs__a222o_1_1/a_386_74# sky130_fd_sc_hs__dfrbp_1_7/a_319_360# sky130_fd_sc_hs__dfxtp_4_7/a_1034_424#
+ sky130_fd_sc_hs__fa_2_21/a_992_347# sky130_fd_sc_hs__dfrtn_1_1/a_922_127# sky130_fd_sc_hs__nor2b_1_43/a_278_368#
+ sky130_fd_sc_hs__dfrtn_1_37/a_1598_93# sky130_fd_sc_hs__dfrbp_1_23/a_125_78# sky130_fd_sc_hs__dfrtp_4_5/a_812_138#
+ sky130_fd_sc_hs__nor2b_1_5/a_27_112# sky130_fd_sc_hs__o21a_1_75/a_83_244# sky130_fd_sc_hs__inv_4_115/Y
+ sky130_fd_sc_hs__a211oi_1_3/a_71_368# sky130_fd_sc_hs__nand2_1_51/Y sky130_fd_sc_hs__o21a_1_69/A2
+ sky130_fd_sc_hs__fa_2_1/a_1119_79# sky130_fd_sc_hs__dfstp_2_5/D sky130_fd_sc_hs__dfrbp_1_1/a_1482_48#
+ sky130_fd_sc_hs__a22oi_1_17/a_339_74# sky130_fd_sc_hs__dfrbp_1_13/a_1224_74# sky130_fd_sc_hs__dfrtp_4_59/a_1827_81#
+ sky130_fd_sc_hs__dfxtp_2_11/a_644_504# sky130_fd_sc_hs__dfrbp_1_17/a_796_463# sky130_fd_sc_hs__dfrtp_4_91/a_1678_395#
+ sky130_fd_sc_hs__dfrtp_4_53/a_1627_493# sky130_fd_sc_hs__dfrtp_4_49/a_789_463# sky130_fd_sc_hs__dfxtp_2_5/a_1125_508#
+ sky130_fd_sc_hs__nor2b_1_43/a_27_112# sky130_fd_sc_hs__dfrbp_1_33/a_498_360# sky130_fd_sc_hs__nand2b_4_1/a_31_74#
+ sky130_fd_sc_hs__dfrtp_4_89/a_789_463# sky130_fd_sc_hs__dfsbp_2_1/a_757_401# sky130_fd_sc_hs__nand2_1_75/a_117_74#
+ sky130_fd_sc_hs__a21oi_1_119/a_117_74# sky130_fd_sc_hs__dfrtp_4_67/a_124_78# sky130_fd_sc_hs__dfrbp_1_21/a_319_360#
+ sky130_fd_sc_hs__fa_2_11/a_1119_79# sky130_fd_sc_hs__dfrtn_1_15/a_1547_508# sky130_fd_sc_hs__dfstp_2_5/a_225_74#
+ sky130_fd_sc_hs__nand2_1_41/a_117_74# sky130_fd_sc_hs__fa_2_23/a_683_347# sky130_fd_sc_hs__dfrtp_4_45/a_494_366#
+ sky130_fd_sc_hs__dfrtp_4_35/a_124_78# sky130_fd_sc_hs__a222oi_1_1/a_369_392# sky130_fd_sc_hs__dfrtn_1_3/a_1934_94#
+ sky130_fd_sc_hs__dfrtn_1_25/a_922_127# sky130_fd_sc_hs__o21a_1_25/a_320_74# sky130_fd_sc_hs__dfrtn_1_1/a_33_74#
+ sky130_fd_sc_hs__dfrtp_4_59/a_1678_395# sky130_fd_sc_hs__a22oi_1_9/a_71_368# sky130_fd_sc_hs__o21a_1_67/X
+ sky130_fd_sc_hs__dfrtp_4_7/a_37_78# sky130_fd_sc_hs__dfrbp_1_11/a_38_78# sky130_fd_sc_hs__xnor2_1_9/a_112_119#
+ sky130_fd_sc_hs__dfrbp_1_25/a_1482_48# sky130_fd_sc_hs__dfrtp_4_73/a_2010_409# sky130_fd_sc_hs__inv_4_7/A
+ sky130_fd_sc_hs__nand2_1_3/a_117_74# sky130_fd_sc_hs__a21oi_1_25/a_29_368# sky130_fd_sc_hs__dfrtn_1_5/a_507_368#
+ sky130_fd_sc_hs__xnor2_1_9/A sky130_fd_sc_hs__dfrtn_1_21/a_817_508# sky130_fd_sc_hs__nor2_1_29/a_116_368#
+ sky130_fd_sc_hs__dfrtp_4_71/a_37_78# sky130_fd_sc_hs__xor2_1_3/a_455_87# sky130_fd_sc_hs__a21oi_1_7/a_29_368#
+ sky130_fd_sc_hs__dfrbp_1_17/D sky130_fd_sc_hs__dfrtp_4_23/a_2010_409# sky130_fd_sc_hs__dfrbp_1_9/a_498_360#
+ sky130_fd_sc_hs__nand2_2_9/B sky130_fd_sc_hs__nor2_1_103/a_116_368# sky130_fd_sc_hs__dfxtp_2_7/a_27_74#
+ sky130_fd_sc_hs__nor2b_1_33/a_278_368# sky130_fd_sc_hs__sdlclkp_1_1/a_709_54# sky130_fd_sc_hs__inv_4_95/A
+ sky130_fd_sc_hs__nand2_2_11/Y sky130_fd_sc_hs__dfxtp_2_3/a_708_101# sky130_fd_sc_hs__dfrtn_1_47/a_856_304#
+ sky130_fd_sc_hs__dfrtn_1_47/a_850_127# sky130_fd_sc_hs__a21oi_1_55/a_117_74# sky130_fd_sc_hs__inv_4_29/Y
+ sky130_fd_sc_hs__o22ai_1_7/a_340_368# sky130_fd_sc_hs__dfrtp_4_43/a_1647_81# sky130_fd_sc_hs__a21oi_1_15/Y
+ sky130_fd_sc_hs__dfrtn_1_27/a_507_368# sky130_fd_sc_hs__dfrtn_1_45/a_714_127# sky130_fd_sc_hs__dfxtp_2_3/a_1125_508#
+ sky130_fd_sc_hs__dfrtn_1_23/a_1736_119# sky130_fd_sc_hs__a31oi_1_1/a_136_368# sky130_fd_sc_hs__o21a_1_77/A2
+ sky130_fd_sc_hs__dfrbp_1_27/a_125_78# sky130_fd_sc_hs__xor2_1_1/a_355_368# sky130_fd_sc_hs__dfrtp_4_79/a_789_463#
+ sky130_fd_sc_hs__nor2b_1_9/a_27_112# sky130_fd_sc_hs__a21oi_1_103/a_29_368# sky130_fd_sc_hs__dfrbp_1_1/a_125_78#
+ sky130_fd_sc_hs__dfrtn_1_23/a_1266_119# sky130_fd_sc_hs__nand2_1_115/a_117_74# sky130_fd_sc_hs__dfrtp_4_43/a_1350_392#
+ sky130_fd_sc_hs__nor2_1_29/B sky130_fd_sc_hs__dfrbp_1_11/a_319_360# sky130_fd_sc_hs__dfrtn_1_13/a_1547_508#
+ sky130_fd_sc_hs__dfrbp_1_9/a_38_78# sky130_fd_sc_hs__nand2_2_3/B sky130_fd_sc_hs__nor2_1_19/B
+ sky130_fd_sc_hs__fa_2_13/a_683_347# sky130_fd_sc_hs__xor2_1_11/a_158_392# sky130_fd_sc_hs__dfrtp_4_35/a_494_366#
+ sky130_fd_sc_hs__fa_2_1/a_27_378# sky130_fd_sc_hs__dfrtn_1_15/a_922_127# sky130_fd_sc_hs__dfrtp_4_73/a_494_366#
+ sky130_fd_sc_hs__dfrtp_4_7/a_124_78# sky130_fd_sc_hs__dfrbp_1_39/a_1434_74# sky130_fd_sc_hs__nor2b_1_47/a_27_112#
+ sky130_fd_sc_hs__dfrbp_1_41/a_1465_471# sky130_fd_sc_hs__nor3_1_13/Y sky130_fd_sc_hs__nand2_1_79/a_117_74#
+ sky130_fd_sc_hs__dfrbp_1_15/a_1482_48# sky130_fd_sc_hs__fa_2_17/a_1202_368# sky130_fd_sc_hs__nor2b_1_13/a_27_112#
+ sky130_fd_sc_hs__o31ai_1_7/A1 sky130_fd_sc_hs__dfstp_2_7/a_225_74# sky130_fd_sc_hs__nand2_1_45/a_117_74#
+ sky130_fd_sc_hs__dfrtp_4_43/a_890_138# sky130_fd_sc_hs__dfrtp_4_39/a_124_78# sky130_fd_sc_hs__o211ai_1_9/a_311_74#
+ sky130_fd_sc_hs__nand2_1_13/a_117_74# sky130_fd_sc_hs__o21a_1_29/a_320_74# sky130_fd_sc_hs__dfrtn_1_11/a_817_508#
+ sky130_fd_sc_hs__dfrbp_1_27/a_910_118# sky130_fd_sc_hs__nor2_1_19/a_116_368# sky130_fd_sc_hs__dfrbp_1_25/a_2026_424#
+ sky130_fd_sc_hs__dfrtp_4_9/a_1627_493# sky130_fd_sc_hs__a22oi_1_11/Y sky130_fd_sc_hs__fa_2_5/a_1094_347#
+ sky130_fd_sc_hs__dfrtp_4_21/a_2010_409# sky130_fd_sc_hs__dfrtp_4_17/a_699_463# sky130_fd_sc_hs__nor3_1_1/a_114_368#
+ sky130_fd_sc_hs__dfrtp_4_83/a_124_78# sky130_fd_sc_hs__fa_2_1/a_701_79# sky130_fd_sc_hs__nand2_1_7/a_117_74#
+ sky130_fd_sc_hs__dfrtp_4_57/a_699_463# sky130_fd_sc_hs__nor2_1_97/a_116_368# sky130_fd_sc_hs__o21a_1_73/a_320_74#
+ sky130_fd_sc_hs__a21oi_1_29/a_29_368# sky130_fd_sc_hs__a21oi_1_101/a_117_74# sky130_fd_sc_hs__or2_1_1/B
+ sky130_fd_sc_hs__o31ai_1_7/a_203_368# sky130_fd_sc_hs__dfxtp_4_5/a_1034_424# sky130_fd_sc_hs__nor2b_1_23/a_278_368#
+ sky130_fd_sc_hs__a31oi_1_1/a_223_74# sky130_fd_sc_hs__a21oi_1_73/a_29_368# sky130_fd_sc_hs__nor3_1_15/Y
+ sky130_fd_sc_hs__dfrtp_4_33/a_1647_81# sky130_fd_sc_hs__dfrtp_4_39/a_1827_81# sky130_fd_sc_hs__dfrtn_1_17/a_507_368#
+ sky130_fd_sc_hs__dfrtn_1_35/a_714_127# sky130_fd_sc_hs__dfrbp_1_33/a_1224_74# sky130_fd_sc_hs__dfrtn_1_21/a_1736_119#
+ sky130_fd_sc_hs__dfrbp_1_37/a_796_463# sky130_fd_sc_hs__dfrtp_4_69/a_789_463# sky130_fd_sc_hs__dfstp_2_7/a_2022_94#
+ sky130_fd_sc_hs__dfrtn_1_21/a_1266_119# sky130_fd_sc_hs__o22ai_1_7/a_142_368# sky130_fd_sc_hs__nor2_1_7/a_116_368#
+ sky130_fd_sc_hs__dfstp_2_1/a_1278_74# sky130_fd_sc_hs__dfrtn_1_39/a_120_74# sky130_fd_sc_hs__dfrtp_4_49/a_37_78#
+ sky130_fd_sc_hs__a21oi_1_59/a_117_74# sky130_fd_sc_hs__dfrtp_4_49/a_834_355# sky130_fd_sc_hs__dfrtp_4_89/a_834_355#
+ sky130_fd_sc_hs__xor2_1_5/a_194_125# sky130_fd_sc_hs__nor3_1_11/a_198_368# sky130_fd_sc_hs__dfrtp_4_63/a_494_366#
+ sky130_fd_sc_hs__dfrtp_4_57/a_1678_395# sky130_fd_sc_hs__a21oi_1_107/a_29_368# sky130_fd_sc_hs__dfrtn_1_5/a_856_304#
+ sky130_fd_sc_hs__nand2_1_119/a_117_74# sky130_fd_sc_hs__dfrtn_1_5/a_850_127# sky130_fd_sc_hs__o21a_1_41/X
+ sky130_fd_sc_hs__dfrtp_4_43/a_313_74# sky130_fd_sc_hs__dfrtp_4_33/a_890_138# sky130_fd_sc_hs__a31oi_2_1/a_114_74#
+ sky130_fd_sc_hs__o21a_1_71/a_376_387# sky130_fd_sc_hs__nand2_4_3/a_27_74# sky130_fd_sc_hs__dfxtp_2_11/a_538_429#
+ sky130_fd_sc_hs__fa_2_5/a_27_378# sky130_fd_sc_hs__dfrtn_1_1/a_714_127# sky130_fd_sc_hs__o21a_1_17/a_83_244#
+ sky130_fd_sc_hs__dfrbp_1_17/a_910_118# sky130_fd_sc_hs__dfrtp_4_3/D sky130_fd_sc_hs__nor2_1_47/a_116_368#
+ sky130_fd_sc_hs__dfrbp_1_9/a_1224_74# sky130_fd_sc_hs__dfrtp_4_65/a_37_78# sky130_fd_sc_hs__o21a_1_61/a_83_244#
+ sky130_fd_sc_hs__a22o_1_13/a_230_79# sky130_fd_sc_hs__nor2_1_87/a_116_368# sky130_fd_sc_hs__dfrbp_1_3/a_796_463#
+ sky130_fd_sc_hs__nand4_1_1/a_373_74# sky130_fd_sc_hs__dfstp_2_5/a_1356_74# sky130_fd_sc_hs__dfrbp_1_21/Q_N
+ sky130_fd_sc_hs__nand2_1_17/a_117_74# sky130_fd_sc_hs__dfstp_2_5/a_1521_508# sky130_fd_sc_hs__dfrtn_1_45/a_1934_94#
+ sky130_fd_sc_hs__nor2_1_89/Y sky130_fd_sc_hs__dfxtp_2_11/a_1019_424# sky130_fd_sc_hs__dfrtp_4_49/a_812_138#
+ sky130_fd_sc_hs__dfrtp_4_87/a_124_78# sky130_fd_sc_hs__dfrtn_1_27/a_856_304# sky130_fd_sc_hs__o31ai_1_5/a_119_368#
+ sky130_fd_sc_hs__dfrtn_1_27/a_850_127# sky130_fd_sc_hs__dfrtp_4_89/a_812_138# sky130_fd_sc_hs__fa_2_5/a_701_79#
+ sky130_fd_sc_hs__nand2_1_61/a_117_74# sky130_fd_sc_hs__o21a_1_77/a_320_74# sky130_fd_sc_hs__nor3_1_3/C
+ sky130_fd_sc_hs__dfrtp_4_53/a_124_78# sky130_fd_sc_hs__xnor2_1_9/a_138_385# sky130_fd_sc_hs__dfrtp_4_23/a_1647_81#
+ sky130_fd_sc_hs__dfrtp_4_29/a_1827_81# sky130_fd_sc_hs__dfxtp_2_9/a_695_459# sky130_fd_sc_hs__dfrtn_1_25/a_714_127#
+ sky130_fd_sc_hs__dfrbp_1_5/a_832_118# sky130_fd_sc_hs__dfrtp_4_51/a_1627_493# sky130_fd_sc_hs__dfrtp_4_67/a_1827_81#
+ sky130_fd_sc_hs__dfxtp_2_1/a_1125_508# sky130_fd_sc_hs__dfrtp_4_59/a_789_463# sky130_fd_sc_hs__fa_2_19/a_27_79#
+ sky130_fd_sc_hs__sdlclkp_1_1/a_566_74# sky130_fd_sc_hs__dfrbp_1_41/a_498_360# sky130_fd_sc_hs__dfrtn_1_39/a_1736_119#
+ sky130_fd_sc_hs__sdlclkp_1_1/a_318_74# sky130_fd_sc_hs__o21ai_1_5/Y sky130_fd_sc_hs__dfrtp_4_41/a_1350_392#
+ sky130_fd_sc_hs__a22o_1_11/a_222_392# sky130_fd_sc_hs__dfrtn_1_39/a_1266_119# sky130_fd_sc_hs__dfrtn_1_11/a_1547_508#
+ sky130_fd_sc_hs__clkbuf_8_1/a_125_368# sky130_fd_sc_hs__fa_2_21/a_1119_79# sky130_fd_sc_hs__dfsbp_2_1/a_595_97#
+ sky130_fd_sc_hs__dfrtn_1_21/a_33_74# sky130_fd_sc_hs__dfrtp_4_79/a_834_355# sky130_fd_sc_hs__dfrtp_4_53/a_494_366#
+ sky130_fd_sc_hs__dfrtp_4_19/a_1627_493# sky130_fd_sc_hs__dfrtp_4_71/a_2010_409#
+ sky130_fd_sc_hs__dfxtp_2_11/a_27_74# sky130_fd_sc_hs__dfrtp_4_19/a_37_78# sky130_fd_sc_hs__dfrbp_1_35/a_1482_48#
+ sky130_fd_sc_hs__dfsbp_2_1/a_1453_118# sky130_fd_sc_hs__dfrbp_1_29/a_832_118# sky130_fd_sc_hs__dfrtp_4_23/a_890_138#
+ sky130_fd_sc_hs__dfxtp_4_9/a_651_503# sky130_fd_sc_hs__a21oi_1_93/Y sky130_fd_sc_hs__o21a_1_61/a_376_387#
+ sky130_fd_sc_hs__nor3_1_5/B sky130_fd_sc_hs__dfrbp_1_23/a_2026_424# sky130_fd_sc_hs__dfsbp_2_1/a_731_97#
+ sky130_fd_sc_hs__dfrtp_4_7/a_1627_493# sky130_fd_sc_hs__fa_2_3/a_1094_347# sky130_fd_sc_hs__dfrbp_1_9/a_125_78#
+ sky130_fd_sc_hs__nor2_1_81/Y sky130_fd_sc_hs__nor2_1_77/a_116_368# sky130_fd_sc_hs__dfrtp_4_39/a_2010_409#
+ sky130_fd_sc_hs__dfrtn_1_21/a_120_74# sky130_fd_sc_hs__a21oi_1_41/a_117_74# sky130_fd_sc_hs__fa_2_5/a_484_347#
+ sky130_fd_sc_hs__a211oi_1_3/a_354_368# sky130_fd_sc_hs__fa_2_9/a_27_378# sky130_fd_sc_hs__a32oi_1_1/a_469_74#
+ sky130_fd_sc_hs__o21ai_2_1/a_27_74# sky130_fd_sc_hs__xnor2_1_7/a_376_368# sky130_fd_sc_hs__dfstp_2_4/a_1521_508#
+ sky130_fd_sc_hs__dfrbp_1_31/a_1624_74# sky130_fd_sc_hs__o21a_1_9/a_320_74# sky130_fd_sc_hs__dfrtn_1_35/a_1934_94#
+ sky130_fd_sc_hs__dfrtp_4_91/a_313_74# sky130_fd_sc_hs__fa_2_3/SUM sky130_fd_sc_hs__dfrtn_1_19/a_1550_119#
+ sky130_fd_sc_hs__dfrtn_1_17/a_856_304# sky130_fd_sc_hs__dfrbp_1_13/a_125_78# sky130_fd_sc_hs__a222o_1_1/a_32_74#
+ sky130_fd_sc_hs__dfrtn_1_17/a_850_127# sky130_fd_sc_hs__dfrtp_4_79/a_812_138# sky130_fd_sc_hs__o21a_1_65/a_83_244#
+ sky130_fd_sc_hs__dfrtp_4_91/a_1350_392# sky130_fd_sc_hs__nand2_1_101/a_117_74# sky130_fd_sc_hs__nand4_1_5/a_373_74#
+ sky130_fd_sc_hs__o211ai_1_11/a_116_368# sky130_fd_sc_hs__dfrtp_4_13/a_1647_81# sky130_fd_sc_hs__dfsbp_2_1/a_27_74#
+ sky130_fd_sc_hs__dfrtp_4_19/a_1827_81# sky130_fd_sc_hs__fa_2_23/a_487_79# sky130_fd_sc_hs__dfrtn_1_15/a_714_127#
+ sky130_fd_sc_hs__dfstp_2_7/a_1266_341# sky130_fd_sc_hs__dfstp_2_5/a_612_74# sky130_fd_sc_hs__dfrtn_1_37/a_507_368#
+ sky130_fd_sc_hs__dfrtn_1_9/a_817_508# sky130_fd_sc_hs__nand2_1_97/a_117_74# sky130_fd_sc_hs__conb_1_3/a_165_290#
+ sky130_fd_sc_hs__dfrtp_4_91/a_1647_81# sky130_fd_sc_hs__dfrtp_4_69/a_1627_493# sky130_fd_sc_hs__dfsbp_2_1/a_1001_74#
+ sky130_fd_sc_hs__nor2b_1_33/a_27_112# sky130_fd_sc_hs__nor2_4_1/a_27_368# sky130_fd_sc_hs__fa_2_9/a_701_79#
+ sky130_fd_sc_hs__nand2_1_65/a_117_74# sky130_fd_sc_hs__xor2_1_3/a_158_392# sky130_fd_sc_hs__dfrbp_1_39/a_706_463#
+ sky130_fd_sc_hs__dfrtp_4_59/a_1350_392# sky130_fd_sc_hs__or3b_2_1/a_27_368# sky130_fd_sc_hs__dfrtp_4_69/a_834_355#
+ sky130_fd_sc_hs__dfrtn_1_29/a_1547_508# sky130_fd_sc_hs__dfrtn_1_1/a_1934_94# sky130_fd_sc_hs__dfrtp_4_55/a_1678_395#
+ sky130_fd_sc_hs__dfrtn_1_3/a_1598_93# sky130_fd_sc_hs__dfrtp_4_17/a_1627_493# sky130_fd_sc_hs__a22oi_1_1/a_159_74#
+ sky130_fd_sc_hs__dfrtp_4_83/a_494_366# sky130_fd_sc_hs__o211ai_1_3/a_116_368# sky130_fd_sc_hs__o21a_1_15/a_320_74#
+ sky130_fd_sc_hs__dfrbp_1_5/a_841_401# sky130_fd_sc_hs__dfrbp_1_7/a_1624_74# sky130_fd_sc_hs__fa_2_15/a_1202_368#
+ sky130_fd_sc_hs__dfxtp_4_7/a_206_368# sky130_fd_sc_hs__o21a_1_11/a_376_387# sky130_fd_sc_hs__dfrbp_1_19/a_832_118#
+ sky130_fd_sc_hs__dfrtp_4_89/a_2010_409# sky130_fd_sc_hs__dfrtp_4_13/a_890_138# sky130_fd_sc_hs__a21oi_1_15/a_29_368#
+ sky130_fd_sc_hs__o21a_1_51/a_376_387# sky130_fd_sc_hs__dfrbp_1_15/D sky130_fd_sc_hs__xnor2_1_15/a_376_368#
+ sky130_fd_sc_hs__dfrtp_4_1/a_37_78# sky130_fd_sc_hs__fa_2_9/a_336_347# sky130_fd_sc_hs__o211ai_1_11/a_31_74#
+ sky130_fd_sc_hs__dfrtp_4_91/a_890_138# sky130_fd_sc_hs__dfrbp_1_37/a_910_118# sky130_fd_sc_hs__nor2_1_27/a_116_368#
+ sky130_fd_sc_hs__nand2_2_7/B sky130_fd_sc_hs__nor2_1_67/a_116_368# sky130_fd_sc_hs__dfrtp_4_27/a_699_463#
+ sky130_fd_sc_hs__fa_2_7/COUT sky130_fd_sc_hs__dfrtp_4_59/a_37_78# sky130_fd_sc_hs__dfrtp_4_37/a_2010_409#
+ sky130_fd_sc_hs__dfxtp_4_3/a_1034_424# sky130_fd_sc_hs__dfrbp_1_29/a_841_401# sky130_fd_sc_hs__a22o_1_29/a_132_392#
+ sky130_fd_sc_hs__nor3_1_5/C sky130_fd_sc_hs__fa_2_19/a_336_347# sky130_fd_sc_hs__dfstp_2_1/a_1521_508#
+ sky130_fd_sc_hs__dfrtn_1_25/a_1934_94# sky130_fd_sc_hs__dfrbp_1_21/a_1624_74# sky130_fd_sc_hs__a22o_1_13/a_52_123#
+ sky130_fd_sc_hs__dfrtn_1_5/a_33_74# sky130_fd_sc_hs__dfrtp_4_69/a_812_138# sky130_fd_sc_hs__a21oi_1_77/a_117_74#
+ sky130_fd_sc_hs__dfrbp_1_13/a_38_78# sky130_fd_sc_hs__a21oi_1_45/a_117_74# sky130_fd_sc_hs__a32oi_1_5/a_469_74#
+ sky130_fd_sc_hs__dfrtp_4_17/a_313_74# sky130_fd_sc_hs__fa_2_1/a_683_347# sky130_fd_sc_hs__dfrtp_4_47/a_1827_81#
+ sky130_fd_sc_hs__a21oi_1_11/a_117_74# sky130_fd_sc_hs__dfrtp_4_81/a_1647_81# sky130_fd_sc_hs__dfrtp_4_39/a_789_463#
+ sky130_fd_sc_hs__dfrbp_1_41/a_1224_74# sky130_fd_sc_hs__dfrtp_4_87/a_1827_81# sky130_fd_sc_hs__dfrtp_4_67/a_1627_493#
+ sky130_fd_sc_hs__dfrbp_1_17/a_125_78# sky130_fd_sc_hs__dfrtp_4_73/a_37_78# sky130_fd_sc_hs__dfrbp_1_45/a_796_463#
+ sky130_fd_sc_hs__o22ai_1_7/a_27_74# sky130_fd_sc_hs__o21a_1_69/a_83_244# sky130_fd_sc_hs__o211ai_1_3/a_31_74#
+ sky130_fd_sc_hs__dfrbp_1_3/a_910_118# sky130_fd_sc_hs__nand2_1_105/a_117_74# sky130_fd_sc_hs__dfxtp_2_5/a_644_504#
+ sky130_fd_sc_hs__o21a_1_35/a_83_244# sky130_fd_sc_hs__dfrtp_4_59/a_834_355# sky130_fd_sc_hs__fa_2_11/a_683_347#
+ sky130_fd_sc_hs__dfrtp_4_9/a_494_366# sky130_fd_sc_hs__dfstp_2_7/a_612_74# sky130_fd_sc_hs__dfrtp_4_53/a_1678_395#
+ sky130_fd_sc_hs__o21ai_1_1/a_162_368# sky130_fd_sc_hs__dfrtn_1_13/a_922_127# sky130_fd_sc_hs__nor2b_1_9/Y
+ sky130_fd_sc_hs__nor2b_1_37/a_27_112# sky130_fd_sc_hs__dfrbp_1_3/a_38_78# sky130_fd_sc_hs__a22o_1_5/a_132_392#
+ sky130_fd_sc_hs__nand2_1_69/a_117_74# sky130_fd_sc_hs__dfxtp_4_7/a_437_503# sky130_fd_sc_hs__o21a_1_41/a_376_387#
+ sky130_fd_sc_hs__dfrbp_1_47/a_832_118# sky130_fd_sc_hs__dfrtp_4_29/a_124_78# sky130_fd_sc_hs__fa_2_9/a_1202_368#
+ sky130_fd_sc_hs__dfrtp_4_81/a_890_138# sky130_fd_sc_hs__fa_2_5/a_27_79# sky130_fd_sc_hs__fa_2_1/a_1094_347#
+ sky130_fd_sc_hs__dfrtp_4_5/a_1627_493# sky130_fd_sc_hs__o21a_1_19/a_320_74# sky130_fd_sc_hs__dfxtp_4_5/a_735_102#
+ sky130_fd_sc_hs__a21oi_1_123/a_117_74# sky130_fd_sc_hs__nor2_1_57/a_116_368# sky130_fd_sc_hs__a21oi_1_19/a_29_368#
+ sky130_fd_sc_hs__o21a_1_63/a_320_74# sky130_fd_sc_hs__dfxtp_4_2/a_1034_424# sky130_fd_sc_hs__dfrbp_1_19/a_841_401#
+ sky130_fd_sc_hs__a22o_1_19/a_132_392# sky130_fd_sc_hs__o31ai_1_5/a_203_368# sky130_fd_sc_hs__dfrtn_1_15/a_1934_94#
+ sky130_fd_sc_hs__dfrbp_1_11/a_1624_74# sky130_fd_sc_hs__dfstp_2_4/a_398_74# sky130_fd_sc_hs__dfrtn_1_17/a_1550_119#
+ sky130_fd_sc_hs__nor2b_1_17/Y sky130_fd_sc_hs__a21oi_1_63/a_29_368# sky130_fd_sc_hs__dfrtp_4_59/a_812_138#
+ sky130_fd_sc_hs__dfrtn_1_37/a_856_304# sky130_fd_sc_hs__dfrbp_1_5/a_1434_74# sky130_fd_sc_hs__dfrtn_1_37/a_850_127#
+ sky130_fd_sc_hs__dfxtp_4_7/a_27_74# sky130_fd_sc_hs__nand2_2_11/a_27_74# sky130_fd_sc_hs__dfrtp_4_7/a_1647_81#
+ sky130_fd_sc_hs__nand2_2_1/a_27_74# sky130_fd_sc_hs__fa_2_5/a_1205_79# sky130_fd_sc_hs__dfrtp_4_37/a_1827_81#
+ sky130_fd_sc_hs__dfrtp_4_3/a_1827_81# sky130_fd_sc_hs__dfrtn_1_39/D sky130_fd_sc_hs__dfrtp_4_29/a_789_463#
+ sky130_fd_sc_hs__dfrtp_4_71/a_1647_81# sky130_fd_sc_hs__dfrtp_4_77/a_1827_81# sky130_fd_sc_hs__dfrtn_1_37/a_1736_119#
+ sky130_fd_sc_hs__dfrbp_1_41/Q_N sky130_fd_sc_hs__o31ai_1_1/a_114_74# sky130_fd_sc_hs__dfrtp_4_67/a_789_463#
+ sky130_fd_sc_hs__dfrtn_1_37/a_1266_119# sky130_fd_sc_hs__dfstp_2_1/a_27_74# sky130_fd_sc_hs__dfrbp_1_33/Q_N
+ sky130_fd_sc_hs__dfrtn_1_29/a_120_74# sky130_fd_sc_hs__dfrtp_4_57/a_1350_392# sky130_fd_sc_hs__a32oi_1_9/a_469_74#
+ sky130_fd_sc_hs__dfrtn_1_27/a_1547_508# sky130_fd_sc_hs__dfrbp_1_23/Q_N sky130_fd_sc_hs__dfrtp_4_15/a_1627_493#
+ sky130_fd_sc_hs__dfrbp_1_29/a_1434_74# sky130_fd_sc_hs__a21oi_1_93/a_117_74# sky130_fd_sc_hs__dfrtp_4_43/a_37_78#
+ sky130_fd_sc_hs__dfrtn_1_43/a_922_127# sky130_fd_sc_hs__fa_2_13/a_1202_368# sky130_fd_sc_hs__a211oi_1_3/a_159_74#
+ sky130_fd_sc_hs__nand2_1_109/a_117_74# sky130_fd_sc_hs__dfrtp_4_87/a_2010_409# sky130_fd_sc_hs__o21a_1_31/a_376_387#
+ sky130_fd_sc_hs__dfrbp_1_43/a_1482_48# sky130_fd_sc_hs__dfrtp_4_33/a_313_74# sky130_fd_sc_hs__dfxtp_2_1/a_206_368#
+ sky130_fd_sc_hs__dfrtp_4_7/a_890_138# sky130_fd_sc_hs__dfrbp_1_21/a_2026_424# sky130_fd_sc_hs__dfrtp_4_71/a_890_138#
+ sky130_fd_sc_hs__xnor2_1_3/Y sky130_fd_sc_hs__dfrbp_1_33/a_125_78# sky130_fd_sc_hs__and2_2_3/a_31_74#
+ sky130_fd_sc_hs__dfrbp_1_39/a_2026_424# sky130_fd_sc_hs__nor3_1_1/A sky130_fd_sc_hs__dfrbp_1_1/a_796_463#
+ sky130_fd_sc_hs__o21a_1_51/a_83_244# sky130_fd_sc_hs__dfrtp_4_85/a_699_463# sky130_fd_sc_hs__dfstp_2_4/a_1356_74#
+ sky130_fd_sc_hs__dfrbp_1_47/a_841_401# sky130_fd_sc_hs__nor2_1_121/a_116_368# sky130_fd_sc_hs__nor3_1_5/a_198_368#
+ sky130_fd_sc_hs__a22oi_1_9/a_159_74# sky130_fd_sc_hs__a22o_1_7/a_222_392# sky130_fd_sc_hs__dfrtp_4_9/a_1678_395#
+ sky130_fd_sc_hs__dfrtn_1_45/a_1598_93# sky130_fd_sc_hs__dfrtp_4_77/a_124_78# sky130_fd_sc_hs__nand2_1_51/a_117_74#
+ sky130_fd_sc_hs__o21a_1_67/a_320_74# sky130_fd_sc_hs__a22oi_1_3/a_339_74# sky130_fd_sc_hs__dfrtp_4_21/a_1647_81#
+ sky130_fd_sc_hs__dfrbp_1_9/a_1465_471# sky130_fd_sc_hs__dfxtp_2_7/a_695_459# sky130_fd_sc_hs__dfrtp_4_11/a_124_78#
+ sky130_fd_sc_hs__dfrtp_4_19/a_789_463# sky130_fd_sc_hs__dfrtp_4_61/a_1647_81# sky130_fd_sc_hs__fa_2_17/a_27_378#
+ sky130_fd_sc_hs__a21oi_1_67/a_29_368# sky130_fd_sc_hs__dfrbp_1_25/a_796_463# sky130_fd_sc_hs__nor2_1_57/B
+ sky130_fd_sc_hs__nand2b_1_1/a_27_112# sky130_fd_sc_hs__dfrtp_4_67/a_37_78# sky130_fd_sc_hs__a21oi_1_33/a_29_368#
+ sky130_fd_sc_hs__sdlclkp_4_1/a_744_74# sky130_fd_sc_hs__dfrtp_4_39/a_834_355# sky130_fd_sc_hs__dfrbp_1_39/a_319_360#
+ sky130_fd_sc_hs__a32oi_1_3/a_391_74# sky130_fd_sc_hs__fa_2_13/a_27_79# sky130_fd_sc_hs__nand4_1_5/D
+ sky130_fd_sc_hs__dfrbp_1_19/a_1434_74# sky130_fd_sc_hs__dfrtn_1_33/a_922_127# sky130_fd_sc_hs__fa_2_11/a_1202_368#
+ sky130_fd_sc_hs__fa_2_7/SUM sky130_fd_sc_hs__xor2_1_11/a_194_125# sky130_fd_sc_hs__o21a_1_21/a_376_387#
+ sky130_fd_sc_hs__dfrbp_1_27/a_832_118# sky130_fd_sc_hs__dfsbp_2_1/a_706_463# sky130_fd_sc_hs__fa_2_23/a_1094_347#
+ sky130_fd_sc_hs__fa_2_17/a_701_79# sky130_fd_sc_hs__dfrtp_4_21/a_890_138# sky130_fd_sc_hs__fa_2_7/a_1202_368#
+ sky130_fd_sc_hs__dfsbp_2_1/a_1261_74# sky130_fd_sc_hs__dfxtp_2_11/a_1172_124# sky130_fd_sc_hs__dfrtp_4_61/a_890_138#
+ sky130_fd_sc_hs__dfrtp_4_5/a_313_74# sky130_fd_sc_hs__nand2_4_9/A sky130_fd_sc_hs__nor3_1_7/Y
+ sky130_fd_sc_hs__a21oi_1_97/a_117_74# sky130_fd_sc_hs__dfrtp_4_83/a_37_78# sky130_fd_sc_hs__dfrtp_4_57/D
+ sky130_fd_sc_hs__dfrtn_1_27/a_300_74# sky130_fd_sc_hs__nor2_1_37/a_116_368# sky130_fd_sc_hs__dfrbp_1_45/a_910_118#
+ sky130_fd_sc_hs__dfrtp_4_35/a_2010_409# sky130_fd_sc_hs__dfrtn_1_45/a_120_74# sky130_fd_sc_hs__nor2_1_75/a_116_368#
+ sky130_fd_sc_hs__dfxtp_2_5/a_538_429# sky130_fd_sc_hs__dfrtn_1_7/a_120_74# sky130_fd_sc_hs__dfrtp_4_1/a_699_463#
+ sky130_fd_sc_hs__dfrtn_1_11/a_120_74# sky130_fd_sc_hs__dfrtp_4_75/a_699_463# sky130_fd_sc_hs__a21oi_1_31/a_117_74#
+ sky130_fd_sc_hs__dfrtn_1_25/a_33_74# sky130_fd_sc_hs__nor2_1_111/a_116_368# sky130_fd_sc_hs__o21ai_1_1/a_27_74#
+ sky130_fd_sc_hs__dfrbp_1_37/a_125_78# sky130_fd_sc_hs__dfrtn_1_35/a_1598_93# sky130_fd_sc_hs__nor2b_1_41/a_278_368#
+ sky130_fd_sc_hs__dfrtp_4_81/a_313_74# sky130_fd_sc_hs__dfrtp_4_39/a_812_138# sky130_fd_sc_hs__dfrtn_1_1/a_300_74#
+ sky130_fd_sc_hs__o21a_1_55/a_83_244# sky130_fd_sc_hs__fa_2_15/a_484_347# sky130_fd_sc_hs__dfrtp_4_17/a_1827_81#
+ sky130_fd_sc_hs__dfstp_2_5/a_1266_341# sky130_fd_sc_hs__fa_2_13/a_487_79# sky130_fd_sc_hs__dfxtp_4_9/a_1226_296#
+ sky130_fd_sc_hs__dfrtn_1_13/a_714_127# sky130_fd_sc_hs__nor2_1_15/B sky130_fd_sc_hs__dfrtp_4_51/a_1647_81#
+ sky130_fd_sc_hs__dfrtp_4_57/a_1827_81# sky130_fd_sc_hs__dfrtp_4_65/a_1627_493# sky130_fd_sc_hs__dfrbp_1_9/Q_N
+ sky130_fd_sc_hs__dfrtn_1_7/a_817_508# sky130_fd_sc_hs__dfrbp_1_15/a_796_463# sky130_fd_sc_hs__dfrtn_1_35/a_1736_119#
+ sky130_fd_sc_hs__nor3_1_15/B sky130_fd_sc_hs__dfrtp_4_47/a_789_463# sky130_fd_sc_hs__nor2b_1_23/a_27_112#
+ sky130_fd_sc_hs__dfrbp_1_31/a_498_360# sky130_fd_sc_hs__dfrtn_1_35/a_1266_119# sky130_fd_sc_hs__dfrtp_4_87/a_789_463#
+ sky130_fd_sc_hs__inv_4_27/Y sky130_fd_sc_hs__dfrtp_4_55/a_1350_392# sky130_fd_sc_hs__nand2_1_55/a_117_74#
+ sky130_fd_sc_hs__dfrbp_1_47/a_38_78# sky130_fd_sc_hs__dfrtp_4_29/a_834_355# sky130_fd_sc_hs__dfrtp_4_47/a_124_78#
+ sky130_fd_sc_hs__a22oi_1_7/a_339_74# sky130_fd_sc_hs__dfrtp_4_67/a_834_355# sky130_fd_sc_hs__fa_2_21/a_683_347#
+ sky130_fd_sc_hs__o21a_1_37/a_320_74# sky130_fd_sc_hs__dfrtp_4_51/a_1678_395# sky130_fd_sc_hs__dfrtp_4_43/a_494_366#
+ sky130_fd_sc_hs__dfrtn_1_23/a_922_127# sky130_fd_sc_hs__dfrtn_1_1/a_1598_93# sky130_fd_sc_hs__a22oi_1_23/a_71_368#
+ sky130_fd_sc_hs__dfrbp_1_47/a_1434_74# sky130_fd_sc_hs__nand2b_1_5/a_27_112# sky130_fd_sc_hs__dfrtp_4_85/a_2010_409#
+ sky130_fd_sc_hs__a21oi_1_37/a_29_368# sky130_fd_sc_hs__dfrbp_1_23/a_1482_48# sky130_fd_sc_hs__xnor2_1_7/a_112_119#
+ sky130_fd_sc_hs__dfrbp_1_17/a_832_118# sky130_fd_sc_hs__a32oi_1_7/a_391_74# sky130_fd_sc_hs__dfrtp_4_51/a_890_138#
+ sky130_fd_sc_hs__dfrtp_4_3/a_1627_493# sky130_fd_sc_hs__a21oi_1_83/a_29_368# sky130_fd_sc_hs__dfrtp_4_19/a_1678_395#
+ sky130_fd_sc_hs__nand3b_2_1/a_27_94# sky130_fd_sc_hs__dfrtn_1_3/a_507_368# sky130_fd_sc_hs__fa_2_9/a_992_347#
+ sky130_fd_sc_hs__dfxtp_4_9/a_696_458# sky130_fd_sc_hs__o21a_1_7/a_376_387# sky130_fd_sc_hs__dfxtp_4_2/Q
+ sky130_fd_sc_hs__a32oi_1_3/a_27_368# sky130_fd_sc_hs__dfrtp_4_25/a_699_463# sky130_fd_sc_hs__nor2b_1_9/a_278_368#
+ sky130_fd_sc_hs__dfrbp_1_7/a_498_360# sky130_fd_sc_hs__or3b_2_1/a_190_260# sky130_fd_sc_hs__dfrtp_4_65/a_699_463#
+ sky130_fd_sc_hs__nor2_1_101/a_116_368# sky130_fd_sc_hs__dfrbp_1_27/a_841_401# sky130_fd_sc_hs__dfrtp_4_9/a_313_74#
+ sky130_fd_sc_hs__dfrbp_1_5/a_706_463# sky130_fd_sc_hs__fa_2_19/a_992_347# sky130_fd_sc_hs__dfrtn_1_15/a_1550_119#
+ sky130_fd_sc_hs__dfrtp_4_7/a_1678_395# sky130_fd_sc_hs__nor2b_1_31/a_278_368# sky130_fd_sc_hs__dfrtn_1_25/a_1598_93#
+ sky130_fd_sc_hs__dfrtp_4_29/a_812_138# sky130_fd_sc_hs__dfrtn_1_49/a_120_74# sky130_fd_sc_hs__maj3_1_3/a_403_136#
+ sky130_fd_sc_hs__dfrtp_4_67/a_812_138# sky130_fd_sc_hs__dfxtp_2_1/a_708_101# sky130_fd_sc_hs__dfstp_2_5/a_781_74#
+ sky130_fd_sc_hs__dfrbp_1_7/a_1465_471# sky130_fd_sc_hs__dfstp_2_4/a_1266_341# sky130_fd_sc_hs__o22ai_1_5/a_340_368#
+ sky130_fd_sc_hs__dfrtp_4_41/a_1647_81# sky130_fd_sc_hs__dfrtp_4_63/a_1627_493# sky130_fd_sc_hs__dfrtn_1_43/a_300_74#
+ sky130_fd_sc_hs__dfrtn_1_43/a_714_127# sky130_fd_sc_hs__a21oi_1_117/a_29_368# sky130_fd_sc_hs__dfrtp_4_37/a_789_463#
+ sky130_fd_sc_hs__dfrtp_4_85/a_313_74# sky130_fd_sc_hs__dfrtp_4_3/a_789_463# sky130_fd_sc_hs__dfrbp_1_21/a_498_360#
+ sky130_fd_sc_hs__nor3_1_15/a_114_368# sky130_fd_sc_hs__dfrtp_4_77/a_789_463# sky130_fd_sc_hs__xnor2_1_15/a_112_119#
+ sky130_fd_sc_hs__o21a_1_59/a_83_244# sky130_fd_sc_hs__dfrtp_4_53/a_1350_392# sky130_fd_sc_hs__dfrbp_1_29/a_706_463#
+ sky130_fd_sc_hs__dfrtp_4_19/a_834_355# sky130_fd_sc_hs__dfrbp_1_1/a_910_118# sky130_fd_sc_hs__dfxtp_2_3/a_644_504#
+ sky130_fd_sc_hs__dfrtn_1_25/a_1547_508# sky130_fd_sc_hs__a21oi_1_91/Y sky130_fd_sc_hs__dfrtp_4_13/a_1627_493#
+ sky130_fd_sc_hs__dfrtp_4_33/a_494_366# sky130_fd_sc_hs__dfstp_2_7/a_1489_118# sky130_fd_sc_hs__dfrtp_4_69/a_1678_395#
+ sky130_fd_sc_hs__nor2b_1_27/a_27_112# sky130_fd_sc_hs__dfrtn_1_7/a_33_74# sky130_fd_sc_hs__a22o_1_23/a_230_79#
+ sky130_fd_sc_hs__inv_4_25/Y sky130_fd_sc_hs__nand2_1_59/a_117_74# sky130_fd_sc_hs__dfrbp_1_13/a_1482_48#
+ sky130_fd_sc_hs__dfxtp_2_3/a_27_74# sky130_fd_sc_hs__fa_2_21/a_1094_347# sky130_fd_sc_hs__inv_4_57/Y
+ sky130_fd_sc_hs__fa_2_5/a_1202_368# sky130_fd_sc_hs__dfrtp_4_41/a_890_138# sky130_fd_sc_hs__dfrtp_4_19/a_124_78#
+ sky130_fd_sc_hs__dfrtp_4_17/a_1678_395# sky130_fd_sc_hs__dfrbp_1_37/a_2026_424#
+ sky130_fd_sc_hs__or2_1_3/a_152_368# sky130_fd_sc_hs__dfrbp_1_25/a_910_118# sky130_fd_sc_hs__o21a_1_55/X
+ sky130_fd_sc_hs__nor2_1_17/a_116_368# sky130_fd_sc_hs__dfrtp_4_33/a_2010_409# sky130_fd_sc_hs__dfxtp_2_9/a_1019_424#
+ sky130_fd_sc_hs__nand2b_1_9/a_27_112# sky130_fd_sc_hs__dfrtp_4_77/a_37_78# sky130_fd_sc_hs__nor2b_1_5/Y
+ sky130_fd_sc_hs__a21oi_1_113/a_117_74# sky130_fd_sc_hs__dfrtp_4_15/a_699_463# sky130_fd_sc_hs__o211ai_1_5/a_31_74#
+ sky130_fd_sc_hs__dfrtp_4_55/a_699_463# sky130_fd_sc_hs__nor2_1_95/a_116_368# sky130_fd_sc_hs__o21a_1_53/a_320_74#
+ sky130_fd_sc_hs__dfrbp_1_17/a_841_401# sky130_fd_sc_hs__nor2b_1_15/Y sky130_fd_sc_hs__dfstp_2_7/a_1057_118#
+ sky130_fd_sc_hs__dfrtn_1_13/a_1550_119# sky130_fd_sc_hs__dfrtn_1_13/a_1934_94# sky130_fd_sc_hs__dfrtn_1_15/a_1598_93#
+ sky130_fd_sc_hs__nor2b_1_21/a_278_368# sky130_fd_sc_hs__dfrbp_1_17/Q_N sky130_fd_sc_hs__dfrtp_4_19/a_812_138#
+ sky130_fd_sc_hs__a32oi_1_7/a_27_368# sky130_fd_sc_hs__dfstp_2_1/a_1266_341# sky130_fd_sc_hs__dfxtp_4_7/a_1226_296#
+ sky130_fd_sc_hs__dfrtp_4_31/a_1647_81# sky130_fd_sc_hs__dfrtn_1_33/a_1736_119# sky130_fd_sc_hs__dfrtn_1_33/a_714_127#
+ sky130_fd_sc_hs__dfrbp_1_31/a_1224_74# sky130_fd_sc_hs__dfrbp_1_11/a_498_360# sky130_fd_sc_hs__dfrtn_1_33/a_1266_119#
+ sky130_fd_sc_hs__dfrbp_1_35/a_796_463# sky130_fd_sc_hs__o22ai_1_5/a_142_368# sky130_fd_sc_hs__dfrbp_1_19/a_706_463#
+ sky130_fd_sc_hs__dfrtn_1_19/a_120_74# sky130_fd_sc_hs__dfstp_2_7/a_781_74# sky130_fd_sc_hs__a21oi_1_39/a_117_74#
+ sky130_fd_sc_hs__a2bb2oi_1_1/a_399_368# sky130_fd_sc_hs__dfrtp_4_47/a_834_355# sky130_fd_sc_hs__o21ai_1_11/a_162_368#
+ sky130_fd_sc_hs__fa_2_15/a_1205_79# sky130_fd_sc_hs__o21a_1_3/a_83_244# sky130_fd_sc_hs__dfrtp_4_23/a_494_366#
+ sky130_fd_sc_hs__dfrtp_4_87/a_834_355# sky130_fd_sc_hs__xor2_1_3/a_194_125# sky130_fd_sc_hs__dfrtp_4_67/a_1678_395#
+ sky130_fd_sc_hs__dfrtp_4_89/a_313_74# sky130_fd_sc_hs__dfrbp_1_27/a_1434_74# sky130_fd_sc_hs__dfrtn_1_41/a_922_127#
+ sky130_fd_sc_hs__dfrtn_1_13/a_300_74# sky130_fd_sc_hs__dfrtp_4_83/a_2010_409# sky130_fd_sc_hs__dfrtn_1_3/a_856_304#
+ sky130_fd_sc_hs__dfrtn_1_3/a_850_127# sky130_fd_sc_hs__nand2_2_13/a_27_74# sky130_fd_sc_hs__dfrbp_1_37/a_832_118#
+ sky130_fd_sc_hs__dfrtp_4_23/a_313_74# sky130_fd_sc_hs__dfrtp_4_31/a_890_138# sky130_fd_sc_hs__dfrtp_4_1/a_1627_493#
+ sky130_fd_sc_hs__dfrbp_1_15/a_910_118# sky130_fd_sc_hs__dfxtp_2_7/a_1019_424# sky130_fd_sc_hs__nor2b_1_3/a_27_112#
+ sky130_fd_sc_hs__a22o_1_27/a_230_79# sky130_fd_sc_hs__dfrbp_1_7/a_1224_74# sky130_fd_sc_hs__dfrtp_4_45/a_699_463#
+ sky130_fd_sc_hs__o21a_1_41/a_83_244# sky130_fd_sc_hs__nor2_1_85/a_116_368# sky130_fd_sc_hs__dfrtp_4_9/a_1350_392#
+ sky130_fd_sc_hs__dfxtp_2_11/a_1217_314# sky130_fd_sc_hs__dfstp_2_1/a_1356_74# sky130_fd_sc_hs__nand4_2_1/a_27_74#
+ sky130_fd_sc_hs__dfrtp_4_3/a_124_78# sky130_fd_sc_hs__dfrtp_4_5/a_1678_395# sky130_fd_sc_hs__nor2b_1_11/a_278_368#
+ sky130_fd_sc_hs__dfrtn_1_43/a_1934_94# sky130_fd_sc_hs__dfrtp_4_77/D sky130_fd_sc_hs__dfrtp_4_47/a_812_138#
+ sky130_fd_sc_hs__dfxtp_2_9/a_431_508# sky130_fd_sc_hs__dfrtp_4_87/a_812_138# sky130_fd_sc_hs__dfstp_2_4/a_225_74#
+ sky130_fd_sc_hs__o21a_1_57/a_320_74# sky130_fd_sc_hs__a32oi_1_3/a_119_74# sky130_fd_sc_hs__xnor2_1_7/a_138_385#
+ sky130_fd_sc_hs__dfrtp_4_27/a_1827_81# sky130_fd_sc_hs__dfrtn_1_23/a_714_127# sky130_fd_sc_hs__dfrtn_1_31/a_1736_119#
+ sky130_fd_sc_hs__dfrbp_1_3/a_832_118# sky130_fd_sc_hs__dfrtp_4_17/a_789_463# sky130_fd_sc_hs__a2bb2oi_1_1/a_488_74#
+ sky130_fd_sc_hs__dfrbp_1_21/a_1224_74# sky130_fd_sc_hs__dfrtn_1_45/a_507_368# sky130_fd_sc_hs__a21oi_1_57/a_29_368#
+ sky130_fd_sc_hs__dfrtn_1_31/a_1266_119# sky130_fd_sc_hs__dfrtp_4_57/a_789_463# sky130_fd_sc_hs__dfrtn_1_23/a_1547_508#
+ sky130_fd_sc_hs__dfrbp_1_47/a_706_463# sky130_fd_sc_hs__dfrtp_4_37/a_834_355# sky130_fd_sc_hs__dfrtp_4_11/a_1627_493#
+ sky130_fd_sc_hs__dfrtp_4_13/a_494_366# sky130_fd_sc_hs__dfrtp_4_3/a_834_355# sky130_fd_sc_hs__dfrtp_4_77/a_834_355#
+ sky130_fd_sc_hs__dfrtp_4_61/a_37_78# sky130_fd_sc_hs__dfrbp_1_17/a_1434_74# sky130_fd_sc_hs__dfrtn_1_31/a_922_127#
+ sky130_fd_sc_hs__dfrtp_4_91/a_494_366# sky130_fd_sc_hs__a2bb2oi_1_1/a_126_112# sky130_fd_sc_hs__xnor2_1_3/a_293_74#
+ sky130_fd_sc_hs__fa_2_3/a_1202_368# sky130_fd_sc_hs__dfrbp_1_33/a_1482_48# sky130_fd_sc_hs__dfxtp_4_7/a_651_503#
+ sky130_fd_sc_hs__o21a_1_7/a_83_244# sky130_fd_sc_hs__a22o_1_23/a_52_123# sky130_fd_sc_hs__dfrtp_4_15/a_1678_395#
+ sky130_fd_sc_hs__dfxtp_4_9/a_544_485# sky130_fd_sc_hs__dfrbp_1_35/a_2026_424# sky130_fd_sc_hs__dfrtp_4_31/a_2010_409#
+ sky130_fd_sc_hs__a21oi_1_87/a_117_74# sky130_fd_sc_hs__dfrtn_1_39/a_817_508# sky130_fd_sc_hs__dfrbp_1_19/a_1465_471#
+ sky130_fd_sc_hs__a222oi_1_1/a_461_74# sky130_fd_sc_hs__dfrtn_1_17/a_300_74# sky130_fd_sc_hs__dfrtn_1_35/a_120_74#
+ sky130_fd_sc_hs__dfrtp_4_49/a_2010_409# sky130_fd_sc_hs__a21oi_1_53/a_117_74# sky130_fd_sc_hs__dfrtp_4_35/a_699_463#
+ sky130_fd_sc_hs__dfxtp_2_3/a_538_429# sky130_fd_sc_hs__xnor2_1_15/a_138_385# sky130_fd_sc_hs__dfrtp_4_27/a_313_74#
+ sky130_fd_sc_hs__dfrtp_4_73/a_699_463# sky130_fd_sc_hs__fa_2_3/a_484_347# sky130_fd_sc_hs__a21oi_1_21/a_117_74#
+ sky130_fd_sc_hs__a211oi_1_1/a_354_368# sky130_fd_sc_hs__dfrtn_1_11/a_1550_119# sky130_fd_sc_hs__o2bb2ai_1_1/a_397_74#
+ sky130_fd_sc_hs__dfrbp_1_37/a_841_401# sky130_fd_sc_hs__o21ai_2_1/a_116_368# sky130_fd_sc_hs__dfrbp_1_39/a_1624_74#
+ sky130_fd_sc_hs__dfrbp_1_5/a_319_360# sky130_fd_sc_hs__xnor2_1_5/a_376_368# sky130_fd_sc_hs__dfrtn_1_33/a_1934_94#
+ sky130_fd_sc_hs__dfrtp_4_71/a_313_74# sky130_fd_sc_hs__dfrtp_4_37/a_812_138# sky130_fd_sc_hs__dfrtn_1_19/D
+ sky130_fd_sc_hs__a21oi_1_3/a_117_74# sky130_fd_sc_hs__dfrtp_4_3/a_812_138# sky130_fd_sc_hs__dfrbp_1_25/a_38_78#
+ sky130_fd_sc_hs__dfrtp_4_77/a_812_138# sky130_fd_sc_hs__o21a_1_45/a_83_244# sky130_fd_sc_hs__dfrbp_1_5/a_1465_471#
+ sky130_fd_sc_hs__dfxtp_4_5/a_1226_296# sky130_fd_sc_hs__dfrtp_4_11/a_1647_81# sky130_fd_sc_hs__fa_2_9/a_1119_79#
+ sky130_fd_sc_hs__dfrtp_4_61/a_1627_493# sky130_fd_sc_hs__dfrbp_1_9/a_1482_48# sky130_fd_sc_hs__o21a_1_11/a_83_244#
+ sky130_fd_sc_hs__nor2b_2_1/a_27_392# sky130_fd_sc_hs__o21a_1_1/a_320_74# sky130_fd_sc_hs__dfrbp_1_11/a_1224_74#
+ sky130_fd_sc_hs__dfrtn_1_35/a_507_368# sky130_fd_sc_hs__conb_1_1/a_165_290# sky130_fd_sc_hs__dfrtp_4_51/a_1350_392#
+ sky130_fd_sc_hs__dfrtn_1_21/a_1547_508# sky130_fd_sc_hs__xor2_1_1/a_158_392# sky130_fd_sc_hs__dfrtp_4_37/a_124_78#
+ sky130_fd_sc_hs__dfrbp_1_29/a_319_360# sky130_fd_sc_hs__a32oi_1_7/a_119_74# sky130_fd_sc_hs__fa_2_19/a_1119_79#
+ sky130_fd_sc_hs__dfrtn_1_27/a_33_74# sky130_fd_sc_hs__o21a_1_27/a_320_74# sky130_fd_sc_hs__dfrtp_4_29/a_1627_493#
+ sky130_fd_sc_hs__dfstp_2_7/a_1596_118# sky130_fd_sc_hs__dfrtn_1_21/a_922_127# sky130_fd_sc_hs__dfrtp_4_81/a_494_366#
+ sky130_fd_sc_hs__o211ai_1_1/a_116_368# sky130_fd_sc_hs__dfrtp_4_81/a_2010_409# sky130_fd_sc_hs__dfrbp_1_3/a_841_401#
+ sky130_fd_sc_hs__a22oi_1_13/a_71_368# sky130_fd_sc_hs__dfxtp_4_5/a_206_368# sky130_fd_sc_hs__dfrtp_4_19/a_1350_392#
+ sky130_fd_sc_hs__dfrtp_4_79/D sky130_fd_sc_hs__dfrtp_4_11/a_890_138# sky130_fd_sc_hs__xnor2_1_13/a_376_368#
+ sky130_fd_sc_hs__fa_2_23/a_27_378# sky130_fd_sc_hs__fa_2_7/a_336_347# sky130_fd_sc_hs__dfrtn_1_1/a_507_368#
+ sky130_fd_sc_hs__dfrbp_1_17/a_1465_471# sky130_fd_sc_hs__dfrtn_1_29/a_817_508# sky130_fd_sc_hs__dfstp_2_7/a_1566_92#
+ sky130_fd_sc_hs__dfrbp_1_35/a_910_118# sky130_fd_sc_hs__dfrtp_4_7/a_1350_392# sky130_fd_sc_hs__nor2_1_65/a_116_368#
+ sky130_fd_sc_hs__xnor2_1_7/a_293_74# sky130_fd_sc_hs__dfrtn_1_43/a_33_74# sky130_fd_sc_hs__dfrtp_4_63/a_699_463#
+ sky130_fd_sc_hs__a22o_1_27/a_52_123# sky130_fd_sc_hs__maj3_1_3/a_406_384# sky130_fd_sc_hs__a22o_1_27/a_132_392#
+ sky130_fd_sc_hs__fa_2_17/a_336_347# sky130_fd_sc_hs__dfrtn_1_23/a_1934_94# sky130_fd_sc_hs__dfrtn_1_29/a_1550_119#
+ sky130_fd_sc_hs__maj3_1_1/a_403_136# sky130_fd_sc_hs__dfrtn_1_45/a_856_304# sky130_fd_sc_hs__fa_2_23/a_701_79#
+ sky130_fd_sc_hs__dfrtn_1_45/a_850_127# sky130_fd_sc_hs__a21oi_1_25/a_117_74# sky130_fd_sc_hs__sdlclkp_1_1/a_667_80#
+ sky130_fd_sc_hs__dfrtn_1_33/a_300_74# sky130_fd_sc_hs__dfrtn_1_25/a_507_368# sky130_fd_sc_hs__dfrtp_4_79/a_1627_493#
+ sky130_fd_sc_hs__dfrtn_1_41/a_714_127# sky130_fd_sc_hs__dfrbp_1_5/a_125_78# sky130_fd_sc_hs__dfrtn_1_49/a_1736_119#
+ sky130_fd_sc_hs__dfrtp_4_75/a_313_74# sky130_fd_sc_hs__dfrbp_1_47/Q_N sky130_fd_sc_hs__dfrtp_4_85/a_1827_81#
+ sky130_fd_sc_hs__xor2_1_9/a_355_368# sky130_fd_sc_hs__a21oi_1_7/a_117_74# sky130_fd_sc_hs__dfrbp_1_43/a_796_463#
+ sky130_fd_sc_hs__dfrtn_1_49/a_1266_119# sky130_fd_sc_hs__o21a_1_49/a_83_244# sky130_fd_sc_hs__dfrtp_4_69/a_1350_392#
+ sky130_fd_sc_hs__dfrbp_1_27/a_706_463# sky130_fd_sc_hs__dfrtp_4_17/a_834_355# sky130_fd_sc_hs__dfrbp_1_19/a_319_360#
+ sky130_fd_sc_hs__a22o_1_3/a_230_79# sky130_fd_sc_hs__dfrtn_1_39/a_1547_508# sky130_fd_sc_hs__dfrtp_4_57/a_834_355#
+ sky130_fd_sc_hs__dfstp_2_5/a_1489_118# sky130_fd_sc_hs__dfrbp_1_41/a_125_78# sky130_fd_sc_hs__dfrtp_4_65/a_1678_395#
+ sky130_fd_sc_hs__dfrtp_4_7/a_494_366# sky130_fd_sc_hs__o21a_1_5/a_320_74# sky130_fd_sc_hs__nor2b_1_49/a_27_112#
+ sky130_fd_sc_hs__dfrtn_1_11/a_922_127# sky130_fd_sc_hs__dfrtp_4_71/a_494_366# sky130_fd_sc_hs__dfrtp_4_55/a_37_78#
+ sky130_fd_sc_hs__and2_2_3/a_118_74# sky130_fd_sc_hs__dfrbp_1_37/a_1434_74# sky130_fd_sc_hs__nor2b_1_17/a_27_112#
+ sky130_fd_sc_hs__dfrtp_4_17/a_1350_392# sky130_fd_sc_hs__a22o_1_3/a_132_392# sky130_fd_sc_hs__nand2_1_49/a_117_74#
+ sky130_fd_sc_hs__fa_2_1/a_1202_368# sky130_fd_sc_hs__a222o_1_1/a_119_74# sky130_fd_sc_hs__dfxtp_4_5/a_437_503#
+ sky130_fd_sc_hs__conb_1_3/LO sky130_fd_sc_hs__nor2b_2_1/a_228_368# sky130_fd_sc_hs__dfrbp_1_45/a_832_118#
+ sky130_fd_sc_hs__dfrbp_1_33/a_2026_424# sky130_fd_sc_hs__nand2_1_93/a_117_74# sky130_fd_sc_hs__dfxtp_2_5/a_1019_424#
+ sky130_fd_sc_hs__dfrtn_1_19/a_817_508# sky130_fd_sc_hs__a22oi_1_17/a_71_368# sky130_fd_sc_hs__sdlclkp_1_1/a_116_424#
+ sky130_fd_sc_hs__nand2_1_9/a_117_74# sky130_fd_sc_hs__nor3_1_9/a_114_368# sky130_fd_sc_hs__dfrtp_4_47/a_2010_409#
+ sky130_fd_sc_hs__a21oi_1_103/a_117_74# sky130_fd_sc_hs__nor2_1_55/a_116_368# sky130_fd_sc_hs__a2bb2oi_1_1/a_117_392#
+ sky130_fd_sc_hs__nor2_1_53/Y sky130_fd_sc_hs__dfrtp_4_53/a_699_463# sky130_fd_sc_hs__dfstp_2_5/a_1057_118#
+ sky130_fd_sc_hs__o21a_1_43/a_320_74# sky130_fd_sc_hs__dfrtp_4_3/a_1678_395# sky130_fd_sc_hs__a22o_1_17/a_132_392#
+ sky130_fd_sc_hs__o22ai_1_3/a_27_74# sky130_fd_sc_hs__dfrtn_1_13/a_1598_93# sky130_fd_sc_hs__dfrtp_4_17/a_812_138#
+ sky130_fd_sc_hs__nor2b_1_27/Y sky130_fd_sc_hs__a21oi_1_43/a_29_368# sky130_fd_sc_hs__nor2_1_13/B
+ sky130_fd_sc_hs__nor4_1_1/Y sky130_fd_sc_hs__dfrtp_4_57/a_812_138# sky130_fd_sc_hs__dfxtp_2_11/a_695_459#
+ sky130_fd_sc_hs__dfrbp_1_3/a_1465_471# sky130_fd_sc_hs__dfrtn_1_35/a_856_304# sky130_fd_sc_hs__dfrtn_1_35/a_850_127#
+ sky130_fd_sc_hs__dfrbp_1_3/a_1434_74# sky130_fd_sc_hs__dfrtn_1_11/a_33_74# sky130_fd_sc_hs__fa_2_3/a_1205_79#
+ sky130_fd_sc_hs__dfrtp_4_5/a_1647_81# sky130_fd_sc_hs__dfrtn_1_15/a_507_368# sky130_fd_sc_hs__dfrtn_1_31/a_714_127#
+ sky130_fd_sc_hs__dfrtp_4_1/a_1827_81# sky130_fd_sc_hs__dfrtp_4_27/a_789_463# sky130_fd_sc_hs__dfrtn_1_47/a_1736_119#
+ sky130_fd_sc_hs__dfrtp_4_75/a_1827_81# sky130_fd_sc_hs__dfrtn_1_47/a_1266_119# sky130_fd_sc_hs__o211ai_1_9/a_31_74#
+ sky130_fd_sc_hs__nor2_1_5/a_116_368# sky130_fd_sc_hs__dfrtp_4_67/a_1350_392# sky130_fd_sc_hs__dfrbp_1_17/a_706_463#
+ sky130_fd_sc_hs__a22o_1_29/a_222_392# sky130_fd_sc_hs__a21oi_1_29/a_117_74# sky130_fd_sc_hs__fa_2_1/a_27_79#
+ sky130_fd_sc_hs__dfrbp_1_47/a_319_360# sky130_fd_sc_hs__dfstp_2_4/a_1489_118# sky130_fd_sc_hs__a211oi_4_1/a_77_368#
+ sky130_fd_sc_hs__dfrtp_4_21/a_494_366# sky130_fd_sc_hs__dfrtp_4_63/a_1678_395# sky130_fd_sc_hs__dfrtp_4_27/a_1627_493#
+ sky130_fd_sc_hs__dfxtp_2_9/a_1172_124# sky130_fd_sc_hs__dfrtn_1_37/a_300_74# sky130_fd_sc_hs__dfrtp_4_61/a_494_366#
+ sky130_fd_sc_hs__dfrtp_4_79/a_313_74# sky130_fd_sc_hs__nor2_2_3/A sky130_fd_sc_hs__a21oi_1_73/a_117_74#
+ sky130_fd_sc_hs__dfrbp_1_35/a_38_78# sky130_fd_sc_hs__dfrtn_1_1/a_856_304# sky130_fd_sc_hs__dfrtn_1_1/a_850_127#
+ sky130_fd_sc_hs__a22o_1_7/a_230_79# sky130_fd_sc_hs__nor2b_1_43/Y sky130_fd_sc_hs__dfrbp_1_41/a_1482_48#
+ sky130_fd_sc_hs__dfrtp_4_13/a_1678_395# sky130_fd_sc_hs__dfrtp_4_13/a_313_74# sky130_fd_sc_hs__dfrbp_1_45/a_125_78#
+ sky130_fd_sc_hs__dfrtp_4_5/a_890_138# sky130_fd_sc_hs__dfxtp_2_3/a_1019_424# sky130_fd_sc_hs__dfrbp_1_15/a_1465_471#
+ sky130_fd_sc_hs__dfrbp_1_3/Q_N sky130_fd_sc_hs__dfrtn_1_49/a_817_508# sky130_fd_sc_hs__a22o_1_17/a_230_79#
+ sky130_fd_sc_hs__or2_1_1/a_63_368# sky130_fd_sc_hs__nor2_1_45/a_116_368# sky130_fd_sc_hs__dfrtp_4_5/a_1350_392#
+ sky130_fd_sc_hs__o21a_1_31/a_83_244# sky130_fd_sc_hs__dfstp_2_4/a_1057_118# sky130_fd_sc_hs__dfrtn_1_37/a_33_74#
+ sky130_fd_sc_hs__dfrtp_4_83/a_699_463# sky130_fd_sc_hs__dfstp_2_4/a_612_74# sky130_fd_sc_hs__a22oi_1_23/a_159_74#
+ sky130_fd_sc_hs__dfrbp_1_45/a_841_401# sky130_fd_sc_hs__dfrtn_1_27/a_1550_119# sky130_fd_sc_hs__nor3_1_3/a_198_368#
+ sky130_fd_sc_hs__dfxtp_4_9/a_1141_508# sky130_fd_sc_hs__a22o_1_5/a_222_392# sky130_fd_sc_hs__dfrtn_1_41/a_1934_94#
+ sky130_fd_sc_hs__dfrtn_1_43/a_1598_93# sky130_fd_sc_hs__nand2_1_63/a_117_74# sky130_fd_sc_hs__a21oi_1_107/a_117_74#
+ sky130_fd_sc_hs__dfrtp_4_57/a_124_78# sky130_fd_sc_hs__dfrbp_1_1/a_1465_471# sky130_fd_sc_hs__dfrtn_1_25/a_856_304#
+ sky130_fd_sc_hs__o31ai_1_3/a_119_368# sky130_fd_sc_hs__dfxtp_2_7/a_431_508# sky130_fd_sc_hs__dfrtn_1_25/a_850_127#
+ sky130_fd_sc_hs__dfxtp_4_3/a_1226_296# sky130_fd_sc_hs__nand2_1_31/a_117_74# sky130_fd_sc_hs__o21a_1_47/a_320_74#
+ sky130_fd_sc_hs__fa_2_23/a_484_347# sky130_fd_sc_hs__a21oi_1_79/a_29_368# sky130_fd_sc_hs__dfrtp_4_25/a_1827_81#
+ sky130_fd_sc_hs__nand2_2_7/a_27_74# sky130_fd_sc_hs__o21a_1_13/a_320_74# sky130_fd_sc_hs__dfrtp_4_77/a_1627_493#
+ sky130_fd_sc_hs__dfrtn_1_21/a_714_127# sky130_fd_sc_hs__dfrbp_1_1/a_832_118# sky130_fd_sc_hs__dfrtp_4_65/a_1827_81#
+ sky130_fd_sc_hs__a21oi_1_47/a_29_368# sky130_fd_sc_hs__dfrbp_1_23/a_796_463# sky130_fd_sc_hs__dfstp_2_5/a_767_384#
+ sky130_fd_sc_hs__a22o_1_19/a_222_392# sky130_fd_sc_hs__dfstp_2_7/a_27_74# sky130_fd_sc_hs__dfstp_2_1/a_1489_118#
+ sky130_fd_sc_hs__a21oi_1_91/a_29_368# sky130_fd_sc_hs__dfrtp_4_25/a_1627_493# sky130_fd_sc_hs__dfxtp_2_7/a_1172_124#
+ sky130_fd_sc_hs__dfrtp_4_51/a_494_366# sky130_fd_sc_hs__fa_2_23/a_1202_368# sky130_fd_sc_hs__a222o_1_1/a_651_74#
+ sky130_fd_sc_hs__a22o_1_3/a_52_123# sky130_fd_sc_hs__dfrtp_4_15/a_1350_392# sky130_fd_sc_hs__fa_2_3/a_487_79#
+ sky130_fd_sc_hs__dfrbp_1_25/a_832_118# sky130_fd_sc_hs__o21a_1_69/a_376_387# sky130_fd_sc_hs__dfrbp_1_31/a_2026_424#
+ sky130_fd_sc_hs__nor2_2_3/B sky130_fd_sc_hs__dfrbp_1_43/a_910_118# sky130_fd_sc_hs__nor2_1_35/a_116_368#
+ sky130_fd_sc_hs__dfrtp_4_49/a_313_74# sky130_fd_sc_hs__dfrtn_1_25/a_120_74# sky130_fd_sc_hs__dfrtp_4_9/a_699_463#
+ sky130_fd_sc_hs__nor2_1_73/a_116_368# sky130_fd_sc_hs__dfstp_2_1/a_1057_118# sky130_fd_sc_hs__dfrtp_4_1/a_1678_395#
+ sky130_fd_sc_hs__dfrtn_1_17/D sky130_fd_sc_hs__dfrtp_4_63/a_37_78# sky130_fd_sc_hs__dfrtn_1_9/a_922_127#
+ sky130_fd_sc_hs__nor2b_1_49/a_278_368# sky130_fd_sc_hs__dfrtn_1_31/a_1934_94# sky130_fd_sc_hs__dfrtn_1_33/a_1598_93#
+ sky130_fd_sc_hs__dfrtp_4_61/a_313_74# sky130_fd_sc_hs__dfrtn_1_15/a_856_304# sky130_fd_sc_hs__dfrtn_1_15/a_850_127#
+ sky130_fd_sc_hs__dfxtp_4_2/a_1226_296# sky130_fd_sc_hs__o21a_1_39/X sky130_fd_sc_hs__fa_2_13/a_484_347#
+ sky130_fd_sc_hs__dfrtp_4_15/a_1827_81# sky130_fd_sc_hs__dfrtn_1_11/a_714_127# sky130_fd_sc_hs__nor2b_1_35/a_27_112#
+ sky130_fd_sc_hs__dfrtp_4_55/a_1827_81# sky130_fd_sc_hs__dfrbp_1_13/a_796_463# sky130_fd_sc_hs__dfrbp_1_39/a_498_360#
+ sky130_fd_sc_hs__dfrtp_4_85/a_789_463# sky130_fd_sc_hs__a22oi_1_21/a_339_74# sky130_fd_sc_hs__nand2_1_35/a_117_74#
+ sky130_fd_sc_hs__o22ai_1_11/a_27_74# sky130_fd_sc_hs__dfrtn_1_37/a_1547_508# sky130_fd_sc_hs__dfrbp_1_37/a_706_463#
+ sky130_fd_sc_hs__dfrtp_4_27/a_834_355# sky130_fd_sc_hs__dfrbp_1_27/a_319_360# sky130_fd_sc_hs__xnor2_1_13/a_293_74#
+ sky130_fd_sc_hs__dfstp_2_5/a_1596_118# sky130_fd_sc_hs__dfrtp_4_41/a_494_366# sky130_fd_sc_hs__dfrbp_1_11/Q_N
+ sky130_fd_sc_hs__dfrbp_1_1/a_841_401# sky130_fd_sc_hs__dfrbp_1_45/a_1434_74# sky130_fd_sc_hs__dfrbp_1_5/a_1624_74#
+ sky130_fd_sc_hs__dfrbp_1_29/a_38_78# sky130_fd_sc_hs__xnor2_1_5/a_112_119# sky130_fd_sc_hs__dfrbp_1_15/a_832_118#
+ sky130_fd_sc_hs__dfrtp_4_11/a_1678_395# sky130_fd_sc_hs__a21oi_1_95/a_29_368# sky130_fd_sc_hs__o21a_1_59/a_376_387#
+ sky130_fd_sc_hs__dfxtp_2_1/a_1019_424# sky130_fd_sc_hs__dfrbp_1_13/a_1465_471# sky130_fd_sc_hs__dfstp_2_1/a_398_74#
+ sky130_fd_sc_hs__fa_2_13/a_27_378# sky130_fd_sc_hs__fa_2_7/a_992_347# sky130_fd_sc_hs__o21a_1_69/X
+ sky130_fd_sc_hs__dfxtp_4_7/a_696_458# sky130_fd_sc_hs__a22o_1_7/a_52_123# sky130_fd_sc_hs__dfrtp_4_45/a_2010_409#
+ sky130_fd_sc_hs__dfrtp_4_89/a_37_78# sky130_fd_sc_hs__dfrtp_4_17/a_37_78# sky130_fd_sc_hs__nor2_1_25/a_116_368#
+ sky130_fd_sc_hs__o21a_1_5/a_376_387# sky130_fd_sc_hs__fa_2_7/a_487_79# sky130_fd_sc_hs__fa_2_17/SUM
+ sky130_fd_sc_hs__nor2b_1_7/a_278_368# sky130_fd_sc_hs__nor2_1_109/a_116_368# sky130_fd_sc_hs__a22o_1_17/a_52_123#
+ sky130_fd_sc_hs__maj3_1_1/a_406_384# sky130_fd_sc_hs__dfrbp_1_25/a_841_401# sky130_fd_sc_hs__dfrbp_1_3/a_706_463#
+ sky130_fd_sc_hs__dfxtp_4_7/a_1141_508# sky130_fd_sc_hs__dfrbp_1_29/a_1624_74# sky130_fd_sc_hs__fa_2_17/a_992_347#
+ sky130_fd_sc_hs__nor2b_1_39/a_278_368# sky130_fd_sc_hs__o21ai_1_7/a_27_74# sky130_fd_sc_hs__dfrtn_1_21/a_1934_94#
+ sky130_fd_sc_hs__dfrtn_1_23/a_1598_93# sky130_fd_sc_hs__dfrtp_4_27/a_812_138# sky130_fd_sc_hs__dfrbp_1_43/a_38_78#
+ sky130_fd_sc_hs__dfstp_2_7/a_716_456# sky130_fd_sc_hs__fa_2_13/a_701_79# sky130_fd_sc_hs__a21oi_1_15/a_117_74#
+ sky130_fd_sc_hs__dfrtp_4_1/a_313_74# sky130_fd_sc_hs__fa_2_9/a_683_347# sky130_fd_sc_hs__dfrtp_4_75/a_1627_493#
+ sky130_fd_sc_hs__o22ai_1_3/a_340_368# sky130_fd_sc_hs__dfrtp_4_49/a_1647_81# sky130_fd_sc_hs__dfrtn_1_45/a_1736_119#
+ sky130_fd_sc_hs__dfrtp_4_45/a_1827_81# sky130_fd_sc_hs__dfrtp_4_33/a_37_78# sky130_fd_sc_hs__dfrtn_1_23/a_300_74#
+ sky130_fd_sc_hs__dfrtp_4_89/a_1647_81# sky130_fd_sc_hs__nand4_1_3/a_259_74# sky130_fd_sc_hs__conb_1_3/HI
+ sky130_fd_sc_hs__dfrtn_1_45/a_1266_119# sky130_fd_sc_hs__dfrtp_4_65/a_313_74# sky130_fd_sc_hs__xor2_1_7/a_355_368#
+ sky130_fd_sc_hs__dfrtp_4_1/a_789_463# sky130_fd_sc_hs__dfrtp_4_65/a_1350_392# sky130_fd_sc_hs__nor3_1_13/a_114_368#
+ sky130_fd_sc_hs__sdlclkp_4_1/a_785_455# sky130_fd_sc_hs__dfrtn_1_3/a_120_74# sky130_fd_sc_hs__xnor2_1_13/a_112_119#
+ sky130_fd_sc_hs__dfrtp_4_75/a_789_463# sky130_fd_sc_hs__o21a_1_39/a_83_244# sky130_fd_sc_hs__dfrbp_1_17/a_319_360#
+ sky130_fd_sc_hs__dfxtp_2_1/a_644_504# sky130_fd_sc_hs__dfrtp_4_61/a_1678_395# sky130_fd_sc_hs__fa_2_19/a_683_347#
+ sky130_fd_sc_hs__dfstp_2_4/a_1596_118# sky130_fd_sc_hs__fa_2_23/a_1205_79# sky130_fd_sc_hs__dfrtp_4_31/a_494_366#
+ sky130_fd_sc_hs__fa_2_21/a_1202_368# sky130_fd_sc_hs__nor2b_1_39/a_27_112# sky130_fd_sc_hs__o21ai_1_9/a_162_368#
+ sky130_fd_sc_hs__o21a_1_11/X sky130_fd_sc_hs__a22oi_1_25/a_339_74# sky130_fd_sc_hs__nand2_1_39/a_117_74#
+ sky130_fd_sc_hs__dfsbp_2_1/a_398_74# sky130_fd_sc_hs__o21a_1_49/a_376_387# sky130_fd_sc_hs__dfxtp_2_9/a_1217_314#
+ sky130_fd_sc_hs__dfrtp_4_49/a_890_138# sky130_fd_sc_hs__dfrtp_4_29/a_1678_395# sky130_fd_sc_hs__dfrbp_1_47/a_2026_424#
+ sky130_fd_sc_hs__dfrtp_4_89/a_890_138# sky130_fd_sc_hs__nand2_1_83/a_117_74# sky130_fd_sc_hs__or2_1_1/a_152_368#
+ sky130_fd_sc_hs__dfrbp_1_23/a_910_118# sky130_fd_sc_hs__nor2_1_15/a_116_368# sky130_fd_sc_hs__dfrtp_4_3/a_1350_392#
+ sky130_fd_sc_hs__dfxtp_4_3/a_735_102# sky130_fd_sc_hs__dfrtp_4_43/a_124_78# sky130_fd_sc_hs__a21oi_1_99/a_29_368#
+ sky130_fd_sc_hs__nor2_1_93/a_116_368# sky130_fd_sc_hs__o21a_1_33/a_320_74# sky130_fd_sc_hs__dfrbp_1_15/a_841_401#
+ sky130_fd_sc_hs__dfrtn_1_25/a_1550_119# sky130_fd_sc_hs__dfrbp_1_19/a_1624_74# sky130_fd_sc_hs__o31ai_1_3/a_203_368#
+ sky130_fd_sc_hs__dfrtn_1_11/a_1934_94# sky130_fd_sc_hs__dfrtn_1_9/a_1736_119# sky130_fd_sc_hs__dfrbp_1_1/a_1434_74#
+ sky130_fd_sc_hs__dfrtn_1_9/a_1266_119# sky130_fd_sc_hs__dfrtp_4_73/a_1627_493# sky130_fd_sc_hs__dfrtp_4_35/a_1827_81#
+ sky130_fd_sc_hs__dfrtn_1_13/a_507_368# sky130_fd_sc_hs__dfrtp_4_79/a_1647_81# sky130_fd_sc_hs__dfrbp_1_39/a_1224_74#
+ sky130_fd_sc_hs__dfrtp_4_9/a_37_78# sky130_fd_sc_hs__dfrtp_4_25/a_789_463# sky130_fd_sc_hs__dfrtp_4_73/a_1827_81#
+ sky130_fd_sc_hs__dfrtp_4_63/a_1350_392# sky130_fd_sc_hs__dfrbp_1_33/a_796_463# sky130_fd_sc_hs__dfrtp_4_65/a_789_463#
+ sky130_fd_sc_hs__dfstp_2_5/a_2022_94# sky130_fd_sc_hs__inv_2_9/Y sky130_fd_sc_hs__dfrtn_1_35/a_1547_508#
+ sky130_fd_sc_hs__o22ai_1_3/a_142_368# sky130_fd_sc_hs__dfrtp_4_23/a_1627_493# sky130_fd_sc_hs__a21oi_1_19/a_117_74#
+ sky130_fd_sc_hs__dfxtp_2_5/a_1172_124# sky130_fd_sc_hs__dfstp_2_1/a_1596_118# sky130_fd_sc_hs__fa_2_13/a_1205_79#
+ sky130_fd_sc_hs__dfrtp_4_79/a_1678_395# sky130_fd_sc_hs__dfrtp_4_85/a_834_355# sky130_fd_sc_hs__xor2_1_1/a_194_125#
+ sky130_fd_sc_hs__dfrtp_4_13/a_1350_392# sky130_fd_sc_hs__dfrtp_4_69/a_313_74# sky130_fd_sc_hs__dfrbp_1_25/a_1434_74#
+ sky130_fd_sc_hs__a21oi_1_63/a_117_74# sky130_fd_sc_hs__o21a_1_39/a_376_387# sky130_fd_sc_hs__dfsbp_2_1/a_1258_341#
+ sky130_fd_sc_hs__dfxtp_2_7/a_1217_314# sky130_fd_sc_hs__dfrtn_1_15/a_33_74# sky130_fd_sc_hs__dfrbp_1_35/a_832_118#
+ sky130_fd_sc_hs__dfrtn_1_9/a_714_127# sky130_fd_sc_hs__dfrtp_4_79/a_890_138# sky130_fd_sc_hs__dfrbp_1_1/a_38_78#
+ sky130_fd_sc_hs__dfrtp_4_43/a_2010_409# sky130_fd_sc_hs__dfrbp_1_13/a_910_118# sky130_fd_sc_hs__dfrtn_1_47/a_817_508#
+ sky130_fd_sc_hs__fa_2_23/SUM sky130_fd_sc_hs__dfrbp_1_9/a_796_463# sky130_fd_sc_hs__dfrtp_4_43/a_699_463#
+ sky130_fd_sc_hs__fa_2_11/a_487_79# sky130_fd_sc_hs__o21a_1_21/a_83_244# sky130_fd_sc_hs__nor2_1_83/a_116_368#
+ sky130_fd_sc_hs__a222oi_1_1/a_697_74# sky130_fd_sc_hs__dfxtp_4_5/a_1141_508# sky130_fd_sc_hs__a22oi_1_13/a_159_74#
+ sky130_fd_sc_hs__nand2_1_87/a_117_74# sky130_fd_sc_hs__dfrbp_1_47/a_1624_74# sky130_fd_sc_hs__conb_1_3/a_21_290#
+ sky130_fd_sc_hs__dfrtn_1_41/a_1598_93# sky130_fd_sc_hs__nand2b_1_1/a_269_74# sky130_fd_sc_hs__a22oi_1_5/a_339_74#
+ sky130_fd_sc_hs__dfrtn_1_7/a_1736_119# sky130_fd_sc_hs__dfrtp_4_85/a_812_138# sky130_fd_sc_hs__nand2_1_21/a_117_74#
+ sky130_fd_sc_hs__dfrtn_1_7/a_1266_119# sky130_fd_sc_hs__xnor2_1_5/a_138_385# sky130_fd_sc_hs__dfrtn_1_43/a_1736_119#
+ sky130_fd_sc_hs__dfrtp_4_91/a_124_78# sky130_fd_sc_hs__dfxtp_2_5/a_695_459# sky130_fd_sc_hs__dfrtp_4_69/a_1647_81#
+ sky130_fd_sc_hs__dfrtn_1_43/a_1266_119# sky130_fd_sc_hs__dfrtp_4_15/a_789_463# sky130_fd_sc_hs__dfrtp_4_63/a_1827_81#
+ sky130_fd_sc_hs__dfrtp_4_27/a_37_78# sky130_fd_sc_hs__dfrtn_1_43/a_507_368# sky130_fd_sc_hs__dfrtp_4_55/a_789_463#
+ sky130_fd_sc_hs__dfstp_2_4/a_767_384# sky130_fd_sc_hs__inv_4_15/A sky130_fd_sc_hs__dfrtp_4_21/a_1627_493#
+ sky130_fd_sc_hs__dfxtp_2_3/a_1172_124# sky130_fd_sc_hs__dfrbp_1_45/a_706_463# sky130_fd_sc_hs__dfrbp_1_37/a_319_360#
+ sky130_fd_sc_hs__a21oi_1_82/a_29_368# sky130_fd_sc_hs__dfrtp_4_11/a_494_366# sky130_fd_sc_hs__dfrtn_1_39/a_33_74#
+ sky130_fd_sc_hs__dfrtp_4_1/a_834_355# sky130_fd_sc_hs__dfrtp_4_75/a_834_355# sky130_fd_sc_hs__nand4_1_1/a_181_74#
+ sky130_fd_sc_hs__dfrbp_1_15/a_1434_74# sky130_fd_sc_hs__o21a_1_29/a_376_387# sky130_fd_sc_hs__dfrbp_1_31/a_1482_48#
+ sky130_fd_sc_hs__dfrbp_1_11/a_1465_471# sky130_fd_sc_hs__dfrtp_4_27/a_1678_395#
+ sky130_fd_sc_hs__dfxtp_4_5/a_651_503# sky130_fd_sc_hs__maj3_1_3/a_595_136# sky130_fd_sc_hs__dfrbp_1_45/a_2026_424#
+ sky130_fd_sc_hs__dfrtp_4_69/a_890_138# sky130_fd_sc_hs__dfxtp_4_7/a_544_485# sky130_fd_sc_hs__dfrtn_1_47/a_120_74#
+ sky130_fd_sc_hs__dfrtp_4_1/a_1350_392# sky130_fd_sc_hs__a21oi_1_67/a_117_74# sky130_fd_sc_hs__dfrtn_1_15/a_120_74#
+ sky130_fd_sc_hs__dfstp_2_4/a_781_74# sky130_fd_sc_hs__a21oi_1_33/a_117_74# sky130_fd_sc_hs__dfrtp_4_33/a_699_463#
+ sky130_fd_sc_hs__xnor2_1_13/a_138_385# sky130_fd_sc_hs__dfxtp_2_1/a_538_429# sky130_fd_sc_hs__nand4_2_1/Y
+ sky130_fd_sc_hs__dfrtn_1_23/a_1550_119# sky130_fd_sc_hs__dfrbp_1_39/a_125_78# sky130_fd_sc_hs__dfrtn_1_41/a_300_74#
+ sky130_fd_sc_hs__fa_2_1/a_484_347# sky130_fd_sc_hs__nor2_1_119/a_116_368# sky130_fd_sc_hs__dfrbp_1_35/a_841_401#
+ sky130_fd_sc_hs__dfrtn_1_5/a_300_74# sky130_fd_sc_hs__dfrbp_1_3/a_319_360# sky130_fd_sc_hs__dfrtn_1_7/a_922_127#
+ sky130_fd_sc_hs__xnor2_1_3/a_376_368# sky130_fd_sc_hs__dfrbp_1_13/Q_N sky130_fd_sc_hs__o211ai_1_11/a_311_74#
+ sky130_fd_sc_hs__dfrtn_1_31/a_1598_93# sky130_fd_sc_hs__dfrtp_4_51/a_313_74# sky130_fd_sc_hs__dfrtn_1_13/a_856_304#
+ sky130_fd_sc_hs__dfrtp_4_1/a_812_138# sky130_fd_sc_hs__dfrtp_4_75/a_812_138# sky130_fd_sc_hs__o2bb2ai_1_1/a_490_368#
+ sky130_fd_sc_hs__dfrtn_1_13/a_850_127# sky130_fd_sc_hs__o21a_1_25/a_83_244# sky130_fd_sc_hs__fa_2_11/a_484_347#
+ sky130_fd_sc_hs__dfrtn_1_41/a_1736_119# sky130_fd_sc_hs__fa_2_7/a_1119_79# sky130_fd_sc_hs__a22oi_1_17/a_159_74#
+ sky130_fd_sc_hs__dfrbp_1_7/a_1482_48# sky130_fd_sc_hs__dfrtp_4_59/a_1647_81# sky130_fd_sc_hs__dfrtn_1_41/a_1266_119#
+ sky130_fd_sc_hs__dfrtp_4_53/a_1827_81# sky130_fd_sc_hs__a22o_1_21/a_230_79# sky130_fd_sc_hs__dfrtn_1_33/a_507_368#
+ sky130_fd_sc_hs__dfrtn_1_5/a_817_508# sky130_fd_sc_hs__dfrtp_4_45/a_789_463# sky130_fd_sc_hs__nor4_1_3/a_342_368#
+ sky130_fd_sc_hs__nand2b_1_5/a_269_74# sky130_fd_sc_hs__dfrtn_1_33/a_1547_508# sky130_fd_sc_hs__a222oi_1_1/a_119_74#
+ sky130_fd_sc_hs__a22oi_1_11/a_339_74# sky130_fd_sc_hs__nand2_1_25/a_117_74# sky130_fd_sc_hs__dfrtp_4_25/a_834_355#
+ sky130_fd_sc_hs__dfrtp_4_17/a_124_78# sky130_fd_sc_hs__fa_2_17/a_1119_79# sky130_fd_sc_hs__dfrtp_4_77/a_1678_395#
+ sky130_fd_sc_hs__dfrtp_4_65/a_834_355# sky130_fd_sc_hs__dfrtn_1_9/a_1934_94# sky130_fd_sc_hs__dfrtp_4_11/a_1350_392#
+ sky130_fd_sc_hs__o21a_1_19/a_376_387# sky130_fd_sc_hs__fa_2_11/a_27_79# sky130_fd_sc_hs__dfrbp_1_21/a_1482_48#
+ sky130_fd_sc_hs__nand2_1_15/Y sky130_fd_sc_hs__dfrtp_4_25/a_1678_395# sky130_fd_sc_hs__a21oi_1_85/a_29_368#
+ sky130_fd_sc_hs__dfrtp_4_59/a_890_138# sky130_fd_sc_hs__xnor2_1_11/a_376_368# sky130_fd_sc_hs__nand4_1_5/a_181_74#
+ sky130_fd_sc_hs__dfrtp_4_41/a_2010_409# sky130_fd_sc_hs__a22oi_1_3/a_71_368# sky130_fd_sc_hs__dfrbp_1_29/a_1465_471#
+ sky130_fd_sc_hs__a21oi_1_51/a_29_368# sky130_fd_sc_hs__fa_2_5/a_336_347# sky130_fd_sc_hs__dfrtn_1_27/a_817_508#
+ sky130_fd_sc_hs__a211oi_4_1/a_92_74# sky130_fd_sc_hs__dfrbp_1_33/a_910_118# sky130_fd_sc_hs__sdlclkp_1_1/a_288_48#
+ sky130_fd_sc_hs__a31oi_2_1/a_27_368# sky130_fd_sc_hs__dfrtp_4_23/a_699_463# sky130_fd_sc_hs__nor2_1_63/a_116_368#
+ sky130_fd_sc_hs__dfrbp_1_5/a_498_360# sky130_fd_sc_hs__dfrtn_1_21/a_1550_119# sky130_fd_sc_hs__dfrtp_4_11/a_37_78#
+ sky130_fd_sc_hs__a21oi_1_1/a_29_368# sky130_fd_sc_hs__a22o_1_25/a_132_392# sky130_fd_sc_hs__dfrbp_1_1/a_706_463#
+ sky130_fd_sc_hs__dfrbp_1_27/a_1624_74# sky130_fd_sc_hs__dfrtn_1_21/a_1598_93# sky130_fd_sc_hs__dfrtp_4_25/a_812_138#
+ sky130_fd_sc_hs__dfrtp_4_65/a_812_138# sky130_fd_sc_hs__a21oi_1_37/a_117_74# sky130_fd_sc_hs__dfrtn_1_43/a_856_304#
+ sky130_fd_sc_hs__dfrtp_4_71/a_1627_493# sky130_fd_sc_hs__dfrtn_1_43/a_850_127# sky130_fd_sc_hs__o21ai_1_11/a_27_74#
+ sky130_fd_sc_hs__dfrtn_1_9/a_300_74# sky130_fd_sc_hs__a21oi_1_83/a_117_74# sky130_fd_sc_hs__dfrtn_1_23/a_507_368#
+ sky130_fd_sc_hs__dfrtp_4_61/a_1350_392# sky130_fd_sc_hs__dfrtp_4_35/a_789_463# sky130_fd_sc_hs__dfrtp_4_55/a_313_74#
+ sky130_fd_sc_hs__dfrbp_1_29/a_498_360# sky130_fd_sc_hs__dfrtp_4_83/a_1827_81# sky130_fd_sc_hs__dfrtn_1_31/a_1547_508#
+ sky130_fd_sc_hs__dfrbp_1_41/a_796_463# sky130_fd_sc_hs__dfrtp_4_73/a_789_463# sky130_fd_sc_hs__o21a_1_29/a_83_244#
+ sky130_fd_sc_hs__fa_2_19/a_487_79# sky130_fd_sc_hs__dfrbp_1_9/a_910_118# sky130_fd_sc_hs__dfrtp_4_21/a_313_74#
+ sky130_fd_sc_hs__dfxtp_2_1/a_1172_124# sky130_fd_sc_hs__dfrbp_1_25/a_706_463# sky130_fd_sc_hs__a222o_1_1/a_337_390#
+ sky130_fd_sc_hs__dfrtp_4_15/a_834_355# sky130_fd_sc_hs__dfrtp_4_39/a_1627_493# sky130_fd_sc_hs__dfrtp_4_55/a_834_355#
+ sky130_fd_sc_hs__nor4_1_3/a_144_368# sky130_fd_sc_hs__dfrtp_4_5/a_494_366# sky130_fd_sc_hs__o21a_1_73/a_83_244#
+ sky130_fd_sc_hs__dfrtp_4_91/a_2010_409# sky130_fd_sc_hs__maj3_1_3/a_223_120# sky130_fd_sc_hs__nand2b_1_9/a_269_74#
+ sky130_fd_sc_hs__dfrtp_4_29/a_1350_392# sky130_fd_sc_hs__dfrbp_1_35/a_1434_74# sky130_fd_sc_hs__a211oi_1_1/a_71_368#
+ sky130_fd_sc_hs__a22o_1_1/a_132_392# sky130_fd_sc_hs__dfxtp_2_5/a_1217_314# sky130_fd_sc_hs__a22oi_1_15/a_339_74#
+ sky130_fd_sc_hs__nand2_1_29/a_117_74# sky130_fd_sc_hs__dfrbp_1_11/a_1482_48# sky130_fd_sc_hs__dfrbp_1_43/a_2026_424#
+ sky130_fd_sc_hs__dfrbp_1_43/a_832_118# sky130_fd_sc_hs__nor2b_1_41/a_27_112# sky130_fd_sc_hs__dfrbp_1_27/a_1465_471#
+ sky130_fd_sc_hs__nand2_1_73/a_117_74# sky130_fd_sc_hs__a21oi_1_117/a_117_74# sky130_fd_sc_hs__dfrtn_1_17/a_817_508#
+ sky130_fd_sc_hs__dfrtp_4_59/a_2010_409# sky130_fd_sc_hs__nor3_1_7/a_114_368# sky130_fd_sc_hs__dfxtp_4_2/a_735_102#
+ sky130_fd_sc_hs__dfstp_2_1/a_225_74# sky130_fd_sc_hs__nand2_4_13/a_27_74# sky130_fd_sc_hs__dfrtp_4_13/a_699_463#
+ sky130_fd_sc_hs__dfrtp_4_33/a_124_78# sky130_fd_sc_hs__nor2_1_53/a_116_368# sky130_fd_sc_hs__o211ai_1_3/a_311_74#
+ sky130_fd_sc_hs__a21oi_1_89/a_29_368# sky130_fd_sc_hs__dfxtp_4_3/a_1141_508# sky130_fd_sc_hs__dfrtn_1_49/a_33_74#
+ sky130_fd_sc_hs__o21a_1_23/a_320_74# sky130_fd_sc_hs__a22o_1_15/a_132_392# sky130_fd_sc_hs__dfrtp_4_91/a_699_463#
+ sky130_fd_sc_hs__dfxtp_2_11/a_431_508# sky130_fd_sc_hs__dfrbp_1_17/a_1624_74# sky130_fd_sc_hs__dfrtn_1_39/a_1550_119#
+ sky130_fd_sc_hs__a22oi_1_7/a_71_368# sky130_fd_sc_hs__nor2b_1_29/a_278_368# sky130_fd_sc_hs__dfrtn_1_11/a_1598_93#
+ sky130_fd_sc_hs__dfrtp_4_15/a_812_138# sky130_fd_sc_hs__nand2_1_1/a_117_74# sky130_fd_sc_hs__a21oi_1_23/a_29_368#
+ sky130_fd_sc_hs__dfrtn_1_5/a_1736_119# sky130_fd_sc_hs__dfrtp_4_55/a_812_138# sky130_fd_sc_hs__dfrtn_1_33/a_856_304#
+ sky130_fd_sc_hs__maj3_1_3/a_84_74# sky130_fd_sc_hs__dfrtn_1_5/a_1266_119# sky130_fd_sc_hs__nor4_1_3/a_228_368#
+ sky130_fd_sc_hs__dfrtn_1_33/a_850_127# sky130_fd_sc_hs__dfrtp_4_51/a_37_78# sky130_fd_sc_hs__dfrtp_4_39/a_1647_81#
+ sky130_fd_sc_hs__xor2_1_1/a_455_87# sky130_fd_sc_hs__a21oi_1_5/a_29_368# sky130_fd_sc_hs__dfrtp_4_89/a_1627_493#
+ sky130_fd_sc_hs__fa_2_1/a_1205_79#
Xsky130_fd_sc_hs__xnor2_1_7 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__xnor2_1_7/A sky130_fd_sc_hs__xnor2_1_7/Y
+ sky130_fd_sc_hs__xnor2_1_7/B sky130_fd_sc_hs__xnor2_1_7/a_376_368# sky130_fd_sc_hs__xnor2_1_7/a_112_119#
+ sky130_fd_sc_hs__xnor2_1_7/a_138_385# sky130_fd_sc_hs__xnor2_1_7/a_293_74# sky130_fd_sc_hs__xnor2_1
Xsky130_fd_sc_hs__nor2b_1_32 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__dfxtp_4_7/Q sky130_fd_sc_hs__nor2b_1_33/Y
+ sky130_fd_sc_hs__dfxtp_4_2/Q sky130_fd_sc_hs__nor2b_1_33/a_278_368# sky130_fd_sc_hs__nor2b_1_33/a_27_112#
+ sky130_fd_sc_hs__nor2b_1
Xsky130_fd_sc_hs__nor2b_1_21 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__fa_2_23/SUM sky130_fd_sc_hs__nor2b_1_21/Y
+ sky130_fd_sc_hs__or2_1_1/A sky130_fd_sc_hs__nor2b_1_21/a_278_368# sky130_fd_sc_hs__nor2b_1_21/a_27_112#
+ sky130_fd_sc_hs__nor2b_1
Xsky130_fd_sc_hs__nor2b_1_10 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__fa_2_9/SUM sky130_fd_sc_hs__nor2b_1_11/Y
+ sky130_fd_sc_hs__or2_1_1/A sky130_fd_sc_hs__nor2b_1_11/a_278_368# sky130_fd_sc_hs__nor2b_1_11/a_27_112#
+ sky130_fd_sc_hs__nor2b_1
Xsky130_fd_sc_hs__nor2b_1_43 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nor2_1_101/Y sky130_fd_sc_hs__nor2b_1_43/Y
+ sky130_fd_sc_hs__inv_4_87/A sky130_fd_sc_hs__nor2b_1_43/a_278_368# sky130_fd_sc_hs__nor2b_1_43/a_27_112#
+ sky130_fd_sc_hs__nor2b_1
Xsky130_fd_sc_hs__inv_4_102 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nor3_1_11/B sky130_fd_sc_hs__inv_4_103/A
+ sky130_fd_sc_hs__inv_4
Xsky130_fd_sc_hs__inv_4_113 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_113/Y sky130_fd_sc_hs__inv_4_113/A
+ sky130_fd_sc_hs__inv_4
Xsky130_fd_sc_hs__inv_4_124 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_125/Y sky130_fd_sc_hs__inv_4_125/A
+ sky130_fd_sc_hs__inv_4
Xsky130_fd_sc_hs__inv_4_135 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_135/Y sky130_fd_sc_hs__inv_4_135/A
+ sky130_fd_sc_hs__inv_4
Xsky130_fd_sc_hs__o22ai_1_2 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_53/Y sky130_fd_sc_hs__inv_4_51/A
+ sky130_fd_sc_hs__o22ai_1_3/Y sky130_fd_sc_hs__inv_4_39/Y sky130_fd_sc_hs__dfrbp_1_1/Q
+ sky130_fd_sc_hs__o22ai_1_3/a_340_368# sky130_fd_sc_hs__o22ai_1_3/a_142_368# sky130_fd_sc_hs__o22ai_1_3/a_27_74#
+ sky130_fd_sc_hs__o22ai_1
Xsky130_fd_sc_hs__nand2_4_13 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_4_13/Y aux_osc_en
+ sky130_fd_sc_hs__nand2_4_7/Y sky130_fd_sc_hs__nand2_4_13/a_27_74# sky130_fd_sc_hs__nand2_4
Xsky130_fd_sc_hs__and2_2_0 DVSS DVDD DVDD DVSS fine_control_avg_window_select[3] fine_control_avg_window_select[4]
+ sky130_fd_sc_hs__and2_2_1/X sky130_fd_sc_hs__and2_2_1/a_31_74# sky130_fd_sc_hs__and2_2_1/a_118_74#
+ sky130_fd_sc_hs__and2_2
Xsky130_fd_sc_hs__inv_4_8 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_9/Y sky130_fd_sc_hs__inv_4_9/A
+ sky130_fd_sc_hs__inv_4
Xsky130_fd_sc_hs__a22o_1_14 DVSS DVDD DVDD DVSS osc_fine_con_final[0] manual_control_osc[0]
+ sky130_fd_sc_hs__inv_4_43/Y sky130_fd_sc_hs__fa_2_9/A fftl_en sky130_fd_sc_hs__a22o_1_15/a_222_392#
+ sky130_fd_sc_hs__a22o_1_15/a_230_79# sky130_fd_sc_hs__a22o_1_15/a_52_123# sky130_fd_sc_hs__a22o_1_15/a_132_392#
+ sky130_fd_sc_hs__a22o_1
Xsky130_fd_sc_hs__a22o_1_25 DVSS DVDD DVDD DVSS osc_fine_con_final[10] manual_control_osc[10]
+ sky130_fd_sc_hs__inv_4_43/Y sky130_fd_sc_hs__fa_2_23/B fftl_en sky130_fd_sc_hs__a22o_1_25/a_222_392#
+ sky130_fd_sc_hs__a22o_1_25/a_230_79# sky130_fd_sc_hs__a22o_1_25/a_52_123# sky130_fd_sc_hs__a22o_1_25/a_132_392#
+ sky130_fd_sc_hs__a22o_1
Xsky130_fd_sc_hs__o21ai_1_1 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__o21ai_1_1/Y sky130_fd_sc_hs__o21ai_1_1/B1
+ sky130_fd_sc_hs__a32oi_1_1/Y fine_control_avg_window_select[0] sky130_fd_sc_hs__o21ai_1_1/a_162_368#
+ sky130_fd_sc_hs__o21ai_1_1/a_27_74# sky130_fd_sc_hs__o21ai_1
Xsky130_fd_sc_hs__nand2_1_14 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_21/Y sky130_fd_sc_hs__nand2_1_15/Y
+ fine_control_avg_window_select[2] sky130_fd_sc_hs__nand2_1_15/a_117_74# sky130_fd_sc_hs__nand2_1
Xsky130_fd_sc_hs__nand2_1_58 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_55/Y sky130_fd_sc_hs__nand2_1_59/Y
+ sky130_fd_sc_hs__nor2_1_59/A sky130_fd_sc_hs__nand2_1_59/a_117_74# sky130_fd_sc_hs__nand2_1
Xsky130_fd_sc_hs__nand2_1_47 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_1_47/B sky130_fd_sc_hs__nor2_1_75/B
+ sky130_fd_sc_hs__nor2b_1_33/Y sky130_fd_sc_hs__nand2_1_47/a_117_74# sky130_fd_sc_hs__nand2_1
Xsky130_fd_sc_hs__nand2_1_36 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nor2_1_29/Y sky130_fd_sc_hs__nor2_1_27/B
+ sky130_fd_sc_hs__inv_4_39/A sky130_fd_sc_hs__nand2_1_37/a_117_74# sky130_fd_sc_hs__nand2_1
Xsky130_fd_sc_hs__nand2_1_25 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nor2_1_13/Y sky130_fd_sc_hs__nor2_1_25/B
+ sky130_fd_sc_hs__o21a_1_21/A1 sky130_fd_sc_hs__nand2_1_25/a_117_74# sky130_fd_sc_hs__nand2_1
Xsky130_fd_sc_hs__nand2_1_69 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nor2_1_47/Y sky130_fd_sc_hs__o21a_1_57/B1
+ sky130_fd_sc_hs__inv_4_93/A sky130_fd_sc_hs__nand2_1_69/a_117_74# sky130_fd_sc_hs__nand2_1
Xsky130_fd_sc_hs__inv_2_5 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_2_5/A sky130_fd_sc_hs__inv_2_5/Y
+ sky130_fd_sc_hs__inv_2
Xsky130_fd_sc_hs__dfxtp_4_4 DVSS DVDD DVDD DVSS out_star sky130_fd_sc_hs__dfxtp_4_5/D
+ clk_out sky130_fd_sc_hs__dfxtp_4_5/a_1226_296# sky130_fd_sc_hs__dfxtp_4_5/a_735_102#
+ sky130_fd_sc_hs__dfxtp_4_5/a_1141_508# sky130_fd_sc_hs__dfxtp_4_5/a_206_368# sky130_fd_sc_hs__dfxtp_4_5/a_437_503#
+ sky130_fd_sc_hs__dfxtp_4_5/a_27_74# sky130_fd_sc_hs__dfxtp_4_5/a_651_503# sky130_fd_sc_hs__dfxtp_4_5/a_696_458#
+ sky130_fd_sc_hs__dfxtp_4_5/a_544_485# sky130_fd_sc_hs__dfxtp_4_5/a_1178_124# sky130_fd_sc_hs__dfxtp_4_5/a_1034_424#
+ sky130_fd_sc_hs__dfxtp_4
Xsky130_fd_sc_hs__nand2_4_9 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_4_9/Y aux_osc_en
+ sky130_fd_sc_hs__nand2_4_9/A sky130_fd_sc_hs__nand2_4_9/a_27_74# sky130_fd_sc_hs__nand2_4
Xsky130_fd_sc_hs__dfxtp_2_1 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__xnor2_1_3/A sky130_fd_sc_hs__dfxtp_4_9/CLK
+ sky130_fd_sc_hs__inv_2_1/Y sky130_fd_sc_hs__dfxtp_2_1/a_431_508# sky130_fd_sc_hs__dfxtp_2_1/a_1125_508#
+ sky130_fd_sc_hs__dfxtp_2_1/a_206_368# sky130_fd_sc_hs__dfxtp_2_1/a_27_74# sky130_fd_sc_hs__dfxtp_2_1/a_708_101#
+ sky130_fd_sc_hs__dfxtp_2_1/a_1019_424# sky130_fd_sc_hs__dfxtp_2_1/a_1172_124# sky130_fd_sc_hs__dfxtp_2_1/a_644_504#
+ sky130_fd_sc_hs__dfxtp_2_1/a_1217_314# sky130_fd_sc_hs__dfxtp_2_1/a_538_429# sky130_fd_sc_hs__dfxtp_2_1/a_695_459#
+ sky130_fd_sc_hs__dfxtp_2
Xsky130_fd_sc_hs__a21oi_1_103 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_123/Y sky130_fd_sc_hs__nand2_1_91/B
+ div_ratio_half[0] sky130_fd_sc_hs__inv_2_5/A sky130_fd_sc_hs__a21oi_1_103/a_117_74#
+ sky130_fd_sc_hs__a21oi_1_103/a_29_368# sky130_fd_sc_hs__a21oi_1
Xsky130_fd_sc_hs__a21oi_1_114 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__o21a_1_59/A2 sky130_fd_sc_hs__dfrtn_1_41/D
+ sky130_fd_sc_hs__o21a_1_71/B1 sky130_fd_sc_hs__inv_4_129/Y sky130_fd_sc_hs__a21oi_1_115/a_117_74#
+ sky130_fd_sc_hs__a21oi_1_115/a_29_368# sky130_fd_sc_hs__a21oi_1
Xsky130_fd_sc_hs__maj3_1_1 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__maj3_1_1/A sky130_fd_sc_hs__maj3_1_1/B
+ sky130_fd_sc_hs__maj3_1_1/X sky130_fd_sc_hs__maj3_1_1/C sky130_fd_sc_hs__maj3_1_1/a_598_384#
+ sky130_fd_sc_hs__maj3_1_1/a_226_384# sky130_fd_sc_hs__maj3_1_1/a_84_74# sky130_fd_sc_hs__maj3_1_1/a_403_136#
+ sky130_fd_sc_hs__maj3_1_1/a_406_384# sky130_fd_sc_hs__maj3_1_1/a_595_136# sky130_fd_sc_hs__maj3_1_1/a_223_120#
+ sky130_fd_sc_hs__maj3_1
Xsky130_fd_sc_hs__nand2_2_6 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_2_7/Y sky130_fd_sc_hs__nand2_2_7/B
+ sky130_fd_sc_hs__inv_2_9/A sky130_fd_sc_hs__nand2_2_7/a_27_74# sky130_fd_sc_hs__nand2_2
Xsky130_fd_sc_hs__nor2_2_2 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nor2_2_3/B sky130_fd_sc_hs__nor2_2_3/Y
+ sky130_fd_sc_hs__nor2_2_3/A sky130_fd_sc_hs__nor2_2_3/a_35_368# sky130_fd_sc_hs__nor2_2
Xsky130_fd_sc_hs__nor2_1_22 DVSS DVDD DVDD DVSS fine_control_avg_window_select[2]
+ sky130_fd_sc_hs__nor2_1_23/Y fine_control_avg_window_select[1] sky130_fd_sc_hs__nor2_1_23/a_116_368#
+ sky130_fd_sc_hs__nor2_1
Xsky130_fd_sc_hs__nor2_1_11 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__o21a_1_5/B1 sky130_fd_sc_hs__nor2_1_11/Y
+ sky130_fd_sc_hs__inv_4_13/Y sky130_fd_sc_hs__nor2_1_11/a_116_368# sky130_fd_sc_hs__nor2_1
Xsky130_fd_sc_hs__nor2_1_55 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_67/Y sky130_fd_sc_hs__nor4_1_1/B
+ sky130_fd_sc_hs__inv_4_63/A sky130_fd_sc_hs__nor2_1_55/a_116_368# sky130_fd_sc_hs__nor2_1
Xsky130_fd_sc_hs__nor2_1_44 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nor2_1_45/B sky130_fd_sc_hs__nor2_1_45/Y
+ sky130_fd_sc_hs__inv_4_63/Y sky130_fd_sc_hs__nor2_1_45/a_116_368# sky130_fd_sc_hs__nor2_1
Xsky130_fd_sc_hs__nor2_1_33 DVSS DVDD DVDD DVSS fine_control_avg_window_select[4]
+ sky130_fd_sc_hs__nor2_1_33/Y fine_control_avg_window_select[3] sky130_fd_sc_hs__nor2_1_33/a_116_368#
+ sky130_fd_sc_hs__nor2_1
Xsky130_fd_sc_hs__nor2_1_99 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nor2_1_99/B sky130_fd_sc_hs__nor2_1_99/Y
+ sky130_fd_sc_hs__nor2_1_99/A sky130_fd_sc_hs__nor2_1_99/a_116_368# sky130_fd_sc_hs__nor2_1
Xsky130_fd_sc_hs__nor2_1_88 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_87/A sky130_fd_sc_hs__nor2_1_89/Y
+ sky130_fd_sc_hs__nor2_1_89/A sky130_fd_sc_hs__nor2_1_89/a_116_368# sky130_fd_sc_hs__nor2_1
Xsky130_fd_sc_hs__nor2_1_77 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_87/A sky130_fd_sc_hs__nor2_1_77/Y
+ sky130_fd_sc_hs__or3b_2_1/X sky130_fd_sc_hs__nor2_1_77/a_116_368# sky130_fd_sc_hs__nor2_1
Xsky130_fd_sc_hs__nor2_1_66 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_65/Y sky130_fd_sc_hs__nor3_1_1/C
+ sky130_fd_sc_hs__inv_4_89/A sky130_fd_sc_hs__nor2_1_67/a_116_368# sky130_fd_sc_hs__nor2_1
Xsky130_fd_sc_hs__xnor2_1_8 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__xnor2_1_9/A sky130_fd_sc_hs__xnor2_1_9/Y
+ sky130_fd_sc_hs__xnor2_1_9/B sky130_fd_sc_hs__xnor2_1_9/a_376_368# sky130_fd_sc_hs__xnor2_1_9/a_112_119#
+ sky130_fd_sc_hs__xnor2_1_9/a_138_385# sky130_fd_sc_hs__xnor2_1_9/a_293_74# sky130_fd_sc_hs__xnor2_1
Xsky130_fd_sc_hs__nor2b_1_22 DVSS DVDD DVDD DVSS fine_control_avg_window_select[4]
+ sky130_fd_sc_hs__nor2b_1_23/Y fine_control_avg_window_select[3] sky130_fd_sc_hs__nor2b_1_23/a_278_368#
+ sky130_fd_sc_hs__nor2b_1_23/a_27_112# sky130_fd_sc_hs__nor2b_1
Xsky130_fd_sc_hs__nor2b_1_11 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__fa_2_9/SUM sky130_fd_sc_hs__nor2b_1_11/Y
+ sky130_fd_sc_hs__or2_1_1/A sky130_fd_sc_hs__nor2b_1_11/a_278_368# sky130_fd_sc_hs__nor2b_1_11/a_27_112#
+ sky130_fd_sc_hs__nor2b_1
Xsky130_fd_sc_hs__nor2b_1_44 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__o21a_1_63/A1 sky130_fd_sc_hs__nor3_1_13/C
+ sky130_fd_sc_hs__o21a_1_59/A1 sky130_fd_sc_hs__nor2b_1_45/a_278_368# sky130_fd_sc_hs__nor2b_1_45/a_27_112#
+ sky130_fd_sc_hs__nor2b_1
Xsky130_fd_sc_hs__nor2b_1_33 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__dfxtp_4_7/Q sky130_fd_sc_hs__nor2b_1_33/Y
+ sky130_fd_sc_hs__dfxtp_4_2/Q sky130_fd_sc_hs__nor2b_1_33/a_278_368# sky130_fd_sc_hs__nor2b_1_33/a_27_112#
+ sky130_fd_sc_hs__nor2b_1
Xsky130_fd_sc_hs__inv_4_103 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nor3_1_11/B sky130_fd_sc_hs__inv_4_103/A
+ sky130_fd_sc_hs__inv_4
Xsky130_fd_sc_hs__inv_4_114 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_115/Y sky130_fd_sc_hs__nor3_1_15/A
+ sky130_fd_sc_hs__inv_4
Xsky130_fd_sc_hs__inv_4_125 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_125/Y sky130_fd_sc_hs__inv_4_125/A
+ sky130_fd_sc_hs__inv_4
Xsky130_fd_sc_hs__inv_4_136 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_137/Y sky130_fd_sc_hs__inv_4_137/A
+ sky130_fd_sc_hs__inv_4
Xsky130_fd_sc_hs__o22ai_1_3 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_53/Y sky130_fd_sc_hs__inv_4_51/A
+ sky130_fd_sc_hs__o22ai_1_3/Y sky130_fd_sc_hs__inv_4_39/Y sky130_fd_sc_hs__dfrbp_1_1/Q
+ sky130_fd_sc_hs__o22ai_1_3/a_340_368# sky130_fd_sc_hs__o22ai_1_3/a_142_368# sky130_fd_sc_hs__o22ai_1_3/a_27_74#
+ sky130_fd_sc_hs__o22ai_1
Xsky130_fd_sc_hs__nand2_4_14 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__o21ai_2_1/B1 div_ratio_half[4]
+ sky130_fd_sc_hs__inv_4_103/A sky130_fd_sc_hs__nand2_4_15/a_27_74# sky130_fd_sc_hs__nand2_4
Xsky130_fd_sc_hs__and2_2_1 DVSS DVDD DVDD DVSS fine_control_avg_window_select[3] fine_control_avg_window_select[4]
+ sky130_fd_sc_hs__and2_2_1/X sky130_fd_sc_hs__and2_2_1/a_31_74# sky130_fd_sc_hs__and2_2_1/a_118_74#
+ sky130_fd_sc_hs__and2_2
Xsky130_fd_sc_hs__inv_4_90 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__or3b_2_1/B sky130_fd_sc_hs__inv_4_91/A
+ sky130_fd_sc_hs__inv_4
Xsky130_fd_sc_hs__inv_4_9 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_9/Y sky130_fd_sc_hs__inv_4_9/A
+ sky130_fd_sc_hs__inv_4
Xsky130_fd_sc_hs__dfxtp_2_10 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__xnor2_1_7/A sky130_fd_sc_hs__dfxtp_4_9/CLK
+ sky130_fd_sc_hs__nor2_1_91/Y sky130_fd_sc_hs__dfxtp_2_11/a_431_508# sky130_fd_sc_hs__dfxtp_2_11/a_1125_508#
+ sky130_fd_sc_hs__dfxtp_2_11/a_206_368# sky130_fd_sc_hs__dfxtp_2_11/a_27_74# sky130_fd_sc_hs__dfxtp_2_11/a_708_101#
+ sky130_fd_sc_hs__dfxtp_2_11/a_1019_424# sky130_fd_sc_hs__dfxtp_2_11/a_1172_124#
+ sky130_fd_sc_hs__dfxtp_2_11/a_644_504# sky130_fd_sc_hs__dfxtp_2_11/a_1217_314# sky130_fd_sc_hs__dfxtp_2_11/a_538_429#
+ sky130_fd_sc_hs__dfxtp_2_11/a_695_459# sky130_fd_sc_hs__dfxtp_2
Xsky130_fd_sc_hs__a22o_1_26 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__a22o_1_27/X sky130_fd_sc_hs__dfrbp_1_1/Q
+ sky130_fd_sc_hs__inv_4_39/Y sky130_fd_sc_hs__inv_4_61/A sky130_fd_sc_hs__inv_4_37/Y
+ sky130_fd_sc_hs__a22o_1_27/a_222_392# sky130_fd_sc_hs__a22o_1_27/a_230_79# sky130_fd_sc_hs__a22o_1_27/a_52_123#
+ sky130_fd_sc_hs__a22o_1_27/a_132_392# sky130_fd_sc_hs__a22o_1
Xsky130_fd_sc_hs__o21ai_1_2 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__o21ai_1_3/Y sky130_fd_sc_hs__o21ai_1_3/B1
+ sky130_fd_sc_hs__nor2_1_33/Y sky130_fd_sc_hs__and2_2_1/X sky130_fd_sc_hs__o21ai_1_3/a_162_368#
+ sky130_fd_sc_hs__o21ai_1_3/a_27_74# sky130_fd_sc_hs__o21ai_1
Xsky130_fd_sc_hs__a22o_1_15 DVSS DVDD DVDD DVSS osc_fine_con_final[0] manual_control_osc[0]
+ sky130_fd_sc_hs__inv_4_43/Y sky130_fd_sc_hs__fa_2_9/A fftl_en sky130_fd_sc_hs__a22o_1_15/a_222_392#
+ sky130_fd_sc_hs__a22o_1_15/a_230_79# sky130_fd_sc_hs__a22o_1_15/a_52_123# sky130_fd_sc_hs__a22o_1_15/a_132_392#
+ sky130_fd_sc_hs__a22o_1
Xsky130_fd_sc_hs__nand2_1_15 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_21/Y sky130_fd_sc_hs__nand2_1_15/Y
+ fine_control_avg_window_select[2] sky130_fd_sc_hs__nand2_1_15/a_117_74# sky130_fd_sc_hs__nand2_1
Xsky130_fd_sc_hs__nand2_1_48 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nor2_1_49/Y sky130_fd_sc_hs__nor2_1_47/B
+ sky130_fd_sc_hs__nor2_1_69/B sky130_fd_sc_hs__nand2_1_49/a_117_74# sky130_fd_sc_hs__nand2_1
Xsky130_fd_sc_hs__nand2_1_37 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nor2_1_29/Y sky130_fd_sc_hs__nor2_1_27/B
+ sky130_fd_sc_hs__inv_4_39/A sky130_fd_sc_hs__nand2_1_37/a_117_74# sky130_fd_sc_hs__nand2_1
Xsky130_fd_sc_hs__nand2_1_26 DVSS DVDD DVDD DVSS fine_control_avg_window_select[2]
+ sky130_fd_sc_hs__o22ai_1_1/A2 fine_control_avg_window_select[1] sky130_fd_sc_hs__nand2_1_27/a_117_74#
+ sky130_fd_sc_hs__nand2_1
Xsky130_fd_sc_hs__nand2_1_59 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_55/Y sky130_fd_sc_hs__nand2_1_59/Y
+ sky130_fd_sc_hs__nor2_1_59/A sky130_fd_sc_hs__nand2_1_59/a_117_74# sky130_fd_sc_hs__nand2_1
Xsky130_fd_sc_hs__dfxtp_4_5 DVSS DVDD DVDD DVSS out_star sky130_fd_sc_hs__dfxtp_4_5/D
+ clk_out sky130_fd_sc_hs__dfxtp_4_5/a_1226_296# sky130_fd_sc_hs__dfxtp_4_5/a_735_102#
+ sky130_fd_sc_hs__dfxtp_4_5/a_1141_508# sky130_fd_sc_hs__dfxtp_4_5/a_206_368# sky130_fd_sc_hs__dfxtp_4_5/a_437_503#
+ sky130_fd_sc_hs__dfxtp_4_5/a_27_74# sky130_fd_sc_hs__dfxtp_4_5/a_651_503# sky130_fd_sc_hs__dfxtp_4_5/a_696_458#
+ sky130_fd_sc_hs__dfxtp_4_5/a_544_485# sky130_fd_sc_hs__dfxtp_4_5/a_1178_124# sky130_fd_sc_hs__dfxtp_4_5/a_1034_424#
+ sky130_fd_sc_hs__dfxtp_4
Xsky130_fd_sc_hs__inv_2_6 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_2_7/A sky130_fd_sc_hs__inv_2_7/Y
+ sky130_fd_sc_hs__inv_2
Xsky130_fd_sc_hs__dfxtp_2_2 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_2_9/B sky130_fd_sc_hs__dfxtp_4_9/CLK
+ sky130_fd_sc_hs__inv_2_1/A sky130_fd_sc_hs__dfxtp_2_3/a_431_508# sky130_fd_sc_hs__dfxtp_2_3/a_1125_508#
+ sky130_fd_sc_hs__dfxtp_2_3/a_206_368# sky130_fd_sc_hs__dfxtp_2_3/a_27_74# sky130_fd_sc_hs__dfxtp_2_3/a_708_101#
+ sky130_fd_sc_hs__dfxtp_2_3/a_1019_424# sky130_fd_sc_hs__dfxtp_2_3/a_1172_124# sky130_fd_sc_hs__dfxtp_2_3/a_644_504#
+ sky130_fd_sc_hs__dfxtp_2_3/a_1217_314# sky130_fd_sc_hs__dfxtp_2_3/a_538_429# sky130_fd_sc_hs__dfxtp_2_3/a_695_459#
+ sky130_fd_sc_hs__dfxtp_2
Xsky130_fd_sc_hs__a21oi_1_104 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_103/A sky130_fd_sc_hs__nor3_1_7/A
+ sky130_fd_sc_hs__nand2_2_9/B sky130_fd_sc_hs__inv_4_121/Y sky130_fd_sc_hs__a21oi_1_105/a_117_74#
+ sky130_fd_sc_hs__a21oi_1_105/a_29_368# sky130_fd_sc_hs__a21oi_1
Xsky130_fd_sc_hs__a21oi_1_115 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__o21a_1_59/A2 sky130_fd_sc_hs__dfrtn_1_41/D
+ sky130_fd_sc_hs__o21a_1_71/B1 sky130_fd_sc_hs__inv_4_129/Y sky130_fd_sc_hs__a21oi_1_115/a_117_74#
+ sky130_fd_sc_hs__a21oi_1_115/a_29_368# sky130_fd_sc_hs__a21oi_1
Xsky130_fd_sc_hs__nand2_1_120 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__o21a_1_77/A2 sky130_fd_sc_hs__o21a_1_77/B1
+ sky130_fd_sc_hs__inv_4_113/A sky130_fd_sc_hs__nand2_1_121/a_117_74# sky130_fd_sc_hs__nand2_1
Xsky130_fd_sc_hs__maj3_1_2 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__maj3_1_3/A sky130_fd_sc_hs__maj3_1_3/B
+ sky130_fd_sc_hs__maj3_1_3/X sky130_fd_sc_hs__maj3_1_3/C sky130_fd_sc_hs__maj3_1_3/a_598_384#
+ sky130_fd_sc_hs__maj3_1_3/a_226_384# sky130_fd_sc_hs__maj3_1_3/a_84_74# sky130_fd_sc_hs__maj3_1_3/a_403_136#
+ sky130_fd_sc_hs__maj3_1_3/a_406_384# sky130_fd_sc_hs__maj3_1_3/a_595_136# sky130_fd_sc_hs__maj3_1_3/a_223_120#
+ sky130_fd_sc_hs__maj3_1
Xsky130_fd_sc_hs__nand2_2_7 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_2_7/Y sky130_fd_sc_hs__nand2_2_7/B
+ sky130_fd_sc_hs__inv_2_9/A sky130_fd_sc_hs__nand2_2_7/a_27_74# sky130_fd_sc_hs__nand2_2
Xsky130_fd_sc_hs__nor2_2_3 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nor2_2_3/B sky130_fd_sc_hs__nor2_2_3/Y
+ sky130_fd_sc_hs__nor2_2_3/A sky130_fd_sc_hs__nor2_2_3/a_35_368# sky130_fd_sc_hs__nor2_2
Xsky130_fd_sc_hs__nor2_1_12 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nor2_1_13/B sky130_fd_sc_hs__nor2_1_13/Y
+ sky130_fd_sc_hs__inv_4_17/Y sky130_fd_sc_hs__nor2_1_13/a_116_368# sky130_fd_sc_hs__nor2_1
Xsky130_fd_sc_hs__nor2_1_56 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nor2_1_57/B sky130_fd_sc_hs__nor2_1_57/Y
+ sky130_fd_sc_hs__inv_4_79/Y sky130_fd_sc_hs__nor2_1_57/a_116_368# sky130_fd_sc_hs__nor2_1
Xsky130_fd_sc_hs__nor2_1_45 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nor2_1_45/B sky130_fd_sc_hs__nor2_1_45/Y
+ sky130_fd_sc_hs__inv_4_63/Y sky130_fd_sc_hs__nor2_1_45/a_116_368# sky130_fd_sc_hs__nor2_1
Xsky130_fd_sc_hs__nor2_1_34 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nor2_1_35/B sky130_fd_sc_hs__nor2_1_35/Y
+ sky130_fd_sc_hs__inv_4_47/Y sky130_fd_sc_hs__nor2_1_35/a_116_368# sky130_fd_sc_hs__nor2_1
Xsky130_fd_sc_hs__nor2_1_23 DVSS DVDD DVDD DVSS fine_control_avg_window_select[2]
+ sky130_fd_sc_hs__nor2_1_23/Y fine_control_avg_window_select[1] sky130_fd_sc_hs__nor2_1_23/a_116_368#
+ sky130_fd_sc_hs__nor2_1
Xsky130_fd_sc_hs__nor2_1_89 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_87/A sky130_fd_sc_hs__nor2_1_89/Y
+ sky130_fd_sc_hs__nor2_1_89/A sky130_fd_sc_hs__nor2_1_89/a_116_368# sky130_fd_sc_hs__nor2_1
Xsky130_fd_sc_hs__nor2_1_78 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_95/Y sky130_fd_sc_hs__nor4_1_1/A
+ sky130_fd_sc_hs__xnor2_1_9/A sky130_fd_sc_hs__nor2_1_79/a_116_368# sky130_fd_sc_hs__nor2_1
Xsky130_fd_sc_hs__nor2_1_67 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_65/Y sky130_fd_sc_hs__nor3_1_1/C
+ sky130_fd_sc_hs__inv_4_89/A sky130_fd_sc_hs__nor2_1_67/a_116_368# sky130_fd_sc_hs__nor2_1
Xsky130_fd_sc_hs__xnor2_1_9 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__xnor2_1_9/A sky130_fd_sc_hs__xnor2_1_9/Y
+ sky130_fd_sc_hs__xnor2_1_9/B sky130_fd_sc_hs__xnor2_1_9/a_376_368# sky130_fd_sc_hs__xnor2_1_9/a_112_119#
+ sky130_fd_sc_hs__xnor2_1_9/a_138_385# sky130_fd_sc_hs__xnor2_1_9/a_293_74# sky130_fd_sc_hs__xnor2_1
Xsky130_fd_sc_hs__nor2b_1_23 DVSS DVDD DVDD DVSS fine_control_avg_window_select[4]
+ sky130_fd_sc_hs__nor2b_1_23/Y fine_control_avg_window_select[3] sky130_fd_sc_hs__nor2b_1_23/a_278_368#
+ sky130_fd_sc_hs__nor2b_1_23/a_27_112# sky130_fd_sc_hs__nor2b_1
Xsky130_fd_sc_hs__nor2b_1_12 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__fa_2_13/SUM sky130_fd_sc_hs__nor2b_1_13/Y
+ sky130_fd_sc_hs__or2_1_1/A sky130_fd_sc_hs__nor2b_1_13/a_278_368# sky130_fd_sc_hs__nor2b_1_13/a_27_112#
+ sky130_fd_sc_hs__nor2b_1
Xsky130_fd_sc_hs__nor2b_1_45 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__o21a_1_63/A1 sky130_fd_sc_hs__nor3_1_13/C
+ sky130_fd_sc_hs__o21a_1_59/A1 sky130_fd_sc_hs__nor2b_1_45/a_278_368# sky130_fd_sc_hs__nor2b_1_45/a_27_112#
+ sky130_fd_sc_hs__nor2b_1
Xsky130_fd_sc_hs__nor2b_1_34 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nor2b_1_29/Y sky130_fd_sc_hs__dfxtp_4_2/D
+ rst sky130_fd_sc_hs__nor2b_1_35/a_278_368# sky130_fd_sc_hs__nor2b_1_35/a_27_112#
+ sky130_fd_sc_hs__nor2b_1
Xsky130_fd_sc_hs__inv_4_104 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nor2_1_95/B sky130_fd_sc_hs__inv_4_105/A
+ sky130_fd_sc_hs__inv_4
Xsky130_fd_sc_hs__inv_4_115 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_115/Y sky130_fd_sc_hs__nor3_1_15/A
+ sky130_fd_sc_hs__inv_4
Xsky130_fd_sc_hs__inv_4_126 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__maj3_1_3/B sky130_fd_sc_hs__inv_4_127/A
+ sky130_fd_sc_hs__inv_4
Xsky130_fd_sc_hs__inv_4_137 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_137/Y sky130_fd_sc_hs__inv_4_137/A
+ sky130_fd_sc_hs__inv_4
Xsky130_fd_sc_hs__o22ai_1_4 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_81/Y sky130_fd_sc_hs__inv_4_71/A
+ sky130_fd_sc_hs__nor4_1_3/A sky130_fd_sc_hs__inv_4_83/Y sky130_fd_sc_hs__dfrbp_1_7/Q
+ sky130_fd_sc_hs__o22ai_1_5/a_340_368# sky130_fd_sc_hs__o22ai_1_5/a_142_368# sky130_fd_sc_hs__o22ai_1_5/a_27_74#
+ sky130_fd_sc_hs__o22ai_1
Xsky130_fd_sc_hs__conb_1_0 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__conb_1_1/LO sky130_fd_sc_hs__conb_1_1/HI
+ sky130_fd_sc_hs__conb_1_1/a_165_290# sky130_fd_sc_hs__conb_1_1/a_21_290# sky130_fd_sc_hs__conb_1
Xsky130_fd_sc_hs__nand2_4_15 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__o21ai_2_1/B1 div_ratio_half[4]
+ sky130_fd_sc_hs__inv_4_103/A sky130_fd_sc_hs__nand2_4_15/a_27_74# sky130_fd_sc_hs__nand2_4
Xsky130_fd_sc_hs__o22ai_1_10 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_113/Y sky130_fd_sc_hs__o21a_1_71/A1
+ sky130_fd_sc_hs__nor4_1_3/D sky130_fd_sc_hs__inv_4_115/Y sky130_fd_sc_hs__inv_4_99/A
+ sky130_fd_sc_hs__o22ai_1_11/a_340_368# sky130_fd_sc_hs__o22ai_1_11/a_142_368# sky130_fd_sc_hs__o22ai_1_11/a_27_74#
+ sky130_fd_sc_hs__o22ai_1
Xsky130_fd_sc_hs__and2_2_2 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_87/Y sky130_fd_sc_hs__nor2_2_1/Y
+ sky130_fd_sc_hs__inv_2_1/A sky130_fd_sc_hs__and2_2_3/a_31_74# sky130_fd_sc_hs__and2_2_3/a_118_74#
+ sky130_fd_sc_hs__and2_2
Xsky130_fd_sc_hs__inv_4_80 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_81/Y sky130_fd_sc_hs__inv_4_81/A
+ sky130_fd_sc_hs__inv_4
Xsky130_fd_sc_hs__inv_4_91 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__or3b_2_1/B sky130_fd_sc_hs__inv_4_91/A
+ sky130_fd_sc_hs__inv_4
Xsky130_fd_sc_hs__dfxtp_2_11 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__xnor2_1_7/A sky130_fd_sc_hs__dfxtp_4_9/CLK
+ sky130_fd_sc_hs__nor2_1_91/Y sky130_fd_sc_hs__dfxtp_2_11/a_431_508# sky130_fd_sc_hs__dfxtp_2_11/a_1125_508#
+ sky130_fd_sc_hs__dfxtp_2_11/a_206_368# sky130_fd_sc_hs__dfxtp_2_11/a_27_74# sky130_fd_sc_hs__dfxtp_2_11/a_708_101#
+ sky130_fd_sc_hs__dfxtp_2_11/a_1019_424# sky130_fd_sc_hs__dfxtp_2_11/a_1172_124#
+ sky130_fd_sc_hs__dfxtp_2_11/a_644_504# sky130_fd_sc_hs__dfxtp_2_11/a_1217_314# sky130_fd_sc_hs__dfxtp_2_11/a_538_429#
+ sky130_fd_sc_hs__dfxtp_2_11/a_695_459# sky130_fd_sc_hs__dfxtp_2
Xsky130_fd_sc_hs__a22o_1_27 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__a22o_1_27/X sky130_fd_sc_hs__dfrbp_1_1/Q
+ sky130_fd_sc_hs__inv_4_39/Y sky130_fd_sc_hs__inv_4_61/A sky130_fd_sc_hs__inv_4_37/Y
+ sky130_fd_sc_hs__a22o_1_27/a_222_392# sky130_fd_sc_hs__a22o_1_27/a_230_79# sky130_fd_sc_hs__a22o_1_27/a_52_123#
+ sky130_fd_sc_hs__a22o_1_27/a_132_392# sky130_fd_sc_hs__a22o_1
Xsky130_fd_sc_hs__a22o_1_16 DVSS DVDD DVDD DVSS osc_fine_con_final[6] manual_control_osc[6]
+ sky130_fd_sc_hs__inv_4_43/Y sky130_fd_sc_hs__fa_2_13/B fftl_en sky130_fd_sc_hs__a22o_1_17/a_222_392#
+ sky130_fd_sc_hs__a22o_1_17/a_230_79# sky130_fd_sc_hs__a22o_1_17/a_52_123# sky130_fd_sc_hs__a22o_1_17/a_132_392#
+ sky130_fd_sc_hs__a22o_1
Xsky130_fd_sc_hs__o21ai_1_3 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__o21ai_1_3/Y sky130_fd_sc_hs__o21ai_1_3/B1
+ sky130_fd_sc_hs__nor2_1_33/Y sky130_fd_sc_hs__and2_2_1/X sky130_fd_sc_hs__o21ai_1_3/a_162_368#
+ sky130_fd_sc_hs__o21ai_1_3/a_27_74# sky130_fd_sc_hs__o21ai_1
Xsky130_fd_sc_hs__nand2_1_49 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nor2_1_49/Y sky130_fd_sc_hs__nor2_1_47/B
+ sky130_fd_sc_hs__nor2_1_69/B sky130_fd_sc_hs__nand2_1_49/a_117_74# sky130_fd_sc_hs__nand2_1
Xsky130_fd_sc_hs__nand2_1_38 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nor2_1_27/Y sky130_fd_sc_hs__nor2_1_49/B
+ sky130_fd_sc_hs__inv_4_55/A sky130_fd_sc_hs__nand2_1_39/a_117_74# sky130_fd_sc_hs__nand2_1
Xsky130_fd_sc_hs__nand2_1_27 DVSS DVDD DVDD DVSS fine_control_avg_window_select[2]
+ sky130_fd_sc_hs__o22ai_1_1/A2 fine_control_avg_window_select[1] sky130_fd_sc_hs__nand2_1_27/a_117_74#
+ sky130_fd_sc_hs__nand2_1
Xsky130_fd_sc_hs__nand2_1_16 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nor2_1_7/Y sky130_fd_sc_hs__nor2_1_35/B
+ sky130_fd_sc_hs__o21a_1_15/A1 sky130_fd_sc_hs__nand2_1_17/a_117_74# sky130_fd_sc_hs__nand2_1
Xsky130_fd_sc_hs__dfxtp_4_6 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__dfxtp_4_7/Q sky130_fd_sc_hs__dfxtp_4_7/D
+ sky130_fd_sc_hs__inv_4_57/Y sky130_fd_sc_hs__dfxtp_4_7/a_1226_296# sky130_fd_sc_hs__dfxtp_4_7/a_735_102#
+ sky130_fd_sc_hs__dfxtp_4_7/a_1141_508# sky130_fd_sc_hs__dfxtp_4_7/a_206_368# sky130_fd_sc_hs__dfxtp_4_7/a_437_503#
+ sky130_fd_sc_hs__dfxtp_4_7/a_27_74# sky130_fd_sc_hs__dfxtp_4_7/a_651_503# sky130_fd_sc_hs__dfxtp_4_7/a_696_458#
+ sky130_fd_sc_hs__dfxtp_4_7/a_544_485# sky130_fd_sc_hs__dfxtp_4_7/a_1178_124# sky130_fd_sc_hs__dfxtp_4_7/a_1034_424#
+ sky130_fd_sc_hs__dfxtp_4
Xsky130_fd_sc_hs__inv_2_7 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_2_7/A sky130_fd_sc_hs__inv_2_7/Y
+ sky130_fd_sc_hs__inv_2
Xsky130_fd_sc_hs__dfxtp_2_3 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_2_9/B sky130_fd_sc_hs__dfxtp_4_9/CLK
+ sky130_fd_sc_hs__inv_2_1/A sky130_fd_sc_hs__dfxtp_2_3/a_431_508# sky130_fd_sc_hs__dfxtp_2_3/a_1125_508#
+ sky130_fd_sc_hs__dfxtp_2_3/a_206_368# sky130_fd_sc_hs__dfxtp_2_3/a_27_74# sky130_fd_sc_hs__dfxtp_2_3/a_708_101#
+ sky130_fd_sc_hs__dfxtp_2_3/a_1019_424# sky130_fd_sc_hs__dfxtp_2_3/a_1172_124# sky130_fd_sc_hs__dfxtp_2_3/a_644_504#
+ sky130_fd_sc_hs__dfxtp_2_3/a_1217_314# sky130_fd_sc_hs__dfxtp_2_3/a_538_429# sky130_fd_sc_hs__dfxtp_2_3/a_695_459#
+ sky130_fd_sc_hs__dfxtp_2
Xsky130_fd_sc_hs__a21oi_1_105 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_103/A sky130_fd_sc_hs__nor3_1_7/A
+ sky130_fd_sc_hs__nand2_2_9/B sky130_fd_sc_hs__inv_4_121/Y sky130_fd_sc_hs__a21oi_1_105/a_117_74#
+ sky130_fd_sc_hs__a21oi_1_105/a_29_368# sky130_fd_sc_hs__a21oi_1
Xsky130_fd_sc_hs__a21oi_1_116 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__o21a_1_69/A2 sky130_fd_sc_hs__dfrtn_1_39/D
+ sky130_fd_sc_hs__o21a_1_67/B1 sky130_fd_sc_hs__inv_4_125/Y sky130_fd_sc_hs__a21oi_1_117/a_117_74#
+ sky130_fd_sc_hs__a21oi_1_117/a_29_368# sky130_fd_sc_hs__a21oi_1
Xsky130_fd_sc_hs__nand2_1_110 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__o21a_1_71/A2 sky130_fd_sc_hs__o21a_1_71/B1
+ sky130_fd_sc_hs__o21a_1_71/A1 sky130_fd_sc_hs__nand2_1_111/a_117_74# sky130_fd_sc_hs__nand2_1
Xsky130_fd_sc_hs__nand2_1_121 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__o21a_1_77/A2 sky130_fd_sc_hs__o21a_1_77/B1
+ sky130_fd_sc_hs__inv_4_113/A sky130_fd_sc_hs__nand2_1_121/a_117_74# sky130_fd_sc_hs__nand2_1
Xsky130_fd_sc_hs__maj3_1_3 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__maj3_1_3/A sky130_fd_sc_hs__maj3_1_3/B
+ sky130_fd_sc_hs__maj3_1_3/X sky130_fd_sc_hs__maj3_1_3/C sky130_fd_sc_hs__maj3_1_3/a_598_384#
+ sky130_fd_sc_hs__maj3_1_3/a_226_384# sky130_fd_sc_hs__maj3_1_3/a_84_74# sky130_fd_sc_hs__maj3_1_3/a_403_136#
+ sky130_fd_sc_hs__maj3_1_3/a_406_384# sky130_fd_sc_hs__maj3_1_3/a_595_136# sky130_fd_sc_hs__maj3_1_3/a_223_120#
+ sky130_fd_sc_hs__maj3_1
Xsky130_fd_sc_hs__nand2_2_8 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand3_1_1/A sky130_fd_sc_hs__nand2_2_9/B
+ sky130_fd_sc_hs__inv_2_7/Y sky130_fd_sc_hs__nand2_2_9/a_27_74# sky130_fd_sc_hs__nand2_2
Xsky130_fd_sc_hs__nor2_1_13 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nor2_1_13/B sky130_fd_sc_hs__nor2_1_13/Y
+ sky130_fd_sc_hs__inv_4_17/Y sky130_fd_sc_hs__nor2_1_13/a_116_368# sky130_fd_sc_hs__nor2_1
Xsky130_fd_sc_hs__nor2_1_46 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nor2_1_47/B sky130_fd_sc_hs__nor2_1_47/Y
+ sky130_fd_sc_hs__inv_4_65/Y sky130_fd_sc_hs__nor2_1_47/a_116_368# sky130_fd_sc_hs__nor2_1
Xsky130_fd_sc_hs__nor2_1_35 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nor2_1_35/B sky130_fd_sc_hs__nor2_1_35/Y
+ sky130_fd_sc_hs__inv_4_47/Y sky130_fd_sc_hs__nor2_1_35/a_116_368# sky130_fd_sc_hs__nor2_1
Xsky130_fd_sc_hs__nor2_1_24 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nor2_1_25/B sky130_fd_sc_hs__nor2_1_25/Y
+ sky130_fd_sc_hs__inv_4_41/Y sky130_fd_sc_hs__nor2_1_25/a_116_368# sky130_fd_sc_hs__nor2_1
Xsky130_fd_sc_hs__nor2_1_79 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_95/Y sky130_fd_sc_hs__nor4_1_1/A
+ sky130_fd_sc_hs__xnor2_1_9/A sky130_fd_sc_hs__nor2_1_79/a_116_368# sky130_fd_sc_hs__nor2_1
Xsky130_fd_sc_hs__nor2_1_68 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nor2_1_69/B sky130_fd_sc_hs__nor3_1_1/B
+ sky130_fd_sc_hs__inv_4_69/Y sky130_fd_sc_hs__nor2_1_69/a_116_368# sky130_fd_sc_hs__nor2_1
Xsky130_fd_sc_hs__nor2_1_57 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nor2_1_57/B sky130_fd_sc_hs__nor2_1_57/Y
+ sky130_fd_sc_hs__inv_4_79/Y sky130_fd_sc_hs__nor2_1_57/a_116_368# sky130_fd_sc_hs__nor2_1
Xsky130_fd_sc_hs__nor2b_1_13 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__fa_2_13/SUM sky130_fd_sc_hs__nor2b_1_13/Y
+ sky130_fd_sc_hs__or2_1_1/A sky130_fd_sc_hs__nor2b_1_13/a_278_368# sky130_fd_sc_hs__nor2b_1_13/a_27_112#
+ sky130_fd_sc_hs__nor2b_1
Xsky130_fd_sc_hs__nor2b_1_46 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__o21a_1_59/A1 sky130_fd_sc_hs__nor3_1_1/A
+ sky130_fd_sc_hs__o21a_1_63/A1 sky130_fd_sc_hs__nor2b_1_47/a_278_368# sky130_fd_sc_hs__nor2b_1_47/a_27_112#
+ sky130_fd_sc_hs__nor2b_1
Xsky130_fd_sc_hs__nor2b_1_35 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nor2b_1_29/Y sky130_fd_sc_hs__dfxtp_4_2/D
+ rst sky130_fd_sc_hs__nor2b_1_35/a_278_368# sky130_fd_sc_hs__nor2b_1_35/a_27_112#
+ sky130_fd_sc_hs__nor2b_1
Xsky130_fd_sc_hs__nor2b_1_24 DVSS DVDD DVDD DVSS fine_control_avg_window_select[3]
+ sky130_fd_sc_hs__nor2b_1_25/Y fine_control_avg_window_select[4] sky130_fd_sc_hs__nor2b_1_25/a_278_368#
+ sky130_fd_sc_hs__nor2b_1_25/a_27_112# sky130_fd_sc_hs__nor2b_1
Xsky130_fd_sc_hs__inv_4_105 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nor2_1_95/B sky130_fd_sc_hs__inv_4_105/A
+ sky130_fd_sc_hs__inv_4
Xsky130_fd_sc_hs__inv_4_116 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_117/Y sky130_fd_sc_hs__nor2_1_97/A
+ sky130_fd_sc_hs__inv_4
Xsky130_fd_sc_hs__inv_4_127 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__maj3_1_3/B sky130_fd_sc_hs__inv_4_127/A
+ sky130_fd_sc_hs__inv_4
Xsky130_fd_sc_hs__o22ai_1_5 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_81/Y sky130_fd_sc_hs__inv_4_71/A
+ sky130_fd_sc_hs__nor4_1_3/A sky130_fd_sc_hs__inv_4_83/Y sky130_fd_sc_hs__dfrbp_1_7/Q
+ sky130_fd_sc_hs__o22ai_1_5/a_340_368# sky130_fd_sc_hs__o22ai_1_5/a_142_368# sky130_fd_sc_hs__o22ai_1_5/a_27_74#
+ sky130_fd_sc_hs__o22ai_1
Xsky130_fd_sc_hs__conb_1_1 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__conb_1_1/LO sky130_fd_sc_hs__conb_1_1/HI
+ sky130_fd_sc_hs__conb_1_1/a_165_290# sky130_fd_sc_hs__conb_1_1/a_21_290# sky130_fd_sc_hs__conb_1
Xsky130_fd_sc_hs__o22ai_1_11 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_113/Y sky130_fd_sc_hs__o21a_1_71/A1
+ sky130_fd_sc_hs__nor4_1_3/D sky130_fd_sc_hs__inv_4_115/Y sky130_fd_sc_hs__inv_4_99/A
+ sky130_fd_sc_hs__o22ai_1_11/a_340_368# sky130_fd_sc_hs__o22ai_1_11/a_142_368# sky130_fd_sc_hs__o22ai_1_11/a_27_74#
+ sky130_fd_sc_hs__o22ai_1
Xsky130_fd_sc_hs__and2_2_3 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_87/Y sky130_fd_sc_hs__nor2_2_1/Y
+ sky130_fd_sc_hs__inv_2_1/A sky130_fd_sc_hs__and2_2_3/a_31_74# sky130_fd_sc_hs__and2_2_3/a_118_74#
+ sky130_fd_sc_hs__and2_2
Xsky130_fd_sc_hs__inv_4_81 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_81/Y sky130_fd_sc_hs__inv_4_81/A
+ sky130_fd_sc_hs__inv_4
Xsky130_fd_sc_hs__inv_4_70 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_71/Y sky130_fd_sc_hs__inv_4_71/A
+ sky130_fd_sc_hs__inv_4
Xsky130_fd_sc_hs__inv_4_92 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__maj3_1_1/C sky130_fd_sc_hs__inv_4_93/A
+ sky130_fd_sc_hs__inv_4
Xsky130_fd_sc_hs__a22o_1_28 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__a22o_1_29/X sky130_fd_sc_hs__o22ai_1_7/A1
+ sky130_fd_sc_hs__inv_4_97/Y sky130_fd_sc_hs__nor2_1_97/A sky130_fd_sc_hs__nor2_1_99/A
+ sky130_fd_sc_hs__a22o_1_29/a_222_392# sky130_fd_sc_hs__a22o_1_29/a_230_79# sky130_fd_sc_hs__a22o_1_29/a_52_123#
+ sky130_fd_sc_hs__a22o_1_29/a_132_392# sky130_fd_sc_hs__a22o_1
Xsky130_fd_sc_hs__a22o_1_17 DVSS DVDD DVDD DVSS osc_fine_con_final[6] manual_control_osc[6]
+ sky130_fd_sc_hs__inv_4_43/Y sky130_fd_sc_hs__fa_2_13/B fftl_en sky130_fd_sc_hs__a22o_1_17/a_222_392#
+ sky130_fd_sc_hs__a22o_1_17/a_230_79# sky130_fd_sc_hs__a22o_1_17/a_52_123# sky130_fd_sc_hs__a22o_1_17/a_132_392#
+ sky130_fd_sc_hs__a22o_1
Xsky130_fd_sc_hs__o21ai_1_4 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__o21ai_1_5/Y sky130_fd_sc_hs__o21ai_1_5/B1
+ sky130_fd_sc_hs__inv_4_51/Y sky130_fd_sc_hs__inv_4_53/A sky130_fd_sc_hs__o21ai_1_5/a_162_368#
+ sky130_fd_sc_hs__o21ai_1_5/a_27_74# sky130_fd_sc_hs__o21ai_1
Xsky130_fd_sc_hs__nand2_1_39 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nor2_1_27/Y sky130_fd_sc_hs__nor2_1_49/B
+ sky130_fd_sc_hs__inv_4_55/A sky130_fd_sc_hs__nand2_1_39/a_117_74# sky130_fd_sc_hs__nand2_1
Xsky130_fd_sc_hs__nand2_1_28 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__and2_2_1/X sky130_fd_sc_hs__inv_4_25/A
+ sky130_fd_sc_hs__o21a_1_23/A1 sky130_fd_sc_hs__nand2_1_29/a_117_74# sky130_fd_sc_hs__nand2_1
Xsky130_fd_sc_hs__nand2_1_17 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nor2_1_7/Y sky130_fd_sc_hs__nor2_1_35/B
+ sky130_fd_sc_hs__o21a_1_15/A1 sky130_fd_sc_hs__nand2_1_17/a_117_74# sky130_fd_sc_hs__nand2_1
Xsky130_fd_sc_hs__nand3_1_0 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand3_1_1/C sky130_fd_sc_hs__nand4_2_1/B
+ sky130_fd_sc_hs__nand3_1_1/B sky130_fd_sc_hs__nand3_1_1/A sky130_fd_sc_hs__nand3_1_1/a_155_74#
+ sky130_fd_sc_hs__nand3_1_1/a_233_74# sky130_fd_sc_hs__nand3_1
Xsky130_fd_sc_hs__dfxtp_4_7 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__dfxtp_4_7/Q sky130_fd_sc_hs__dfxtp_4_7/D
+ sky130_fd_sc_hs__inv_4_57/Y sky130_fd_sc_hs__dfxtp_4_7/a_1226_296# sky130_fd_sc_hs__dfxtp_4_7/a_735_102#
+ sky130_fd_sc_hs__dfxtp_4_7/a_1141_508# sky130_fd_sc_hs__dfxtp_4_7/a_206_368# sky130_fd_sc_hs__dfxtp_4_7/a_437_503#
+ sky130_fd_sc_hs__dfxtp_4_7/a_27_74# sky130_fd_sc_hs__dfxtp_4_7/a_651_503# sky130_fd_sc_hs__dfxtp_4_7/a_696_458#
+ sky130_fd_sc_hs__dfxtp_4_7/a_544_485# sky130_fd_sc_hs__dfxtp_4_7/a_1178_124# sky130_fd_sc_hs__dfxtp_4_7/a_1034_424#
+ sky130_fd_sc_hs__dfxtp_4
Xsky130_fd_sc_hs__inv_2_8 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_2_9/A sky130_fd_sc_hs__inv_2_9/Y
+ sky130_fd_sc_hs__inv_2
Xsky130_fd_sc_hs__dfxtp_2_4 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_2_3/A sky130_fd_sc_hs__dfxtp_4_9/CLK
+ sky130_fd_sc_hs__dfxtp_2_5/D sky130_fd_sc_hs__dfxtp_2_5/a_431_508# sky130_fd_sc_hs__dfxtp_2_5/a_1125_508#
+ sky130_fd_sc_hs__dfxtp_2_5/a_206_368# sky130_fd_sc_hs__dfxtp_2_5/a_27_74# sky130_fd_sc_hs__dfxtp_2_5/a_708_101#
+ sky130_fd_sc_hs__dfxtp_2_5/a_1019_424# sky130_fd_sc_hs__dfxtp_2_5/a_1172_124# sky130_fd_sc_hs__dfxtp_2_5/a_644_504#
+ sky130_fd_sc_hs__dfxtp_2_5/a_1217_314# sky130_fd_sc_hs__dfxtp_2_5/a_538_429# sky130_fd_sc_hs__dfxtp_2_5/a_695_459#
+ sky130_fd_sc_hs__dfxtp_2
Xsky130_fd_sc_hs__a21oi_1_106 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__o21a_1_67/A2 sky130_fd_sc_hs__dfrtn_1_33/D
+ sky130_fd_sc_hs__o21a_1_57/B1 sky130_fd_sc_hs__nor2_1_95/B sky130_fd_sc_hs__a21oi_1_107/a_117_74#
+ sky130_fd_sc_hs__a21oi_1_107/a_29_368# sky130_fd_sc_hs__a21oi_1
Xsky130_fd_sc_hs__a21oi_1_117 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__o21a_1_69/A2 sky130_fd_sc_hs__dfrtn_1_39/D
+ sky130_fd_sc_hs__o21a_1_67/B1 sky130_fd_sc_hs__inv_4_125/Y sky130_fd_sc_hs__a21oi_1_117/a_117_74#
+ sky130_fd_sc_hs__a21oi_1_117/a_29_368# sky130_fd_sc_hs__a21oi_1
Xsky130_fd_sc_hs__nand2_1_100 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__o21a_1_67/A2 sky130_fd_sc_hs__o21a_1_67/B1
+ sky130_fd_sc_hs__inv_4_133/A sky130_fd_sc_hs__nand2_1_101/a_117_74# sky130_fd_sc_hs__nand2_1
Xsky130_fd_sc_hs__nand2_1_111 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__o21a_1_71/A2 sky130_fd_sc_hs__o21a_1_71/B1
+ sky130_fd_sc_hs__o21a_1_71/A1 sky130_fd_sc_hs__nand2_1_111/a_117_74# sky130_fd_sc_hs__nand2_1
Xsky130_fd_sc_hs__nand2_2_9 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand3_1_1/A sky130_fd_sc_hs__nand2_2_9/B
+ sky130_fd_sc_hs__inv_2_7/Y sky130_fd_sc_hs__nand2_2_9/a_27_74# sky130_fd_sc_hs__nand2_2
Xsky130_fd_sc_hs__nor2_1_47 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nor2_1_47/B sky130_fd_sc_hs__nor2_1_47/Y
+ sky130_fd_sc_hs__inv_4_65/Y sky130_fd_sc_hs__nor2_1_47/a_116_368# sky130_fd_sc_hs__nor2_1
Xsky130_fd_sc_hs__nor2_1_36 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nor2_1_37/B sky130_fd_sc_hs__nor2_1_37/Y
+ sky130_fd_sc_hs__inv_4_35/Y sky130_fd_sc_hs__nor2_1_37/a_116_368# sky130_fd_sc_hs__nor2_1
Xsky130_fd_sc_hs__nor2_1_25 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nor2_1_25/B sky130_fd_sc_hs__nor2_1_25/Y
+ sky130_fd_sc_hs__inv_4_41/Y sky130_fd_sc_hs__nor2_1_25/a_116_368# sky130_fd_sc_hs__nor2_1
Xsky130_fd_sc_hs__nor2_1_14 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nor2_1_15/B sky130_fd_sc_hs__nor2_1_15/Y
+ sky130_fd_sc_hs__inv_4_19/Y sky130_fd_sc_hs__nor2_1_15/a_116_368# sky130_fd_sc_hs__nor2_1
Xsky130_fd_sc_hs__nor2_1_69 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nor2_1_69/B sky130_fd_sc_hs__nor3_1_1/B
+ sky130_fd_sc_hs__inv_4_69/Y sky130_fd_sc_hs__nor2_1_69/a_116_368# sky130_fd_sc_hs__nor2_1
Xsky130_fd_sc_hs__nor2_1_58 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_55/Y sky130_fd_sc_hs__nor4_1_1/D
+ sky130_fd_sc_hs__nor2_1_59/A sky130_fd_sc_hs__nor2_1_59/a_116_368# sky130_fd_sc_hs__nor2_1
Xsky130_fd_sc_hs__nor2b_1_14 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__fa_2_15/SUM sky130_fd_sc_hs__nor2b_1_15/Y
+ sky130_fd_sc_hs__or2_1_1/A sky130_fd_sc_hs__nor2b_1_15/a_278_368# sky130_fd_sc_hs__nor2b_1_15/a_27_112#
+ sky130_fd_sc_hs__nor2b_1
Xsky130_fd_sc_hs__nor2b_1_47 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__o21a_1_59/A1 sky130_fd_sc_hs__nor3_1_1/A
+ sky130_fd_sc_hs__o21a_1_63/A1 sky130_fd_sc_hs__nor2b_1_47/a_278_368# sky130_fd_sc_hs__nor2b_1_47/a_27_112#
+ sky130_fd_sc_hs__nor2b_1
Xsky130_fd_sc_hs__nor2b_1_36 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nor2b_1_29/Y sky130_fd_sc_hs__dfxtp_4_7/D
+ rst sky130_fd_sc_hs__nor2b_1_37/a_278_368# sky130_fd_sc_hs__nor2b_1_37/a_27_112#
+ sky130_fd_sc_hs__nor2b_1
Xsky130_fd_sc_hs__nor2b_1_25 DVSS DVDD DVDD DVSS fine_control_avg_window_select[3]
+ sky130_fd_sc_hs__nor2b_1_25/Y fine_control_avg_window_select[4] sky130_fd_sc_hs__nor2b_1_25/a_278_368#
+ sky130_fd_sc_hs__nor2b_1_25/a_27_112# sky130_fd_sc_hs__nor2b_1
Xsky130_fd_sc_hs__inv_4_106 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_107/Y sky130_fd_sc_hs__nor2_1_95/A
+ sky130_fd_sc_hs__inv_4
Xsky130_fd_sc_hs__inv_4_117 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_117/Y sky130_fd_sc_hs__nor2_1_97/A
+ sky130_fd_sc_hs__inv_4
Xsky130_fd_sc_hs__inv_4_128 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_129/Y sky130_fd_sc_hs__inv_4_129/A
+ sky130_fd_sc_hs__inv_4
Xsky130_fd_sc_hs__o22ai_1_6 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_75/Y sky130_fd_sc_hs__inv_4_85/A
+ sky130_fd_sc_hs__nor4_1_3/C sky130_fd_sc_hs__inv_4_97/Y sky130_fd_sc_hs__o22ai_1_7/A1
+ sky130_fd_sc_hs__o22ai_1_7/a_340_368# sky130_fd_sc_hs__o22ai_1_7/a_142_368# sky130_fd_sc_hs__o22ai_1_7/a_27_74#
+ sky130_fd_sc_hs__o22ai_1
Xsky130_fd_sc_hs__conb_1_2 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__conb_1_3/LO sky130_fd_sc_hs__conb_1_3/HI
+ sky130_fd_sc_hs__conb_1_3/a_165_290# sky130_fd_sc_hs__conb_1_3/a_21_290# sky130_fd_sc_hs__conb_1
Xsky130_fd_sc_hs__dfrtp_4_0 DVSS DVDD sky130_fd_sc_hs__clkbuf_8_1/X DVDD DVSS sky130_fd_sc_hs__inv_4_1/Y
+ sky130_fd_sc_hs__nand2_1_47/B sky130_fd_sc_hs__inv_4_1/A sky130_fd_sc_hs__dfrtp_4_1/a_37_78#
+ sky130_fd_sc_hs__dfrtp_4_1/a_494_366# sky130_fd_sc_hs__dfrtp_4_1/a_699_463# sky130_fd_sc_hs__dfrtp_4_1/a_313_74#
+ sky130_fd_sc_hs__dfrtp_4_1/a_1627_493# sky130_fd_sc_hs__dfrtp_4_1/a_1678_395# sky130_fd_sc_hs__dfrtp_4_1/a_1827_81#
+ sky130_fd_sc_hs__dfrtp_4_1/a_789_463# sky130_fd_sc_hs__dfrtp_4_1/a_1350_392# sky130_fd_sc_hs__dfrtp_4_1/a_834_355#
+ sky130_fd_sc_hs__dfrtp_4_1/a_812_138# sky130_fd_sc_hs__dfrtp_4_1/a_124_78# sky130_fd_sc_hs__dfrtp_4_1/a_1647_81#
+ sky130_fd_sc_hs__dfrtp_4_1/a_2010_409# sky130_fd_sc_hs__dfrtp_4_1/a_890_138# sky130_fd_sc_hs__dfrtp_4
Xsky130_fd_sc_hs__and2_2_4 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_2_3/A sky130_fd_sc_hs__inv_2_5/A
+ sky130_fd_sc_hs__and2_2_5/X sky130_fd_sc_hs__and2_2_5/a_31_74# sky130_fd_sc_hs__and2_2_5/a_118_74#
+ sky130_fd_sc_hs__and2_2
Xsky130_fd_sc_hs__inv_4_71 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_71/Y sky130_fd_sc_hs__inv_4_71/A
+ sky130_fd_sc_hs__inv_4
Xsky130_fd_sc_hs__inv_4_60 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_61/Y sky130_fd_sc_hs__inv_4_61/A
+ sky130_fd_sc_hs__inv_4
Xsky130_fd_sc_hs__inv_4_93 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__maj3_1_1/C sky130_fd_sc_hs__inv_4_93/A
+ sky130_fd_sc_hs__inv_4
Xsky130_fd_sc_hs__inv_4_82 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_83/Y sky130_fd_sc_hs__inv_4_83/A
+ sky130_fd_sc_hs__inv_4
Xsky130_fd_sc_hs__a22o_1_29 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__a22o_1_29/X sky130_fd_sc_hs__o22ai_1_7/A1
+ sky130_fd_sc_hs__inv_4_97/Y sky130_fd_sc_hs__nor2_1_97/A sky130_fd_sc_hs__nor2_1_99/A
+ sky130_fd_sc_hs__a22o_1_29/a_222_392# sky130_fd_sc_hs__a22o_1_29/a_230_79# sky130_fd_sc_hs__a22o_1_29/a_52_123#
+ sky130_fd_sc_hs__a22o_1_29/a_132_392# sky130_fd_sc_hs__a22o_1
Xsky130_fd_sc_hs__a22o_1_18 DVSS DVDD DVDD DVSS osc_fine_con_final[7] manual_control_osc[7]
+ sky130_fd_sc_hs__inv_4_43/Y sky130_fd_sc_hs__fa_2_17/B fftl_en sky130_fd_sc_hs__a22o_1_19/a_222_392#
+ sky130_fd_sc_hs__a22o_1_19/a_230_79# sky130_fd_sc_hs__a22o_1_19/a_52_123# sky130_fd_sc_hs__a22o_1_19/a_132_392#
+ sky130_fd_sc_hs__a22o_1
Xsky130_fd_sc_hs__o21ai_1_5 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__o21ai_1_5/Y sky130_fd_sc_hs__o21ai_1_5/B1
+ sky130_fd_sc_hs__inv_4_51/Y sky130_fd_sc_hs__inv_4_53/A sky130_fd_sc_hs__o21ai_1_5/a_162_368#
+ sky130_fd_sc_hs__o21ai_1_5/a_27_74# sky130_fd_sc_hs__o21ai_1
Xsky130_fd_sc_hs__nand2_1_29 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__and2_2_1/X sky130_fd_sc_hs__inv_4_25/A
+ sky130_fd_sc_hs__o21a_1_23/A1 sky130_fd_sc_hs__nand2_1_29/a_117_74# sky130_fd_sc_hs__nand2_1
Xsky130_fd_sc_hs__nand2_1_18 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nor2_1_21/Y sky130_fd_sc_hs__nor2_1_15/B
+ sky130_fd_sc_hs__o21a_1_17/A1 sky130_fd_sc_hs__nand2_1_19/a_117_74# sky130_fd_sc_hs__nand2_1
Xsky130_fd_sc_hs__nand3_1_1 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand3_1_1/C sky130_fd_sc_hs__nand4_2_1/B
+ sky130_fd_sc_hs__nand3_1_1/B sky130_fd_sc_hs__nand3_1_1/A sky130_fd_sc_hs__nand3_1_1/a_155_74#
+ sky130_fd_sc_hs__nand3_1_1/a_233_74# sky130_fd_sc_hs__nand3_1
Xsky130_fd_sc_hs__inv_2_9 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_2_9/A sky130_fd_sc_hs__inv_2_9/Y
+ sky130_fd_sc_hs__inv_2
Xsky130_fd_sc_hs__dfxtp_4_8 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_103/A sky130_fd_sc_hs__nor2_1_89/Y
+ sky130_fd_sc_hs__dfxtp_4_9/CLK sky130_fd_sc_hs__dfxtp_4_9/a_1226_296# sky130_fd_sc_hs__dfxtp_4_9/a_735_102#
+ sky130_fd_sc_hs__dfxtp_4_9/a_1141_508# sky130_fd_sc_hs__dfxtp_4_9/a_206_368# sky130_fd_sc_hs__dfxtp_4_9/a_437_503#
+ sky130_fd_sc_hs__dfxtp_4_9/a_27_74# sky130_fd_sc_hs__dfxtp_4_9/a_651_503# sky130_fd_sc_hs__dfxtp_4_9/a_696_458#
+ sky130_fd_sc_hs__dfxtp_4_9/a_544_485# sky130_fd_sc_hs__dfxtp_4_9/a_1178_124# sky130_fd_sc_hs__dfxtp_4_9/a_1034_424#
+ sky130_fd_sc_hs__dfxtp_4
Xsky130_fd_sc_hs__dfxtp_2_5 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_2_3/A sky130_fd_sc_hs__dfxtp_4_9/CLK
+ sky130_fd_sc_hs__dfxtp_2_5/D sky130_fd_sc_hs__dfxtp_2_5/a_431_508# sky130_fd_sc_hs__dfxtp_2_5/a_1125_508#
+ sky130_fd_sc_hs__dfxtp_2_5/a_206_368# sky130_fd_sc_hs__dfxtp_2_5/a_27_74# sky130_fd_sc_hs__dfxtp_2_5/a_708_101#
+ sky130_fd_sc_hs__dfxtp_2_5/a_1019_424# sky130_fd_sc_hs__dfxtp_2_5/a_1172_124# sky130_fd_sc_hs__dfxtp_2_5/a_644_504#
+ sky130_fd_sc_hs__dfxtp_2_5/a_1217_314# sky130_fd_sc_hs__dfxtp_2_5/a_538_429# sky130_fd_sc_hs__dfxtp_2_5/a_695_459#
+ sky130_fd_sc_hs__dfxtp_2
Xsky130_fd_sc_hs__a21oi_1_107 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__o21a_1_67/A2 sky130_fd_sc_hs__dfrtn_1_33/D
+ sky130_fd_sc_hs__o21a_1_57/B1 sky130_fd_sc_hs__nor2_1_95/B sky130_fd_sc_hs__a21oi_1_107/a_117_74#
+ sky130_fd_sc_hs__a21oi_1_107/a_29_368# sky130_fd_sc_hs__a21oi_1
Xsky130_fd_sc_hs__a21oi_1_118 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__o21a_1_77/A2 sky130_fd_sc_hs__dfrbp_1_37/D
+ sky130_fd_sc_hs__o21a_1_73/B1 sky130_fd_sc_hs__inv_4_115/Y sky130_fd_sc_hs__a21oi_1_119/a_117_74#
+ sky130_fd_sc_hs__a21oi_1_119/a_29_368# sky130_fd_sc_hs__a21oi_1
Xsky130_fd_sc_hs__nand2_1_101 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__o21a_1_67/A2 sky130_fd_sc_hs__o21a_1_67/B1
+ sky130_fd_sc_hs__inv_4_133/A sky130_fd_sc_hs__nand2_1_101/a_117_74# sky130_fd_sc_hs__nand2_1
Xsky130_fd_sc_hs__nand2_1_112 DVSS DVDD DVDD DVSS div_ratio_half[3] sky130_fd_sc_hs__nand4_2_1/D
+ sky130_fd_sc_hs__inv_2_7/Y sky130_fd_sc_hs__nand2_1_113/a_117_74# sky130_fd_sc_hs__nand2_1
Xsky130_fd_sc_hs__nor2_1_37 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nor2_1_37/B sky130_fd_sc_hs__nor2_1_37/Y
+ sky130_fd_sc_hs__inv_4_35/Y sky130_fd_sc_hs__nor2_1_37/a_116_368# sky130_fd_sc_hs__nor2_1
Xsky130_fd_sc_hs__nor2_1_26 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nor2_1_27/B sky130_fd_sc_hs__nor2_1_27/Y
+ sky130_fd_sc_hs__inv_4_37/Y sky130_fd_sc_hs__nor2_1_27/a_116_368# sky130_fd_sc_hs__nor2_1
Xsky130_fd_sc_hs__nor2_1_15 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nor2_1_15/B sky130_fd_sc_hs__nor2_1_15/Y
+ sky130_fd_sc_hs__inv_4_19/Y sky130_fd_sc_hs__nor2_1_15/a_116_368# sky130_fd_sc_hs__nor2_1
Xsky130_fd_sc_hs__nor2_1_59 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_55/Y sky130_fd_sc_hs__nor4_1_1/D
+ sky130_fd_sc_hs__nor2_1_59/A sky130_fd_sc_hs__nor2_1_59/a_116_368# sky130_fd_sc_hs__nor2_1
Xsky130_fd_sc_hs__nor2_1_48 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nor2_1_49/B sky130_fd_sc_hs__nor2_1_49/Y
+ sky130_fd_sc_hs__inv_4_59/Y sky130_fd_sc_hs__nor2_1_49/a_116_368# sky130_fd_sc_hs__nor2_1
Xsky130_fd_sc_hs__nor2b_1_37 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nor2b_1_29/Y sky130_fd_sc_hs__dfxtp_4_7/D
+ rst sky130_fd_sc_hs__nor2b_1_37/a_278_368# sky130_fd_sc_hs__nor2b_1_37/a_27_112#
+ sky130_fd_sc_hs__nor2b_1
Xsky130_fd_sc_hs__nor2b_1_26 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__fa_2_19/SUM sky130_fd_sc_hs__nor2b_1_27/Y
+ sky130_fd_sc_hs__or2_1_1/A sky130_fd_sc_hs__nor2b_1_27/a_278_368# sky130_fd_sc_hs__nor2b_1_27/a_27_112#
+ sky130_fd_sc_hs__nor2b_1
Xsky130_fd_sc_hs__nor2b_1_15 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__fa_2_15/SUM sky130_fd_sc_hs__nor2b_1_15/Y
+ sky130_fd_sc_hs__or2_1_1/A sky130_fd_sc_hs__nor2b_1_15/a_278_368# sky130_fd_sc_hs__nor2b_1_15/a_27_112#
+ sky130_fd_sc_hs__nor2b_1
Xsky130_fd_sc_hs__nor2b_1_48 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__o21a_1_71/A1 sky130_fd_sc_hs__nor3_1_13/A
+ sky130_fd_sc_hs__inv_4_113/A sky130_fd_sc_hs__nor2b_1_49/a_278_368# sky130_fd_sc_hs__nor2b_1_49/a_27_112#
+ sky130_fd_sc_hs__nor2b_1
Xsky130_fd_sc_hs__inv_4_107 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_107/Y sky130_fd_sc_hs__nor2_1_95/A
+ sky130_fd_sc_hs__inv_4
Xsky130_fd_sc_hs__inv_4_118 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_87/A sky130_fd_sc_hs__nand4_2_1/Y
+ sky130_fd_sc_hs__inv_4
Xsky130_fd_sc_hs__inv_4_129 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_129/Y sky130_fd_sc_hs__inv_4_129/A
+ sky130_fd_sc_hs__inv_4
Xsky130_fd_sc_hs__o22ai_1_7 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_75/Y sky130_fd_sc_hs__inv_4_85/A
+ sky130_fd_sc_hs__nor4_1_3/C sky130_fd_sc_hs__inv_4_97/Y sky130_fd_sc_hs__o22ai_1_7/A1
+ sky130_fd_sc_hs__o22ai_1_7/a_340_368# sky130_fd_sc_hs__o22ai_1_7/a_142_368# sky130_fd_sc_hs__o22ai_1_7/a_27_74#
+ sky130_fd_sc_hs__o22ai_1
Xsky130_fd_sc_hs__conb_1_3 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__conb_1_3/LO sky130_fd_sc_hs__conb_1_3/HI
+ sky130_fd_sc_hs__conb_1_3/a_165_290# sky130_fd_sc_hs__conb_1_3/a_21_290# sky130_fd_sc_hs__conb_1
Xsky130_fd_sc_hs__dfrtp_4_1 DVSS DVDD sky130_fd_sc_hs__clkbuf_8_1/X DVDD DVSS sky130_fd_sc_hs__inv_4_1/Y
+ sky130_fd_sc_hs__nand2_1_47/B sky130_fd_sc_hs__inv_4_1/A sky130_fd_sc_hs__dfrtp_4_1/a_37_78#
+ sky130_fd_sc_hs__dfrtp_4_1/a_494_366# sky130_fd_sc_hs__dfrtp_4_1/a_699_463# sky130_fd_sc_hs__dfrtp_4_1/a_313_74#
+ sky130_fd_sc_hs__dfrtp_4_1/a_1627_493# sky130_fd_sc_hs__dfrtp_4_1/a_1678_395# sky130_fd_sc_hs__dfrtp_4_1/a_1827_81#
+ sky130_fd_sc_hs__dfrtp_4_1/a_789_463# sky130_fd_sc_hs__dfrtp_4_1/a_1350_392# sky130_fd_sc_hs__dfrtp_4_1/a_834_355#
+ sky130_fd_sc_hs__dfrtp_4_1/a_812_138# sky130_fd_sc_hs__dfrtp_4_1/a_124_78# sky130_fd_sc_hs__dfrtp_4_1/a_1647_81#
+ sky130_fd_sc_hs__dfrtp_4_1/a_2010_409# sky130_fd_sc_hs__dfrtp_4_1/a_890_138# sky130_fd_sc_hs__dfrtp_4
Xsky130_fd_sc_hs__and2_2_5 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_2_3/A sky130_fd_sc_hs__inv_2_5/A
+ sky130_fd_sc_hs__and2_2_5/X sky130_fd_sc_hs__and2_2_5/a_31_74# sky130_fd_sc_hs__and2_2_5/a_118_74#
+ sky130_fd_sc_hs__and2_2
Xsky130_fd_sc_hs__inv_4_72 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_73/Y sky130_fd_sc_hs__inv_4_73/A
+ sky130_fd_sc_hs__inv_4
Xsky130_fd_sc_hs__inv_4_61 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_61/Y sky130_fd_sc_hs__inv_4_61/A
+ sky130_fd_sc_hs__inv_4
Xsky130_fd_sc_hs__inv_4_50 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_51/Y sky130_fd_sc_hs__inv_4_51/A
+ sky130_fd_sc_hs__inv_4
Xsky130_fd_sc_hs__inv_4_94 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_95/Y sky130_fd_sc_hs__inv_4_95/A
+ sky130_fd_sc_hs__inv_4
Xsky130_fd_sc_hs__inv_4_83 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_83/Y sky130_fd_sc_hs__inv_4_83/A
+ sky130_fd_sc_hs__inv_4
Xsky130_fd_sc_hs__a22o_1_19 DVSS DVDD DVDD DVSS osc_fine_con_final[7] manual_control_osc[7]
+ sky130_fd_sc_hs__inv_4_43/Y sky130_fd_sc_hs__fa_2_17/B fftl_en sky130_fd_sc_hs__a22o_1_19/a_222_392#
+ sky130_fd_sc_hs__a22o_1_19/a_230_79# sky130_fd_sc_hs__a22o_1_19/a_52_123# sky130_fd_sc_hs__a22o_1_19/a_132_392#
+ sky130_fd_sc_hs__a22o_1
Xsky130_fd_sc_hs__o21ai_1_6 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__o21ai_1_7/Y sky130_fd_sc_hs__inv_4_91/A
+ sky130_fd_sc_hs__and2_2_5/X sky130_fd_sc_hs__nand2_2_5/B sky130_fd_sc_hs__o21ai_1_7/a_162_368#
+ sky130_fd_sc_hs__o21ai_1_7/a_27_74# sky130_fd_sc_hs__o21ai_1
Xsky130_fd_sc_hs__nand2_1_19 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nor2_1_21/Y sky130_fd_sc_hs__nor2_1_15/B
+ sky130_fd_sc_hs__o21a_1_17/A1 sky130_fd_sc_hs__nand2_1_19/a_117_74# sky130_fd_sc_hs__nand2_1
Xsky130_fd_sc_hs__dfxtp_4_9 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_103/A sky130_fd_sc_hs__nor2_1_89/Y
+ sky130_fd_sc_hs__dfxtp_4_9/CLK sky130_fd_sc_hs__dfxtp_4_9/a_1226_296# sky130_fd_sc_hs__dfxtp_4_9/a_735_102#
+ sky130_fd_sc_hs__dfxtp_4_9/a_1141_508# sky130_fd_sc_hs__dfxtp_4_9/a_206_368# sky130_fd_sc_hs__dfxtp_4_9/a_437_503#
+ sky130_fd_sc_hs__dfxtp_4_9/a_27_74# sky130_fd_sc_hs__dfxtp_4_9/a_651_503# sky130_fd_sc_hs__dfxtp_4_9/a_696_458#
+ sky130_fd_sc_hs__dfxtp_4_9/a_544_485# sky130_fd_sc_hs__dfxtp_4_9/a_1178_124# sky130_fd_sc_hs__dfxtp_4_9/a_1034_424#
+ sky130_fd_sc_hs__dfxtp_4
Xsky130_fd_sc_hs__dfxtp_2_6 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_2_5/B sky130_fd_sc_hs__dfxtp_4_9/CLK
+ sky130_fd_sc_hs__nor2b_2_1/Y sky130_fd_sc_hs__dfxtp_2_7/a_431_508# sky130_fd_sc_hs__dfxtp_2_7/a_1125_508#
+ sky130_fd_sc_hs__dfxtp_2_7/a_206_368# sky130_fd_sc_hs__dfxtp_2_7/a_27_74# sky130_fd_sc_hs__dfxtp_2_7/a_708_101#
+ sky130_fd_sc_hs__dfxtp_2_7/a_1019_424# sky130_fd_sc_hs__dfxtp_2_7/a_1172_124# sky130_fd_sc_hs__dfxtp_2_7/a_644_504#
+ sky130_fd_sc_hs__dfxtp_2_7/a_1217_314# sky130_fd_sc_hs__dfxtp_2_7/a_538_429# sky130_fd_sc_hs__dfxtp_2_7/a_695_459#
+ sky130_fd_sc_hs__dfxtp_2
Xsky130_fd_sc_hs__a21oi_1_108 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__o21a_1_75/A2 sky130_fd_sc_hs__dfrbp_1_31/D
+ sky130_fd_sc_hs__o21a_1_51/B1 sky130_fd_sc_hs__inv_4_107/Y sky130_fd_sc_hs__a21oi_1_109/a_117_74#
+ sky130_fd_sc_hs__a21oi_1_109/a_29_368# sky130_fd_sc_hs__a21oi_1
Xsky130_fd_sc_hs__a21oi_1_119 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__o21a_1_77/A2 sky130_fd_sc_hs__dfrbp_1_37/D
+ sky130_fd_sc_hs__o21a_1_73/B1 sky130_fd_sc_hs__inv_4_115/Y sky130_fd_sc_hs__a21oi_1_119/a_117_74#
+ sky130_fd_sc_hs__a21oi_1_119/a_29_368# sky130_fd_sc_hs__a21oi_1
Xsky130_fd_sc_hs__o31ai_1_0 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__o31ai_1_1/A3 fine_control_avg_window_select[2]
+ sky130_fd_sc_hs__o31ai_1_1/B1 fine_control_avg_window_select[1] sky130_fd_sc_hs__o31ai_1_1/Y
+ sky130_fd_sc_hs__o31ai_1_1/a_114_74# sky130_fd_sc_hs__o31ai_1_1/a_119_368# sky130_fd_sc_hs__o31ai_1_1/a_203_368#
+ sky130_fd_sc_hs__o31ai_1
Xsky130_fd_sc_hs__nand2_1_102 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_133/Y sky130_fd_sc_hs__o211ai_1_9/C1
+ sky130_fd_sc_hs__o21a_1_75/A1 sky130_fd_sc_hs__nand2_1_103/a_117_74# sky130_fd_sc_hs__nand2_1
Xsky130_fd_sc_hs__dfrtn_1_40 DVSS DVDD sky130_fd_sc_hs__clkbuf_8_1/X DVDD DVSS ref_clk
+ sky130_fd_sc_hs__inv_4_129/A sky130_fd_sc_hs__dfrtn_1_41/D sky130_fd_sc_hs__dfrtn_1_41/a_1266_119#
+ sky130_fd_sc_hs__dfrtn_1_41/a_1736_119# sky130_fd_sc_hs__dfrtn_1_41/a_817_508# sky130_fd_sc_hs__dfrtn_1_41/a_120_74#
+ sky130_fd_sc_hs__dfrtn_1_41/a_1547_508# sky130_fd_sc_hs__dfrtn_1_41/a_922_127# sky130_fd_sc_hs__dfrtn_1_41/a_33_74#
+ sky130_fd_sc_hs__dfrtn_1_41/a_714_127# sky130_fd_sc_hs__dfrtn_1_41/a_1934_94# sky130_fd_sc_hs__dfrtn_1_41/a_1550_119#
+ sky130_fd_sc_hs__dfrtn_1_41/a_1598_93# sky130_fd_sc_hs__dfrtn_1_41/a_300_74# sky130_fd_sc_hs__dfrtn_1_41/a_507_368#
+ sky130_fd_sc_hs__dfrtn_1_41/a_856_304# sky130_fd_sc_hs__dfrtn_1_41/a_850_127# sky130_fd_sc_hs__dfrtn_1
Xsky130_fd_sc_hs__nand2_1_113 DVSS DVDD DVDD DVSS div_ratio_half[3] sky130_fd_sc_hs__nand4_2_1/D
+ sky130_fd_sc_hs__inv_2_7/Y sky130_fd_sc_hs__nand2_1_113/a_117_74# sky130_fd_sc_hs__nand2_1
Xsky130_fd_sc_hs__nor2_1_38 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_37/Y sky130_fd_sc_hs__nor4_1_1/C
+ sky130_fd_sc_hs__inv_4_61/A sky130_fd_sc_hs__nor2_1_39/a_116_368# sky130_fd_sc_hs__nor2_1
Xsky130_fd_sc_hs__nor2_1_27 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nor2_1_27/B sky130_fd_sc_hs__nor2_1_27/Y
+ sky130_fd_sc_hs__inv_4_37/Y sky130_fd_sc_hs__nor2_1_27/a_116_368# sky130_fd_sc_hs__nor2_1
Xsky130_fd_sc_hs__nor2_1_16 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__o21a_1_9/B1 sky130_fd_sc_hs__nor2_1_17/Y
+ sky130_fd_sc_hs__inv_4_15/Y sky130_fd_sc_hs__nor2_1_17/a_116_368# sky130_fd_sc_hs__nor2_1
Xsky130_fd_sc_hs__nor2_1_49 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nor2_1_49/B sky130_fd_sc_hs__nor2_1_49/Y
+ sky130_fd_sc_hs__inv_4_59/Y sky130_fd_sc_hs__nor2_1_49/a_116_368# sky130_fd_sc_hs__nor2_1
Xsky130_fd_sc_hs__nor2b_1_38 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nor2_1_65/A sky130_fd_sc_hs__nor3_1_5/B
+ sky130_fd_sc_hs__inv_4_73/A sky130_fd_sc_hs__nor2b_1_39/a_278_368# sky130_fd_sc_hs__nor2b_1_39/a_27_112#
+ sky130_fd_sc_hs__nor2b_1
Xsky130_fd_sc_hs__nor2b_1_27 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__fa_2_19/SUM sky130_fd_sc_hs__nor2b_1_27/Y
+ sky130_fd_sc_hs__or2_1_1/A sky130_fd_sc_hs__nor2b_1_27/a_278_368# sky130_fd_sc_hs__nor2b_1_27/a_27_112#
+ sky130_fd_sc_hs__nor2b_1
Xsky130_fd_sc_hs__nor2b_1_16 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__fa_2_17/SUM sky130_fd_sc_hs__nor2b_1_17/Y
+ sky130_fd_sc_hs__or2_1_1/A sky130_fd_sc_hs__nor2b_1_17/a_278_368# sky130_fd_sc_hs__nor2b_1_17/a_27_112#
+ sky130_fd_sc_hs__nor2b_1
Xsky130_fd_sc_hs__nor2b_1_49 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__o21a_1_71/A1 sky130_fd_sc_hs__nor3_1_13/A
+ sky130_fd_sc_hs__inv_4_113/A sky130_fd_sc_hs__nor2b_1_49/a_278_368# sky130_fd_sc_hs__nor2b_1_49/a_27_112#
+ sky130_fd_sc_hs__nor2b_1
Xsky130_fd_sc_hs__inv_4_108 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_109/Y sky130_fd_sc_hs__inv_4_109/A
+ sky130_fd_sc_hs__inv_4
Xsky130_fd_sc_hs__inv_4_119 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_87/A sky130_fd_sc_hs__nand4_2_1/Y
+ sky130_fd_sc_hs__inv_4
Xsky130_fd_sc_hs__o22ai_1_8 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__maj3_1_1/X sky130_fd_sc_hs__o22ai_1_9/B1
+ sky130_fd_sc_hs__o22ai_1_9/Y sky130_fd_sc_hs__inv_4_109/Y sky130_fd_sc_hs__o22ai_1_9/A1
+ sky130_fd_sc_hs__o22ai_1_9/a_340_368# sky130_fd_sc_hs__o22ai_1_9/a_142_368# sky130_fd_sc_hs__o22ai_1_9/a_27_74#
+ sky130_fd_sc_hs__o22ai_1
Xsky130_fd_sc_hs__dfstp_2_0 DVSS DVDD sky130_fd_sc_hs__inv_4_49/Y DVDD DVSS sky130_fd_sc_hs__dfstp_2_1/CLK
+ sky130_fd_sc_hs__or2_1_1/X sky130_fd_sc_hs__xor2_1_9/A sky130_fd_sc_hs__dfstp_2_1/a_1566_92#
+ sky130_fd_sc_hs__dfstp_2_1/a_1521_508# sky130_fd_sc_hs__dfstp_2_1/a_716_456# sky130_fd_sc_hs__dfstp_2_1/a_1266_341#
+ sky130_fd_sc_hs__dfstp_2_1/a_1278_74# sky130_fd_sc_hs__dfstp_2_1/a_398_74# sky130_fd_sc_hs__dfstp_2_1/a_1057_118#
+ sky130_fd_sc_hs__dfstp_2_1/a_1489_118# sky130_fd_sc_hs__dfstp_2_1/a_27_74# sky130_fd_sc_hs__dfstp_2_1/a_1596_118#
+ sky130_fd_sc_hs__dfstp_2_1/a_225_74# sky130_fd_sc_hs__dfstp_2_1/a_1356_74# sky130_fd_sc_hs__dfstp_2_1/a_612_74#
+ sky130_fd_sc_hs__dfstp_2_1/a_781_74# sky130_fd_sc_hs__dfstp_2_1/a_767_384# sky130_fd_sc_hs__dfstp_2_1/a_2022_94#
+ sky130_fd_sc_hs__dfstp_2
Xsky130_fd_sc_hs__dfrtp_4_2 DVSS DVDD sky130_fd_sc_hs__clkbuf_8_1/A DVDD DVSS sky130_fd_sc_hs__dfrtp_4_3/D
+ sky130_fd_sc_hs__nand2_1_47/B sky130_fd_sc_hs__inv_4_3/A sky130_fd_sc_hs__dfrtp_4_3/a_37_78#
+ sky130_fd_sc_hs__dfrtp_4_3/a_494_366# sky130_fd_sc_hs__dfrtp_4_3/a_699_463# sky130_fd_sc_hs__dfrtp_4_3/a_313_74#
+ sky130_fd_sc_hs__dfrtp_4_3/a_1627_493# sky130_fd_sc_hs__dfrtp_4_3/a_1678_395# sky130_fd_sc_hs__dfrtp_4_3/a_1827_81#
+ sky130_fd_sc_hs__dfrtp_4_3/a_789_463# sky130_fd_sc_hs__dfrtp_4_3/a_1350_392# sky130_fd_sc_hs__dfrtp_4_3/a_834_355#
+ sky130_fd_sc_hs__dfrtp_4_3/a_812_138# sky130_fd_sc_hs__dfrtp_4_3/a_124_78# sky130_fd_sc_hs__dfrtp_4_3/a_1647_81#
+ sky130_fd_sc_hs__dfrtp_4_3/a_2010_409# sky130_fd_sc_hs__dfrtp_4_3/a_890_138# sky130_fd_sc_hs__dfrtp_4
Xsky130_fd_sc_hs__inv_4_62 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_63/Y sky130_fd_sc_hs__inv_4_63/A
+ sky130_fd_sc_hs__inv_4
Xsky130_fd_sc_hs__inv_4_51 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_51/Y sky130_fd_sc_hs__inv_4_51/A
+ sky130_fd_sc_hs__inv_4
Xsky130_fd_sc_hs__inv_4_40 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_41/Y sky130_fd_sc_hs__inv_4_41/A
+ sky130_fd_sc_hs__inv_4
Xsky130_fd_sc_hs__inv_4_95 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_95/Y sky130_fd_sc_hs__inv_4_95/A
+ sky130_fd_sc_hs__inv_4
Xsky130_fd_sc_hs__inv_4_84 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_85/Y sky130_fd_sc_hs__inv_4_85/A
+ sky130_fd_sc_hs__inv_4
Xsky130_fd_sc_hs__inv_4_73 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_73/Y sky130_fd_sc_hs__inv_4_73/A
+ sky130_fd_sc_hs__inv_4
Xsky130_fd_sc_hs__o21ai_1_7 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__o21ai_1_7/Y sky130_fd_sc_hs__inv_4_91/A
+ sky130_fd_sc_hs__and2_2_5/X sky130_fd_sc_hs__nand2_2_5/B sky130_fd_sc_hs__o21ai_1_7/a_162_368#
+ sky130_fd_sc_hs__o21ai_1_7/a_27_74# sky130_fd_sc_hs__o21ai_1
Xsky130_fd_sc_hs__dfrbp_1_40 DVSS DVDD sky130_fd_sc_hs__clkbuf_8_1/X DVDD DVSS sky130_fd_sc_hs__inv_4_135/A
+ ref_clk sky130_fd_sc_hs__dfrbp_1_41/D sky130_fd_sc_hs__dfrbp_1_41/Q_N sky130_fd_sc_hs__dfrbp_1_41/a_498_360#
+ sky130_fd_sc_hs__dfrbp_1_41/a_1224_74# sky130_fd_sc_hs__dfrbp_1_41/a_2026_424# sky130_fd_sc_hs__dfrbp_1_41/a_1482_48#
+ sky130_fd_sc_hs__dfrbp_1_41/a_125_78# sky130_fd_sc_hs__dfrbp_1_41/a_796_463# sky130_fd_sc_hs__dfrbp_1_41/a_910_118#
+ sky130_fd_sc_hs__dfrbp_1_41/a_1465_471# sky130_fd_sc_hs__dfrbp_1_41/a_832_118# sky130_fd_sc_hs__dfrbp_1_41/a_841_401#
+ sky130_fd_sc_hs__dfrbp_1_41/a_38_78# sky130_fd_sc_hs__dfrbp_1_41/a_1434_74# sky130_fd_sc_hs__dfrbp_1_41/a_706_463#
+ sky130_fd_sc_hs__dfrbp_1_41/a_319_360# sky130_fd_sc_hs__dfrbp_1_41/a_1624_74# sky130_fd_sc_hs__dfrbp_1
Xsky130_fd_sc_hs__dfxtp_2_7 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_2_5/B sky130_fd_sc_hs__dfxtp_4_9/CLK
+ sky130_fd_sc_hs__nor2b_2_1/Y sky130_fd_sc_hs__dfxtp_2_7/a_431_508# sky130_fd_sc_hs__dfxtp_2_7/a_1125_508#
+ sky130_fd_sc_hs__dfxtp_2_7/a_206_368# sky130_fd_sc_hs__dfxtp_2_7/a_27_74# sky130_fd_sc_hs__dfxtp_2_7/a_708_101#
+ sky130_fd_sc_hs__dfxtp_2_7/a_1019_424# sky130_fd_sc_hs__dfxtp_2_7/a_1172_124# sky130_fd_sc_hs__dfxtp_2_7/a_644_504#
+ sky130_fd_sc_hs__dfxtp_2_7/a_1217_314# sky130_fd_sc_hs__dfxtp_2_7/a_538_429# sky130_fd_sc_hs__dfxtp_2_7/a_695_459#
+ sky130_fd_sc_hs__dfxtp_2
Xsky130_fd_sc_hs__a21oi_1_109 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__o21a_1_75/A2 sky130_fd_sc_hs__dfrbp_1_31/D
+ sky130_fd_sc_hs__o21a_1_51/B1 sky130_fd_sc_hs__inv_4_107/Y sky130_fd_sc_hs__a21oi_1_109/a_117_74#
+ sky130_fd_sc_hs__a21oi_1_109/a_29_368# sky130_fd_sc_hs__a21oi_1
Xsky130_fd_sc_hs__o31ai_1_1 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__o31ai_1_1/A3 fine_control_avg_window_select[2]
+ sky130_fd_sc_hs__o31ai_1_1/B1 fine_control_avg_window_select[1] sky130_fd_sc_hs__o31ai_1_1/Y
+ sky130_fd_sc_hs__o31ai_1_1/a_114_74# sky130_fd_sc_hs__o31ai_1_1/a_119_368# sky130_fd_sc_hs__o31ai_1_1/a_203_368#
+ sky130_fd_sc_hs__o31ai_1
Xsky130_fd_sc_hs__dfrtn_1_30 DVSS DVDD sky130_fd_sc_hs__clkbuf_8_1/X DVDD DVSS ref_clk
+ sky130_fd_sc_hs__inv_4_99/A sky130_fd_sc_hs__dfrtn_1_31/D sky130_fd_sc_hs__dfrtn_1_31/a_1266_119#
+ sky130_fd_sc_hs__dfrtn_1_31/a_1736_119# sky130_fd_sc_hs__dfrtn_1_31/a_817_508# sky130_fd_sc_hs__dfrtn_1_31/a_120_74#
+ sky130_fd_sc_hs__dfrtn_1_31/a_1547_508# sky130_fd_sc_hs__dfrtn_1_31/a_922_127# sky130_fd_sc_hs__dfrtn_1_31/a_33_74#
+ sky130_fd_sc_hs__dfrtn_1_31/a_714_127# sky130_fd_sc_hs__dfrtn_1_31/a_1934_94# sky130_fd_sc_hs__dfrtn_1_31/a_1550_119#
+ sky130_fd_sc_hs__dfrtn_1_31/a_1598_93# sky130_fd_sc_hs__dfrtn_1_31/a_300_74# sky130_fd_sc_hs__dfrtn_1_31/a_507_368#
+ sky130_fd_sc_hs__dfrtn_1_31/a_856_304# sky130_fd_sc_hs__dfrtn_1_31/a_850_127# sky130_fd_sc_hs__dfrtn_1
Xsky130_fd_sc_hs__nand2_1_103 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_133/Y sky130_fd_sc_hs__o211ai_1_9/C1
+ sky130_fd_sc_hs__o21a_1_75/A1 sky130_fd_sc_hs__nand2_1_103/a_117_74# sky130_fd_sc_hs__nand2_1
Xsky130_fd_sc_hs__dfrtn_1_41 DVSS DVDD sky130_fd_sc_hs__clkbuf_8_1/X DVDD DVSS ref_clk
+ sky130_fd_sc_hs__inv_4_129/A sky130_fd_sc_hs__dfrtn_1_41/D sky130_fd_sc_hs__dfrtn_1_41/a_1266_119#
+ sky130_fd_sc_hs__dfrtn_1_41/a_1736_119# sky130_fd_sc_hs__dfrtn_1_41/a_817_508# sky130_fd_sc_hs__dfrtn_1_41/a_120_74#
+ sky130_fd_sc_hs__dfrtn_1_41/a_1547_508# sky130_fd_sc_hs__dfrtn_1_41/a_922_127# sky130_fd_sc_hs__dfrtn_1_41/a_33_74#
+ sky130_fd_sc_hs__dfrtn_1_41/a_714_127# sky130_fd_sc_hs__dfrtn_1_41/a_1934_94# sky130_fd_sc_hs__dfrtn_1_41/a_1550_119#
+ sky130_fd_sc_hs__dfrtn_1_41/a_1598_93# sky130_fd_sc_hs__dfrtn_1_41/a_300_74# sky130_fd_sc_hs__dfrtn_1_41/a_507_368#
+ sky130_fd_sc_hs__dfrtn_1_41/a_856_304# sky130_fd_sc_hs__dfrtn_1_41/a_850_127# sky130_fd_sc_hs__dfrtn_1
Xsky130_fd_sc_hs__nand2_1_114 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__o21a_1_73/A2 sky130_fd_sc_hs__o21a_1_73/B1
+ sky130_fd_sc_hs__or2_1_3/A sky130_fd_sc_hs__nand2_1_115/a_117_74# sky130_fd_sc_hs__nand2_1
Xsky130_fd_sc_hs__a222o_1_0 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nor2b_1_23/Y sky130_fd_sc_hs__a222o_1_1/X
+ sky130_fd_sc_hs__inv_4_29/A sky130_fd_sc_hs__nor2b_1_25/Y sky130_fd_sc_hs__and2_2_1/X
+ sky130_fd_sc_hs__inv_4_35/A sky130_fd_sc_hs__inv_4_31/A sky130_fd_sc_hs__a222o_1_1/a_27_390#
+ sky130_fd_sc_hs__a222o_1_1/a_386_74# sky130_fd_sc_hs__a222o_1_1/a_119_74# sky130_fd_sc_hs__a222o_1_1/a_651_74#
+ sky130_fd_sc_hs__a222o_1_1/a_32_74# sky130_fd_sc_hs__a222o_1_1/a_337_390# sky130_fd_sc_hs__a222o_1
Xsky130_fd_sc_hs__nor2_1_28 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nor2_1_29/B sky130_fd_sc_hs__nor2_1_29/Y
+ sky130_fd_sc_hs__inv_4_53/Y sky130_fd_sc_hs__nor2_1_29/a_116_368# sky130_fd_sc_hs__nor2_1
Xsky130_fd_sc_hs__nor2_1_17 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__o21a_1_9/B1 sky130_fd_sc_hs__nor2_1_17/Y
+ sky130_fd_sc_hs__inv_4_15/Y sky130_fd_sc_hs__nor2_1_17/a_116_368# sky130_fd_sc_hs__nor2_1
Xsky130_fd_sc_hs__nor2_1_39 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_37/Y sky130_fd_sc_hs__nor4_1_1/C
+ sky130_fd_sc_hs__inv_4_61/A sky130_fd_sc_hs__nor2_1_39/a_116_368# sky130_fd_sc_hs__nor2_1
Xsky130_fd_sc_hs__nor2b_1_28 DVSS DVDD DVDD DVSS aux_clk_out sky130_fd_sc_hs__nor2b_1_29/Y
+ sky130_fd_sc_hs__nor2b_1_33/Y sky130_fd_sc_hs__nor2b_1_29/a_278_368# sky130_fd_sc_hs__nor2b_1_29/a_27_112#
+ sky130_fd_sc_hs__nor2b_1
Xsky130_fd_sc_hs__nor2b_1_17 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__fa_2_17/SUM sky130_fd_sc_hs__nor2b_1_17/Y
+ sky130_fd_sc_hs__or2_1_1/A sky130_fd_sc_hs__nor2b_1_17/a_278_368# sky130_fd_sc_hs__nor2b_1_17/a_27_112#
+ sky130_fd_sc_hs__nor2b_1
Xsky130_fd_sc_hs__nor2b_1_39 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nor2_1_65/A sky130_fd_sc_hs__nor3_1_5/B
+ sky130_fd_sc_hs__inv_4_73/A sky130_fd_sc_hs__nor2b_1_39/a_278_368# sky130_fd_sc_hs__nor2b_1_39/a_27_112#
+ sky130_fd_sc_hs__nor2b_1
Xsky130_fd_sc_hs__inv_4_109 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_109/Y sky130_fd_sc_hs__inv_4_109/A
+ sky130_fd_sc_hs__inv_4
Xsky130_fd_sc_hs__o22ai_1_9 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__maj3_1_1/X sky130_fd_sc_hs__o22ai_1_9/B1
+ sky130_fd_sc_hs__o22ai_1_9/Y sky130_fd_sc_hs__inv_4_109/Y sky130_fd_sc_hs__o22ai_1_9/A1
+ sky130_fd_sc_hs__o22ai_1_9/a_340_368# sky130_fd_sc_hs__o22ai_1_9/a_142_368# sky130_fd_sc_hs__o22ai_1_9/a_27_74#
+ sky130_fd_sc_hs__o22ai_1
Xsky130_fd_sc_hs__dfstp_2_1 DVSS DVDD sky130_fd_sc_hs__inv_4_49/Y DVDD DVSS sky130_fd_sc_hs__dfstp_2_1/CLK
+ sky130_fd_sc_hs__or2_1_1/X sky130_fd_sc_hs__xor2_1_9/A sky130_fd_sc_hs__dfstp_2_1/a_1566_92#
+ sky130_fd_sc_hs__dfstp_2_1/a_1521_508# sky130_fd_sc_hs__dfstp_2_1/a_716_456# sky130_fd_sc_hs__dfstp_2_1/a_1266_341#
+ sky130_fd_sc_hs__dfstp_2_1/a_1278_74# sky130_fd_sc_hs__dfstp_2_1/a_398_74# sky130_fd_sc_hs__dfstp_2_1/a_1057_118#
+ sky130_fd_sc_hs__dfstp_2_1/a_1489_118# sky130_fd_sc_hs__dfstp_2_1/a_27_74# sky130_fd_sc_hs__dfstp_2_1/a_1596_118#
+ sky130_fd_sc_hs__dfstp_2_1/a_225_74# sky130_fd_sc_hs__dfstp_2_1/a_1356_74# sky130_fd_sc_hs__dfstp_2_1/a_612_74#
+ sky130_fd_sc_hs__dfstp_2_1/a_781_74# sky130_fd_sc_hs__dfstp_2_1/a_767_384# sky130_fd_sc_hs__dfstp_2_1/a_2022_94#
+ sky130_fd_sc_hs__dfstp_2
Xsky130_fd_sc_hs__dfrtp_4_3 DVSS DVDD sky130_fd_sc_hs__clkbuf_8_1/A DVDD DVSS sky130_fd_sc_hs__dfrtp_4_3/D
+ sky130_fd_sc_hs__nand2_1_47/B sky130_fd_sc_hs__inv_4_3/A sky130_fd_sc_hs__dfrtp_4_3/a_37_78#
+ sky130_fd_sc_hs__dfrtp_4_3/a_494_366# sky130_fd_sc_hs__dfrtp_4_3/a_699_463# sky130_fd_sc_hs__dfrtp_4_3/a_313_74#
+ sky130_fd_sc_hs__dfrtp_4_3/a_1627_493# sky130_fd_sc_hs__dfrtp_4_3/a_1678_395# sky130_fd_sc_hs__dfrtp_4_3/a_1827_81#
+ sky130_fd_sc_hs__dfrtp_4_3/a_789_463# sky130_fd_sc_hs__dfrtp_4_3/a_1350_392# sky130_fd_sc_hs__dfrtp_4_3/a_834_355#
+ sky130_fd_sc_hs__dfrtp_4_3/a_812_138# sky130_fd_sc_hs__dfrtp_4_3/a_124_78# sky130_fd_sc_hs__dfrtp_4_3/a_1647_81#
+ sky130_fd_sc_hs__dfrtp_4_3/a_2010_409# sky130_fd_sc_hs__dfrtp_4_3/a_890_138# sky130_fd_sc_hs__dfrtp_4
Xsky130_fd_sc_hs__inv_4_63 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_63/Y sky130_fd_sc_hs__inv_4_63/A
+ sky130_fd_sc_hs__inv_4
Xsky130_fd_sc_hs__inv_4_52 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_53/Y sky130_fd_sc_hs__inv_4_53/A
+ sky130_fd_sc_hs__inv_4
Xsky130_fd_sc_hs__inv_4_41 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_41/Y sky130_fd_sc_hs__inv_4_41/A
+ sky130_fd_sc_hs__inv_4
Xsky130_fd_sc_hs__inv_4_30 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_31/Y sky130_fd_sc_hs__inv_4_31/A
+ sky130_fd_sc_hs__inv_4
Xsky130_fd_sc_hs__inv_4_96 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_97/Y sky130_fd_sc_hs__inv_4_97/A
+ sky130_fd_sc_hs__inv_4
Xsky130_fd_sc_hs__inv_4_85 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_85/Y sky130_fd_sc_hs__inv_4_85/A
+ sky130_fd_sc_hs__inv_4
Xsky130_fd_sc_hs__inv_4_74 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_75/Y sky130_fd_sc_hs__inv_4_75/A
+ sky130_fd_sc_hs__inv_4
Xsky130_fd_sc_hs__o21ai_1_8 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__o21ai_1_9/Y sky130_fd_sc_hs__nand2_2_7/Y
+ sky130_fd_sc_hs__nand2_2_7/B sky130_fd_sc_hs__inv_2_9/A sky130_fd_sc_hs__o21ai_1_9/a_162_368#
+ sky130_fd_sc_hs__o21ai_1_9/a_27_74# sky130_fd_sc_hs__o21ai_1
Xsky130_fd_sc_hs__nor3_1_0 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nor3_1_1/Y sky130_fd_sc_hs__nor3_1_1/C
+ sky130_fd_sc_hs__nor3_1_1/B sky130_fd_sc_hs__nor3_1_1/A sky130_fd_sc_hs__nor3_1_1/a_198_368#
+ sky130_fd_sc_hs__nor3_1_1/a_114_368# sky130_fd_sc_hs__nor3_1
Xsky130_fd_sc_hs__a22oi_1_0 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nor2_1_33/Y sky130_fd_sc_hs__a22oi_1_1/Y
+ sky130_fd_sc_hs__inv_4_3/A sky130_fd_sc_hs__and2_2_1/X sky130_fd_sc_hs__inv_4_9/A
+ sky130_fd_sc_hs__a22oi_1_1/a_71_368# sky130_fd_sc_hs__a22oi_1_1/a_159_74# sky130_fd_sc_hs__a22oi_1_1/a_339_74#
+ sky130_fd_sc_hs__a22oi_1
Xsky130_fd_sc_hs__dfrbp_1_30 DVSS DVDD sky130_fd_sc_hs__clkbuf_8_1/X DVDD DVSS sky130_fd_sc_hs__nor2_1_95/A
+ ref_clk sky130_fd_sc_hs__dfrbp_1_31/D sky130_fd_sc_hs__dfrbp_1_31/Q_N sky130_fd_sc_hs__dfrbp_1_31/a_498_360#
+ sky130_fd_sc_hs__dfrbp_1_31/a_1224_74# sky130_fd_sc_hs__dfrbp_1_31/a_2026_424# sky130_fd_sc_hs__dfrbp_1_31/a_1482_48#
+ sky130_fd_sc_hs__dfrbp_1_31/a_125_78# sky130_fd_sc_hs__dfrbp_1_31/a_796_463# sky130_fd_sc_hs__dfrbp_1_31/a_910_118#
+ sky130_fd_sc_hs__dfrbp_1_31/a_1465_471# sky130_fd_sc_hs__dfrbp_1_31/a_832_118# sky130_fd_sc_hs__dfrbp_1_31/a_841_401#
+ sky130_fd_sc_hs__dfrbp_1_31/a_38_78# sky130_fd_sc_hs__dfrbp_1_31/a_1434_74# sky130_fd_sc_hs__dfrbp_1_31/a_706_463#
+ sky130_fd_sc_hs__dfrbp_1_31/a_319_360# sky130_fd_sc_hs__dfrbp_1_31/a_1624_74# sky130_fd_sc_hs__dfrbp_1
Xsky130_fd_sc_hs__dfrbp_1_41 DVSS DVDD sky130_fd_sc_hs__clkbuf_8_1/X DVDD DVSS sky130_fd_sc_hs__inv_4_135/A
+ ref_clk sky130_fd_sc_hs__dfrbp_1_41/D sky130_fd_sc_hs__dfrbp_1_41/Q_N sky130_fd_sc_hs__dfrbp_1_41/a_498_360#
+ sky130_fd_sc_hs__dfrbp_1_41/a_1224_74# sky130_fd_sc_hs__dfrbp_1_41/a_2026_424# sky130_fd_sc_hs__dfrbp_1_41/a_1482_48#
+ sky130_fd_sc_hs__dfrbp_1_41/a_125_78# sky130_fd_sc_hs__dfrbp_1_41/a_796_463# sky130_fd_sc_hs__dfrbp_1_41/a_910_118#
+ sky130_fd_sc_hs__dfrbp_1_41/a_1465_471# sky130_fd_sc_hs__dfrbp_1_41/a_832_118# sky130_fd_sc_hs__dfrbp_1_41/a_841_401#
+ sky130_fd_sc_hs__dfrbp_1_41/a_38_78# sky130_fd_sc_hs__dfrbp_1_41/a_1434_74# sky130_fd_sc_hs__dfrbp_1_41/a_706_463#
+ sky130_fd_sc_hs__dfrbp_1_41/a_319_360# sky130_fd_sc_hs__dfrbp_1_41/a_1624_74# sky130_fd_sc_hs__dfrbp_1
Xsky130_fd_sc_hs__dfxtp_2_8 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_2_5/A sky130_fd_sc_hs__dfxtp_4_9/CLK
+ sky130_fd_sc_hs__nor2_1_77/Y sky130_fd_sc_hs__dfxtp_2_9/a_431_508# sky130_fd_sc_hs__dfxtp_2_9/a_1125_508#
+ sky130_fd_sc_hs__dfxtp_2_9/a_206_368# sky130_fd_sc_hs__dfxtp_2_9/a_27_74# sky130_fd_sc_hs__dfxtp_2_9/a_708_101#
+ sky130_fd_sc_hs__dfxtp_2_9/a_1019_424# sky130_fd_sc_hs__dfxtp_2_9/a_1172_124# sky130_fd_sc_hs__dfxtp_2_9/a_644_504#
+ sky130_fd_sc_hs__dfxtp_2_9/a_1217_314# sky130_fd_sc_hs__dfxtp_2_9/a_538_429# sky130_fd_sc_hs__dfxtp_2_9/a_695_459#
+ sky130_fd_sc_hs__dfxtp_2
Xsky130_fd_sc_hs__o31ai_1_2 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_63/Y sky130_fd_sc_hs__nor2_1_65/Y
+ sky130_fd_sc_hs__o31ai_1_3/B1 sky130_fd_sc_hs__inv_4_67/A sky130_fd_sc_hs__o31ai_1_3/Y
+ sky130_fd_sc_hs__o31ai_1_3/a_114_74# sky130_fd_sc_hs__o31ai_1_3/a_119_368# sky130_fd_sc_hs__o31ai_1_3/a_203_368#
+ sky130_fd_sc_hs__o31ai_1
Xsky130_fd_sc_hs__dfrtn_1_20 DVSS DVDD sky130_fd_sc_hs__clkbuf_8_1/X DVDD DVSS sky130_fd_sc_hs__clkbuf_2_1/X
+ sky130_fd_sc_hs__inv_4_83/A sky130_fd_sc_hs__o21a_1_49/X sky130_fd_sc_hs__dfrtn_1_21/a_1266_119#
+ sky130_fd_sc_hs__dfrtn_1_21/a_1736_119# sky130_fd_sc_hs__dfrtn_1_21/a_817_508# sky130_fd_sc_hs__dfrtn_1_21/a_120_74#
+ sky130_fd_sc_hs__dfrtn_1_21/a_1547_508# sky130_fd_sc_hs__dfrtn_1_21/a_922_127# sky130_fd_sc_hs__dfrtn_1_21/a_33_74#
+ sky130_fd_sc_hs__dfrtn_1_21/a_714_127# sky130_fd_sc_hs__dfrtn_1_21/a_1934_94# sky130_fd_sc_hs__dfrtn_1_21/a_1550_119#
+ sky130_fd_sc_hs__dfrtn_1_21/a_1598_93# sky130_fd_sc_hs__dfrtn_1_21/a_300_74# sky130_fd_sc_hs__dfrtn_1_21/a_507_368#
+ sky130_fd_sc_hs__dfrtn_1_21/a_856_304# sky130_fd_sc_hs__dfrtn_1_21/a_850_127# sky130_fd_sc_hs__dfrtn_1
Xsky130_fd_sc_hs__dfrtn_1_31 DVSS DVDD sky130_fd_sc_hs__clkbuf_8_1/X DVDD DVSS ref_clk
+ sky130_fd_sc_hs__inv_4_99/A sky130_fd_sc_hs__dfrtn_1_31/D sky130_fd_sc_hs__dfrtn_1_31/a_1266_119#
+ sky130_fd_sc_hs__dfrtn_1_31/a_1736_119# sky130_fd_sc_hs__dfrtn_1_31/a_817_508# sky130_fd_sc_hs__dfrtn_1_31/a_120_74#
+ sky130_fd_sc_hs__dfrtn_1_31/a_1547_508# sky130_fd_sc_hs__dfrtn_1_31/a_922_127# sky130_fd_sc_hs__dfrtn_1_31/a_33_74#
+ sky130_fd_sc_hs__dfrtn_1_31/a_714_127# sky130_fd_sc_hs__dfrtn_1_31/a_1934_94# sky130_fd_sc_hs__dfrtn_1_31/a_1550_119#
+ sky130_fd_sc_hs__dfrtn_1_31/a_1598_93# sky130_fd_sc_hs__dfrtn_1_31/a_300_74# sky130_fd_sc_hs__dfrtn_1_31/a_507_368#
+ sky130_fd_sc_hs__dfrtn_1_31/a_856_304# sky130_fd_sc_hs__dfrtn_1_31/a_850_127# sky130_fd_sc_hs__dfrtn_1
Xsky130_fd_sc_hs__nand2_1_104 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_135/Y sky130_fd_sc_hs__maj3_1_3/C
+ sky130_fd_sc_hs__inv_4_125/A sky130_fd_sc_hs__nand2_1_105/a_117_74# sky130_fd_sc_hs__nand2_1
Xsky130_fd_sc_hs__dfrtn_1_42 DVSS DVDD sky130_fd_sc_hs__clkbuf_8_1/X DVDD DVSS ref_clk
+ sky130_fd_sc_hs__inv_4_101/A sky130_fd_sc_hs__o21a_1_65/X sky130_fd_sc_hs__dfrtn_1_43/a_1266_119#
+ sky130_fd_sc_hs__dfrtn_1_43/a_1736_119# sky130_fd_sc_hs__dfrtn_1_43/a_817_508# sky130_fd_sc_hs__dfrtn_1_43/a_120_74#
+ sky130_fd_sc_hs__dfrtn_1_43/a_1547_508# sky130_fd_sc_hs__dfrtn_1_43/a_922_127# sky130_fd_sc_hs__dfrtn_1_43/a_33_74#
+ sky130_fd_sc_hs__dfrtn_1_43/a_714_127# sky130_fd_sc_hs__dfrtn_1_43/a_1934_94# sky130_fd_sc_hs__dfrtn_1_43/a_1550_119#
+ sky130_fd_sc_hs__dfrtn_1_43/a_1598_93# sky130_fd_sc_hs__dfrtn_1_43/a_300_74# sky130_fd_sc_hs__dfrtn_1_43/a_507_368#
+ sky130_fd_sc_hs__dfrtn_1_43/a_856_304# sky130_fd_sc_hs__dfrtn_1_43/a_850_127# sky130_fd_sc_hs__dfrtn_1
Xsky130_fd_sc_hs__nand2_1_115 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__o21a_1_73/A2 sky130_fd_sc_hs__o21a_1_73/B1
+ sky130_fd_sc_hs__or2_1_3/A sky130_fd_sc_hs__nand2_1_115/a_117_74# sky130_fd_sc_hs__nand2_1
Xsky130_fd_sc_hs__a222o_1_1 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nor2b_1_23/Y sky130_fd_sc_hs__a222o_1_1/X
+ sky130_fd_sc_hs__inv_4_29/A sky130_fd_sc_hs__nor2b_1_25/Y sky130_fd_sc_hs__and2_2_1/X
+ sky130_fd_sc_hs__inv_4_35/A sky130_fd_sc_hs__inv_4_31/A sky130_fd_sc_hs__a222o_1_1/a_27_390#
+ sky130_fd_sc_hs__a222o_1_1/a_386_74# sky130_fd_sc_hs__a222o_1_1/a_119_74# sky130_fd_sc_hs__a222o_1_1/a_651_74#
+ sky130_fd_sc_hs__a222o_1_1/a_32_74# sky130_fd_sc_hs__a222o_1_1/a_337_390# sky130_fd_sc_hs__a222o_1
Xsky130_fd_sc_hs__nor2_1_29 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nor2_1_29/B sky130_fd_sc_hs__nor2_1_29/Y
+ sky130_fd_sc_hs__inv_4_53/Y sky130_fd_sc_hs__nor2_1_29/a_116_368# sky130_fd_sc_hs__nor2_1
Xsky130_fd_sc_hs__nor2_1_18 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nor2_1_19/B sky130_fd_sc_hs__o21a_1_7/A2
+ sky130_fd_sc_hs__inv_4_29/Y sky130_fd_sc_hs__nor2_1_19/a_116_368# sky130_fd_sc_hs__nor2_1
Xsky130_fd_sc_hs__nor2b_1_29 DVSS DVDD DVDD DVSS aux_clk_out sky130_fd_sc_hs__nor2b_1_29/Y
+ sky130_fd_sc_hs__nor2b_1_33/Y sky130_fd_sc_hs__nor2b_1_29/a_278_368# sky130_fd_sc_hs__nor2b_1_29/a_27_112#
+ sky130_fd_sc_hs__nor2b_1
Xsky130_fd_sc_hs__nor2b_1_18 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__fa_2_21/SUM sky130_fd_sc_hs__nor2b_1_19/Y
+ sky130_fd_sc_hs__or2_1_1/A sky130_fd_sc_hs__nor2b_1_19/a_278_368# sky130_fd_sc_hs__nor2b_1_19/a_27_112#
+ sky130_fd_sc_hs__nor2b_1
Xsky130_fd_sc_hs__dfstp_2_2 DVSS DVDD sky130_fd_sc_hs__inv_4_49/Y DVDD DVSS sky130_fd_sc_hs__o21ai_1_1/Y
+ sky130_fd_sc_hs__nor3_1_3/Y sky130_fd_sc_hs__dfstp_2_5/D sky130_fd_sc_hs__dfstp_2_4/a_1566_92#
+ sky130_fd_sc_hs__dfstp_2_4/a_1521_508# sky130_fd_sc_hs__dfstp_2_4/a_716_456# sky130_fd_sc_hs__dfstp_2_4/a_1266_341#
+ sky130_fd_sc_hs__dfstp_2_4/a_1278_74# sky130_fd_sc_hs__dfstp_2_4/a_398_74# sky130_fd_sc_hs__dfstp_2_4/a_1057_118#
+ sky130_fd_sc_hs__dfstp_2_4/a_1489_118# sky130_fd_sc_hs__dfstp_2_4/a_27_74# sky130_fd_sc_hs__dfstp_2_4/a_1596_118#
+ sky130_fd_sc_hs__dfstp_2_4/a_225_74# sky130_fd_sc_hs__dfstp_2_4/a_1356_74# sky130_fd_sc_hs__dfstp_2_4/a_612_74#
+ sky130_fd_sc_hs__dfstp_2_4/a_781_74# sky130_fd_sc_hs__dfstp_2_4/a_767_384# sky130_fd_sc_hs__dfstp_2_4/a_2022_94#
+ sky130_fd_sc_hs__dfstp_2
Xsky130_fd_sc_hs__dfrtp_4_4 DVSS DVDD sky130_fd_sc_hs__clkbuf_8_1/X DVDD DVSS sky130_fd_sc_hs__dfrtp_4_5/D
+ sky130_fd_sc_hs__nand2_1_47/B sky130_fd_sc_hs__inv_4_7/A sky130_fd_sc_hs__dfrtp_4_5/a_37_78#
+ sky130_fd_sc_hs__dfrtp_4_5/a_494_366# sky130_fd_sc_hs__dfrtp_4_5/a_699_463# sky130_fd_sc_hs__dfrtp_4_5/a_313_74#
+ sky130_fd_sc_hs__dfrtp_4_5/a_1627_493# sky130_fd_sc_hs__dfrtp_4_5/a_1678_395# sky130_fd_sc_hs__dfrtp_4_5/a_1827_81#
+ sky130_fd_sc_hs__dfrtp_4_5/a_789_463# sky130_fd_sc_hs__dfrtp_4_5/a_1350_392# sky130_fd_sc_hs__dfrtp_4_5/a_834_355#
+ sky130_fd_sc_hs__dfrtp_4_5/a_812_138# sky130_fd_sc_hs__dfrtp_4_5/a_124_78# sky130_fd_sc_hs__dfrtp_4_5/a_1647_81#
+ sky130_fd_sc_hs__dfrtp_4_5/a_2010_409# sky130_fd_sc_hs__dfrtp_4_5/a_890_138# sky130_fd_sc_hs__dfrtp_4
Xsky130_fd_sc_hs__inv_4_20 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_21/Y fine_control_avg_window_select[1]
+ sky130_fd_sc_hs__inv_4
Xsky130_fd_sc_hs__inv_4_53 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_53/Y sky130_fd_sc_hs__inv_4_53/A
+ sky130_fd_sc_hs__inv_4
Xsky130_fd_sc_hs__inv_4_42 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_43/Y fftl_en
+ sky130_fd_sc_hs__inv_4
Xsky130_fd_sc_hs__inv_4_31 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_31/Y sky130_fd_sc_hs__inv_4_31/A
+ sky130_fd_sc_hs__inv_4
Xsky130_fd_sc_hs__inv_4_86 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_87/Y sky130_fd_sc_hs__inv_4_87/A
+ sky130_fd_sc_hs__inv_4
Xsky130_fd_sc_hs__inv_4_75 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_75/Y sky130_fd_sc_hs__inv_4_75/A
+ sky130_fd_sc_hs__inv_4
Xsky130_fd_sc_hs__inv_4_64 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_65/Y sky130_fd_sc_hs__inv_4_65/A
+ sky130_fd_sc_hs__inv_4
Xsky130_fd_sc_hs__inv_4_97 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_97/Y sky130_fd_sc_hs__inv_4_97/A
+ sky130_fd_sc_hs__inv_4
Xsky130_fd_sc_hs__o21ai_1_9 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__o21ai_1_9/Y sky130_fd_sc_hs__nand2_2_7/Y
+ sky130_fd_sc_hs__nand2_2_7/B sky130_fd_sc_hs__inv_2_9/A sky130_fd_sc_hs__o21ai_1_9/a_162_368#
+ sky130_fd_sc_hs__o21ai_1_9/a_27_74# sky130_fd_sc_hs__o21ai_1
Xsky130_fd_sc_hs__nor3_1_1 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nor3_1_1/Y sky130_fd_sc_hs__nor3_1_1/C
+ sky130_fd_sc_hs__nor3_1_1/B sky130_fd_sc_hs__nor3_1_1/A sky130_fd_sc_hs__nor3_1_1/a_198_368#
+ sky130_fd_sc_hs__nor3_1_1/a_114_368# sky130_fd_sc_hs__nor3_1
Xsky130_fd_sc_hs__a211oi_1_0 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_27/Y sky130_fd_sc_hs__a211oi_1_1/Y
+ sky130_fd_sc_hs__inv_4_25/Y sky130_fd_sc_hs__nor2b_1_23/Y sky130_fd_sc_hs__o21a_1_15/A1
+ sky130_fd_sc_hs__a211oi_1_1/a_354_368# sky130_fd_sc_hs__a211oi_1_1/a_71_368# sky130_fd_sc_hs__a211oi_1_1/a_159_74#
+ sky130_fd_sc_hs__a211oi_1
Xsky130_fd_sc_hs__a22oi_1_1 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nor2_1_33/Y sky130_fd_sc_hs__a22oi_1_1/Y
+ sky130_fd_sc_hs__inv_4_3/A sky130_fd_sc_hs__and2_2_1/X sky130_fd_sc_hs__inv_4_9/A
+ sky130_fd_sc_hs__a22oi_1_1/a_71_368# sky130_fd_sc_hs__a22oi_1_1/a_159_74# sky130_fd_sc_hs__a22oi_1_1/a_339_74#
+ sky130_fd_sc_hs__a22oi_1
Xsky130_fd_sc_hs__dfrbp_1_20 DVSS DVDD sky130_fd_sc_hs__clkbuf_8_1/X DVDD DVSS sky130_fd_sc_hs__inv_4_85/A
+ sky130_fd_sc_hs__clkbuf_2_1/X sky130_fd_sc_hs__dfrbp_1_21/D sky130_fd_sc_hs__dfrbp_1_21/Q_N
+ sky130_fd_sc_hs__dfrbp_1_21/a_498_360# sky130_fd_sc_hs__dfrbp_1_21/a_1224_74# sky130_fd_sc_hs__dfrbp_1_21/a_2026_424#
+ sky130_fd_sc_hs__dfrbp_1_21/a_1482_48# sky130_fd_sc_hs__dfrbp_1_21/a_125_78# sky130_fd_sc_hs__dfrbp_1_21/a_796_463#
+ sky130_fd_sc_hs__dfrbp_1_21/a_910_118# sky130_fd_sc_hs__dfrbp_1_21/a_1465_471# sky130_fd_sc_hs__dfrbp_1_21/a_832_118#
+ sky130_fd_sc_hs__dfrbp_1_21/a_841_401# sky130_fd_sc_hs__dfrbp_1_21/a_38_78# sky130_fd_sc_hs__dfrbp_1_21/a_1434_74#
+ sky130_fd_sc_hs__dfrbp_1_21/a_706_463# sky130_fd_sc_hs__dfrbp_1_21/a_319_360# sky130_fd_sc_hs__dfrbp_1_21/a_1624_74#
+ sky130_fd_sc_hs__dfrbp_1
Xsky130_fd_sc_hs__dfrbp_1_31 DVSS DVDD sky130_fd_sc_hs__clkbuf_8_1/X DVDD DVSS sky130_fd_sc_hs__nor2_1_95/A
+ ref_clk sky130_fd_sc_hs__dfrbp_1_31/D sky130_fd_sc_hs__dfrbp_1_31/Q_N sky130_fd_sc_hs__dfrbp_1_31/a_498_360#
+ sky130_fd_sc_hs__dfrbp_1_31/a_1224_74# sky130_fd_sc_hs__dfrbp_1_31/a_2026_424# sky130_fd_sc_hs__dfrbp_1_31/a_1482_48#
+ sky130_fd_sc_hs__dfrbp_1_31/a_125_78# sky130_fd_sc_hs__dfrbp_1_31/a_796_463# sky130_fd_sc_hs__dfrbp_1_31/a_910_118#
+ sky130_fd_sc_hs__dfrbp_1_31/a_1465_471# sky130_fd_sc_hs__dfrbp_1_31/a_832_118# sky130_fd_sc_hs__dfrbp_1_31/a_841_401#
+ sky130_fd_sc_hs__dfrbp_1_31/a_38_78# sky130_fd_sc_hs__dfrbp_1_31/a_1434_74# sky130_fd_sc_hs__dfrbp_1_31/a_706_463#
+ sky130_fd_sc_hs__dfrbp_1_31/a_319_360# sky130_fd_sc_hs__dfrbp_1_31/a_1624_74# sky130_fd_sc_hs__dfrbp_1
Xsky130_fd_sc_hs__dfrbp_1_42 DVSS DVDD sky130_fd_sc_hs__clkbuf_8_1/X DVDD DVSS sky130_fd_sc_hs__inv_4_137/A
+ ref_clk sky130_fd_sc_hs__dfrbp_1_43/D sky130_fd_sc_hs__dfrbp_1_43/Q_N sky130_fd_sc_hs__dfrbp_1_43/a_498_360#
+ sky130_fd_sc_hs__dfrbp_1_43/a_1224_74# sky130_fd_sc_hs__dfrbp_1_43/a_2026_424# sky130_fd_sc_hs__dfrbp_1_43/a_1482_48#
+ sky130_fd_sc_hs__dfrbp_1_43/a_125_78# sky130_fd_sc_hs__dfrbp_1_43/a_796_463# sky130_fd_sc_hs__dfrbp_1_43/a_910_118#
+ sky130_fd_sc_hs__dfrbp_1_43/a_1465_471# sky130_fd_sc_hs__dfrbp_1_43/a_832_118# sky130_fd_sc_hs__dfrbp_1_43/a_841_401#
+ sky130_fd_sc_hs__dfrbp_1_43/a_38_78# sky130_fd_sc_hs__dfrbp_1_43/a_1434_74# sky130_fd_sc_hs__dfrbp_1_43/a_706_463#
+ sky130_fd_sc_hs__dfrbp_1_43/a_319_360# sky130_fd_sc_hs__dfrbp_1_43/a_1624_74# sky130_fd_sc_hs__dfrbp_1
Xsky130_fd_sc_hs__nand2_2_10 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_2_11/Y sky130_fd_sc_hs__nand2_2_7/Y
+ sky130_fd_sc_hs__o21ai_1_11/Y sky130_fd_sc_hs__nand2_2_11/a_27_74# sky130_fd_sc_hs__nand2_2
Xsky130_fd_sc_hs__dfxtp_2_9 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_2_5/A sky130_fd_sc_hs__dfxtp_4_9/CLK
+ sky130_fd_sc_hs__nor2_1_77/Y sky130_fd_sc_hs__dfxtp_2_9/a_431_508# sky130_fd_sc_hs__dfxtp_2_9/a_1125_508#
+ sky130_fd_sc_hs__dfxtp_2_9/a_206_368# sky130_fd_sc_hs__dfxtp_2_9/a_27_74# sky130_fd_sc_hs__dfxtp_2_9/a_708_101#
+ sky130_fd_sc_hs__dfxtp_2_9/a_1019_424# sky130_fd_sc_hs__dfxtp_2_9/a_1172_124# sky130_fd_sc_hs__dfxtp_2_9/a_644_504#
+ sky130_fd_sc_hs__dfxtp_2_9/a_1217_314# sky130_fd_sc_hs__dfxtp_2_9/a_538_429# sky130_fd_sc_hs__dfxtp_2_9/a_695_459#
+ sky130_fd_sc_hs__dfxtp_2
Xsky130_fd_sc_hs__o31ai_1_3 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_63/Y sky130_fd_sc_hs__nor2_1_65/Y
+ sky130_fd_sc_hs__o31ai_1_3/B1 sky130_fd_sc_hs__inv_4_67/A sky130_fd_sc_hs__o31ai_1_3/Y
+ sky130_fd_sc_hs__o31ai_1_3/a_114_74# sky130_fd_sc_hs__o31ai_1_3/a_119_368# sky130_fd_sc_hs__o31ai_1_3/a_203_368#
+ sky130_fd_sc_hs__o31ai_1
Xsky130_fd_sc_hs__a21oi_1_0 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nor2_1_1/Y sky130_fd_sc_hs__a21oi_1_1/Y
+ sky130_fd_sc_hs__inv_4_1/Y sky130_fd_sc_hs__inv_4_5/Y sky130_fd_sc_hs__a21oi_1_1/a_117_74#
+ sky130_fd_sc_hs__a21oi_1_1/a_29_368# sky130_fd_sc_hs__a21oi_1
Xsky130_fd_sc_hs__nand4_2_0 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand4_2_1/Y sky130_fd_sc_hs__nand4_2_1/C
+ sky130_fd_sc_hs__nand4_2_1/D sky130_fd_sc_hs__nand4_2_1/B sky130_fd_sc_hs__nor2_2_3/Y
+ sky130_fd_sc_hs__nand4_2_1/a_304_74# sky130_fd_sc_hs__nand4_2_1/a_27_74# sky130_fd_sc_hs__nand4_2_1/a_515_74#
+ sky130_fd_sc_hs__nand4_2
Xsky130_fd_sc_hs__dfrtn_1_10 DVSS DVDD sky130_fd_sc_hs__clkbuf_8_1/X DVDD DVSS sky130_fd_sc_hs__clkbuf_2_1/X
+ sky130_fd_sc_hs__nor2_1_69/B sky130_fd_sc_hs__o21a_1_39/X sky130_fd_sc_hs__dfrtn_1_11/a_1266_119#
+ sky130_fd_sc_hs__dfrtn_1_11/a_1736_119# sky130_fd_sc_hs__dfrtn_1_11/a_817_508# sky130_fd_sc_hs__dfrtn_1_11/a_120_74#
+ sky130_fd_sc_hs__dfrtn_1_11/a_1547_508# sky130_fd_sc_hs__dfrtn_1_11/a_922_127# sky130_fd_sc_hs__dfrtn_1_11/a_33_74#
+ sky130_fd_sc_hs__dfrtn_1_11/a_714_127# sky130_fd_sc_hs__dfrtn_1_11/a_1934_94# sky130_fd_sc_hs__dfrtn_1_11/a_1550_119#
+ sky130_fd_sc_hs__dfrtn_1_11/a_1598_93# sky130_fd_sc_hs__dfrtn_1_11/a_300_74# sky130_fd_sc_hs__dfrtn_1_11/a_507_368#
+ sky130_fd_sc_hs__dfrtn_1_11/a_856_304# sky130_fd_sc_hs__dfrtn_1_11/a_850_127# sky130_fd_sc_hs__dfrtn_1
Xsky130_fd_sc_hs__dfrtn_1_32 DVSS DVDD sky130_fd_sc_hs__clkbuf_8_1/X DVDD DVSS ref_clk
+ sky130_fd_sc_hs__inv_4_105/A sky130_fd_sc_hs__dfrtn_1_33/D sky130_fd_sc_hs__dfrtn_1_33/a_1266_119#
+ sky130_fd_sc_hs__dfrtn_1_33/a_1736_119# sky130_fd_sc_hs__dfrtn_1_33/a_817_508# sky130_fd_sc_hs__dfrtn_1_33/a_120_74#
+ sky130_fd_sc_hs__dfrtn_1_33/a_1547_508# sky130_fd_sc_hs__dfrtn_1_33/a_922_127# sky130_fd_sc_hs__dfrtn_1_33/a_33_74#
+ sky130_fd_sc_hs__dfrtn_1_33/a_714_127# sky130_fd_sc_hs__dfrtn_1_33/a_1934_94# sky130_fd_sc_hs__dfrtn_1_33/a_1550_119#
+ sky130_fd_sc_hs__dfrtn_1_33/a_1598_93# sky130_fd_sc_hs__dfrtn_1_33/a_300_74# sky130_fd_sc_hs__dfrtn_1_33/a_507_368#
+ sky130_fd_sc_hs__dfrtn_1_33/a_856_304# sky130_fd_sc_hs__dfrtn_1_33/a_850_127# sky130_fd_sc_hs__dfrtn_1
Xsky130_fd_sc_hs__nand2_1_105 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_135/Y sky130_fd_sc_hs__maj3_1_3/C
+ sky130_fd_sc_hs__inv_4_125/A sky130_fd_sc_hs__nand2_1_105/a_117_74# sky130_fd_sc_hs__nand2_1
Xsky130_fd_sc_hs__dfrtn_1_43 DVSS DVDD sky130_fd_sc_hs__clkbuf_8_1/X DVDD DVSS ref_clk
+ sky130_fd_sc_hs__inv_4_101/A sky130_fd_sc_hs__o21a_1_65/X sky130_fd_sc_hs__dfrtn_1_43/a_1266_119#
+ sky130_fd_sc_hs__dfrtn_1_43/a_1736_119# sky130_fd_sc_hs__dfrtn_1_43/a_817_508# sky130_fd_sc_hs__dfrtn_1_43/a_120_74#
+ sky130_fd_sc_hs__dfrtn_1_43/a_1547_508# sky130_fd_sc_hs__dfrtn_1_43/a_922_127# sky130_fd_sc_hs__dfrtn_1_43/a_33_74#
+ sky130_fd_sc_hs__dfrtn_1_43/a_714_127# sky130_fd_sc_hs__dfrtn_1_43/a_1934_94# sky130_fd_sc_hs__dfrtn_1_43/a_1550_119#
+ sky130_fd_sc_hs__dfrtn_1_43/a_1598_93# sky130_fd_sc_hs__dfrtn_1_43/a_300_74# sky130_fd_sc_hs__dfrtn_1_43/a_507_368#
+ sky130_fd_sc_hs__dfrtn_1_43/a_856_304# sky130_fd_sc_hs__dfrtn_1_43/a_850_127# sky130_fd_sc_hs__dfrtn_1
Xsky130_fd_sc_hs__nand2_1_116 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_2_7/Y sky130_fd_sc_hs__nand3_1_1/B
+ sky130_fd_sc_hs__inv_2_7/A sky130_fd_sc_hs__nand2_1_117/a_117_74# sky130_fd_sc_hs__nand2_1
Xsky130_fd_sc_hs__dfrtn_1_21 DVSS DVDD sky130_fd_sc_hs__clkbuf_8_1/X DVDD DVSS sky130_fd_sc_hs__clkbuf_2_1/X
+ sky130_fd_sc_hs__inv_4_83/A sky130_fd_sc_hs__o21a_1_49/X sky130_fd_sc_hs__dfrtn_1_21/a_1266_119#
+ sky130_fd_sc_hs__dfrtn_1_21/a_1736_119# sky130_fd_sc_hs__dfrtn_1_21/a_817_508# sky130_fd_sc_hs__dfrtn_1_21/a_120_74#
+ sky130_fd_sc_hs__dfrtn_1_21/a_1547_508# sky130_fd_sc_hs__dfrtn_1_21/a_922_127# sky130_fd_sc_hs__dfrtn_1_21/a_33_74#
+ sky130_fd_sc_hs__dfrtn_1_21/a_714_127# sky130_fd_sc_hs__dfrtn_1_21/a_1934_94# sky130_fd_sc_hs__dfrtn_1_21/a_1550_119#
+ sky130_fd_sc_hs__dfrtn_1_21/a_1598_93# sky130_fd_sc_hs__dfrtn_1_21/a_300_74# sky130_fd_sc_hs__dfrtn_1_21/a_507_368#
+ sky130_fd_sc_hs__dfrtn_1_21/a_856_304# sky130_fd_sc_hs__dfrtn_1_21/a_850_127# sky130_fd_sc_hs__dfrtn_1
Xsky130_fd_sc_hs__nor2_1_19 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nor2_1_19/B sky130_fd_sc_hs__o21a_1_7/A2
+ sky130_fd_sc_hs__inv_4_29/Y sky130_fd_sc_hs__nor2_1_19/a_116_368# sky130_fd_sc_hs__nor2_1
Xsky130_fd_sc_hs__nor2b_1_19 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__fa_2_21/SUM sky130_fd_sc_hs__nor2b_1_19/Y
+ sky130_fd_sc_hs__or2_1_1/A sky130_fd_sc_hs__nor2b_1_19/a_278_368# sky130_fd_sc_hs__nor2b_1_19/a_27_112#
+ sky130_fd_sc_hs__nor2b_1
Xsky130_fd_sc_hs__dfstp_2_3 DVSS DVDD sky130_fd_sc_hs__inv_4_49/Y DVDD DVSS sky130_fd_sc_hs__o21ai_1_1/Y
+ sky130_fd_sc_hs__dfstp_2_5/D sky130_fd_sc_hs__or2_1_1/A sky130_fd_sc_hs__dfstp_2_5/a_1566_92#
+ sky130_fd_sc_hs__dfstp_2_5/a_1521_508# sky130_fd_sc_hs__dfstp_2_5/a_716_456# sky130_fd_sc_hs__dfstp_2_5/a_1266_341#
+ sky130_fd_sc_hs__dfstp_2_5/a_1278_74# sky130_fd_sc_hs__dfstp_2_5/a_398_74# sky130_fd_sc_hs__dfstp_2_5/a_1057_118#
+ sky130_fd_sc_hs__dfstp_2_5/a_1489_118# sky130_fd_sc_hs__dfstp_2_5/a_27_74# sky130_fd_sc_hs__dfstp_2_5/a_1596_118#
+ sky130_fd_sc_hs__dfstp_2_5/a_225_74# sky130_fd_sc_hs__dfstp_2_5/a_1356_74# sky130_fd_sc_hs__dfstp_2_5/a_612_74#
+ sky130_fd_sc_hs__dfstp_2_5/a_781_74# sky130_fd_sc_hs__dfstp_2_5/a_767_384# sky130_fd_sc_hs__dfstp_2_5/a_2022_94#
+ sky130_fd_sc_hs__dfstp_2
Xsky130_fd_sc_hs__dfrtp_4_5 DVSS DVDD sky130_fd_sc_hs__clkbuf_8_1/X DVDD DVSS sky130_fd_sc_hs__dfrtp_4_5/D
+ sky130_fd_sc_hs__nand2_1_47/B sky130_fd_sc_hs__inv_4_7/A sky130_fd_sc_hs__dfrtp_4_5/a_37_78#
+ sky130_fd_sc_hs__dfrtp_4_5/a_494_366# sky130_fd_sc_hs__dfrtp_4_5/a_699_463# sky130_fd_sc_hs__dfrtp_4_5/a_313_74#
+ sky130_fd_sc_hs__dfrtp_4_5/a_1627_493# sky130_fd_sc_hs__dfrtp_4_5/a_1678_395# sky130_fd_sc_hs__dfrtp_4_5/a_1827_81#
+ sky130_fd_sc_hs__dfrtp_4_5/a_789_463# sky130_fd_sc_hs__dfrtp_4_5/a_1350_392# sky130_fd_sc_hs__dfrtp_4_5/a_834_355#
+ sky130_fd_sc_hs__dfrtp_4_5/a_812_138# sky130_fd_sc_hs__dfrtp_4_5/a_124_78# sky130_fd_sc_hs__dfrtp_4_5/a_1647_81#
+ sky130_fd_sc_hs__dfrtp_4_5/a_2010_409# sky130_fd_sc_hs__dfrtp_4_5/a_890_138# sky130_fd_sc_hs__dfrtp_4
Xsky130_fd_sc_hs__inv_4_10 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nor2_1_7/A sky130_fd_sc_hs__inv_4_11/A
+ sky130_fd_sc_hs__inv_4
Xsky130_fd_sc_hs__inv_4_54 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_55/Y sky130_fd_sc_hs__inv_4_55/A
+ sky130_fd_sc_hs__inv_4
Xsky130_fd_sc_hs__inv_4_43 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_43/Y fftl_en
+ sky130_fd_sc_hs__inv_4
Xsky130_fd_sc_hs__inv_4_32 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_33/Y fine_control_avg_window_select[0]
+ sky130_fd_sc_hs__inv_4
Xsky130_fd_sc_hs__inv_4_21 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_21/Y fine_control_avg_window_select[1]
+ sky130_fd_sc_hs__inv_4
Xsky130_fd_sc_hs__inv_4_87 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_87/Y sky130_fd_sc_hs__inv_4_87/A
+ sky130_fd_sc_hs__inv_4
Xsky130_fd_sc_hs__inv_4_76 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_77/Y sky130_fd_sc_hs__nor3_1_1/B
+ sky130_fd_sc_hs__inv_4
Xsky130_fd_sc_hs__inv_4_65 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_65/Y sky130_fd_sc_hs__inv_4_65/A
+ sky130_fd_sc_hs__inv_4
Xsky130_fd_sc_hs__inv_4_98 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_99/Y sky130_fd_sc_hs__inv_4_99/A
+ sky130_fd_sc_hs__inv_4
Xsky130_fd_sc_hs__nor3_1_2 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nor3_1_3/Y sky130_fd_sc_hs__nor3_1_3/C
+ sky130_fd_sc_hs__nor3_1_3/B sky130_fd_sc_hs__nor3_1_3/A sky130_fd_sc_hs__nor3_1_3/a_198_368#
+ sky130_fd_sc_hs__nor3_1_3/a_114_368# sky130_fd_sc_hs__nor3_1
Xsky130_fd_sc_hs__xnor2_1_10 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__o21ai_1_9/Y sky130_fd_sc_hs__xnor2_1_11/Y
+ sky130_fd_sc_hs__nand2_2_5/B sky130_fd_sc_hs__xnor2_1_11/a_376_368# sky130_fd_sc_hs__xnor2_1_11/a_112_119#
+ sky130_fd_sc_hs__xnor2_1_11/a_138_385# sky130_fd_sc_hs__xnor2_1_11/a_293_74# sky130_fd_sc_hs__xnor2_1
Xsky130_fd_sc_hs__a211oi_1_1 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_27/Y sky130_fd_sc_hs__a211oi_1_1/Y
+ sky130_fd_sc_hs__inv_4_25/Y sky130_fd_sc_hs__nor2b_1_23/Y sky130_fd_sc_hs__o21a_1_15/A1
+ sky130_fd_sc_hs__a211oi_1_1/a_354_368# sky130_fd_sc_hs__a211oi_1_1/a_71_368# sky130_fd_sc_hs__a211oi_1_1/a_159_74#
+ sky130_fd_sc_hs__a211oi_1
Xsky130_fd_sc_hs__a22oi_1_2 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nor2b_1_25/Y sky130_fd_sc_hs__nand2_2_1/A
+ sky130_fd_sc_hs__nand2_1_9/A sky130_fd_sc_hs__nor2b_1_23/Y sky130_fd_sc_hs__o21a_1_1/A1
+ sky130_fd_sc_hs__a22oi_1_3/a_71_368# sky130_fd_sc_hs__a22oi_1_3/a_159_74# sky130_fd_sc_hs__a22oi_1_3/a_339_74#
+ sky130_fd_sc_hs__a22oi_1
Xsky130_fd_sc_hs__dfrbp_1_21 DVSS DVDD sky130_fd_sc_hs__clkbuf_8_1/X DVDD DVSS sky130_fd_sc_hs__inv_4_85/A
+ sky130_fd_sc_hs__clkbuf_2_1/X sky130_fd_sc_hs__dfrbp_1_21/D sky130_fd_sc_hs__dfrbp_1_21/Q_N
+ sky130_fd_sc_hs__dfrbp_1_21/a_498_360# sky130_fd_sc_hs__dfrbp_1_21/a_1224_74# sky130_fd_sc_hs__dfrbp_1_21/a_2026_424#
+ sky130_fd_sc_hs__dfrbp_1_21/a_1482_48# sky130_fd_sc_hs__dfrbp_1_21/a_125_78# sky130_fd_sc_hs__dfrbp_1_21/a_796_463#
+ sky130_fd_sc_hs__dfrbp_1_21/a_910_118# sky130_fd_sc_hs__dfrbp_1_21/a_1465_471# sky130_fd_sc_hs__dfrbp_1_21/a_832_118#
+ sky130_fd_sc_hs__dfrbp_1_21/a_841_401# sky130_fd_sc_hs__dfrbp_1_21/a_38_78# sky130_fd_sc_hs__dfrbp_1_21/a_1434_74#
+ sky130_fd_sc_hs__dfrbp_1_21/a_706_463# sky130_fd_sc_hs__dfrbp_1_21/a_319_360# sky130_fd_sc_hs__dfrbp_1_21/a_1624_74#
+ sky130_fd_sc_hs__dfrbp_1
Xsky130_fd_sc_hs__dfrbp_1_10 DVSS DVDD sky130_fd_sc_hs__clkbuf_8_1/X DVDD DVSS sky130_fd_sc_hs__inv_4_79/A
+ sky130_fd_sc_hs__clkbuf_2_1/X sky130_fd_sc_hs__dfrbp_1_11/D sky130_fd_sc_hs__dfrbp_1_11/Q_N
+ sky130_fd_sc_hs__dfrbp_1_11/a_498_360# sky130_fd_sc_hs__dfrbp_1_11/a_1224_74# sky130_fd_sc_hs__dfrbp_1_11/a_2026_424#
+ sky130_fd_sc_hs__dfrbp_1_11/a_1482_48# sky130_fd_sc_hs__dfrbp_1_11/a_125_78# sky130_fd_sc_hs__dfrbp_1_11/a_796_463#
+ sky130_fd_sc_hs__dfrbp_1_11/a_910_118# sky130_fd_sc_hs__dfrbp_1_11/a_1465_471# sky130_fd_sc_hs__dfrbp_1_11/a_832_118#
+ sky130_fd_sc_hs__dfrbp_1_11/a_841_401# sky130_fd_sc_hs__dfrbp_1_11/a_38_78# sky130_fd_sc_hs__dfrbp_1_11/a_1434_74#
+ sky130_fd_sc_hs__dfrbp_1_11/a_706_463# sky130_fd_sc_hs__dfrbp_1_11/a_319_360# sky130_fd_sc_hs__dfrbp_1_11/a_1624_74#
+ sky130_fd_sc_hs__dfrbp_1
Xsky130_fd_sc_hs__dfrbp_1_32 DVSS DVDD sky130_fd_sc_hs__clkbuf_8_1/X DVDD DVSS sky130_fd_sc_hs__maj3_1_3/A
+ ref_clk sky130_fd_sc_hs__o21a_1_61/X sky130_fd_sc_hs__dfrbp_1_33/Q_N sky130_fd_sc_hs__dfrbp_1_33/a_498_360#
+ sky130_fd_sc_hs__dfrbp_1_33/a_1224_74# sky130_fd_sc_hs__dfrbp_1_33/a_2026_424# sky130_fd_sc_hs__dfrbp_1_33/a_1482_48#
+ sky130_fd_sc_hs__dfrbp_1_33/a_125_78# sky130_fd_sc_hs__dfrbp_1_33/a_796_463# sky130_fd_sc_hs__dfrbp_1_33/a_910_118#
+ sky130_fd_sc_hs__dfrbp_1_33/a_1465_471# sky130_fd_sc_hs__dfrbp_1_33/a_832_118# sky130_fd_sc_hs__dfrbp_1_33/a_841_401#
+ sky130_fd_sc_hs__dfrbp_1_33/a_38_78# sky130_fd_sc_hs__dfrbp_1_33/a_1434_74# sky130_fd_sc_hs__dfrbp_1_33/a_706_463#
+ sky130_fd_sc_hs__dfrbp_1_33/a_319_360# sky130_fd_sc_hs__dfrbp_1_33/a_1624_74# sky130_fd_sc_hs__dfrbp_1
Xsky130_fd_sc_hs__dfrbp_1_43 DVSS DVDD sky130_fd_sc_hs__clkbuf_8_1/X DVDD DVSS sky130_fd_sc_hs__inv_4_137/A
+ ref_clk sky130_fd_sc_hs__dfrbp_1_43/D sky130_fd_sc_hs__dfrbp_1_43/Q_N sky130_fd_sc_hs__dfrbp_1_43/a_498_360#
+ sky130_fd_sc_hs__dfrbp_1_43/a_1224_74# sky130_fd_sc_hs__dfrbp_1_43/a_2026_424# sky130_fd_sc_hs__dfrbp_1_43/a_1482_48#
+ sky130_fd_sc_hs__dfrbp_1_43/a_125_78# sky130_fd_sc_hs__dfrbp_1_43/a_796_463# sky130_fd_sc_hs__dfrbp_1_43/a_910_118#
+ sky130_fd_sc_hs__dfrbp_1_43/a_1465_471# sky130_fd_sc_hs__dfrbp_1_43/a_832_118# sky130_fd_sc_hs__dfrbp_1_43/a_841_401#
+ sky130_fd_sc_hs__dfrbp_1_43/a_38_78# sky130_fd_sc_hs__dfrbp_1_43/a_1434_74# sky130_fd_sc_hs__dfrbp_1_43/a_706_463#
+ sky130_fd_sc_hs__dfrbp_1_43/a_319_360# sky130_fd_sc_hs__dfrbp_1_43/a_1624_74# sky130_fd_sc_hs__dfrbp_1
Xsky130_fd_sc_hs__nand2_2_11 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_2_11/Y sky130_fd_sc_hs__nand2_2_7/Y
+ sky130_fd_sc_hs__o21ai_1_11/Y sky130_fd_sc_hs__nand2_2_11/a_27_74# sky130_fd_sc_hs__nand2_2
Xsky130_fd_sc_hs__o31ai_1_4 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_59/Y sky130_fd_sc_hs__nor3_1_1/B
+ sky130_fd_sc_hs__nand4_1_1/D sky130_fd_sc_hs__inv_4_79/A sky130_fd_sc_hs__o31ai_1_5/Y
+ sky130_fd_sc_hs__o31ai_1_5/a_114_74# sky130_fd_sc_hs__o31ai_1_5/a_119_368# sky130_fd_sc_hs__o31ai_1_5/a_203_368#
+ sky130_fd_sc_hs__o31ai_1
Xsky130_fd_sc_hs__a21oi_1_1 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nor2_1_1/Y sky130_fd_sc_hs__a21oi_1_1/Y
+ sky130_fd_sc_hs__inv_4_1/Y sky130_fd_sc_hs__inv_4_5/Y sky130_fd_sc_hs__a21oi_1_1/a_117_74#
+ sky130_fd_sc_hs__a21oi_1_1/a_29_368# sky130_fd_sc_hs__a21oi_1
Xsky130_fd_sc_hs__nand4_2_1 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand4_2_1/Y sky130_fd_sc_hs__nand4_2_1/C
+ sky130_fd_sc_hs__nand4_2_1/D sky130_fd_sc_hs__nand4_2_1/B sky130_fd_sc_hs__nor2_2_3/Y
+ sky130_fd_sc_hs__nand4_2_1/a_304_74# sky130_fd_sc_hs__nand4_2_1/a_27_74# sky130_fd_sc_hs__nand4_2_1/a_515_74#
+ sky130_fd_sc_hs__nand4_2
Xsky130_fd_sc_hs__dfrtn_1_11 DVSS DVDD sky130_fd_sc_hs__clkbuf_8_1/X DVDD DVSS sky130_fd_sc_hs__clkbuf_2_1/X
+ sky130_fd_sc_hs__nor2_1_69/B sky130_fd_sc_hs__o21a_1_39/X sky130_fd_sc_hs__dfrtn_1_11/a_1266_119#
+ sky130_fd_sc_hs__dfrtn_1_11/a_1736_119# sky130_fd_sc_hs__dfrtn_1_11/a_817_508# sky130_fd_sc_hs__dfrtn_1_11/a_120_74#
+ sky130_fd_sc_hs__dfrtn_1_11/a_1547_508# sky130_fd_sc_hs__dfrtn_1_11/a_922_127# sky130_fd_sc_hs__dfrtn_1_11/a_33_74#
+ sky130_fd_sc_hs__dfrtn_1_11/a_714_127# sky130_fd_sc_hs__dfrtn_1_11/a_1934_94# sky130_fd_sc_hs__dfrtn_1_11/a_1550_119#
+ sky130_fd_sc_hs__dfrtn_1_11/a_1598_93# sky130_fd_sc_hs__dfrtn_1_11/a_300_74# sky130_fd_sc_hs__dfrtn_1_11/a_507_368#
+ sky130_fd_sc_hs__dfrtn_1_11/a_856_304# sky130_fd_sc_hs__dfrtn_1_11/a_850_127# sky130_fd_sc_hs__dfrtn_1
Xsky130_fd_sc_hs__dfrtn_1_33 DVSS DVDD sky130_fd_sc_hs__clkbuf_8_1/X DVDD DVSS ref_clk
+ sky130_fd_sc_hs__inv_4_105/A sky130_fd_sc_hs__dfrtn_1_33/D sky130_fd_sc_hs__dfrtn_1_33/a_1266_119#
+ sky130_fd_sc_hs__dfrtn_1_33/a_1736_119# sky130_fd_sc_hs__dfrtn_1_33/a_817_508# sky130_fd_sc_hs__dfrtn_1_33/a_120_74#
+ sky130_fd_sc_hs__dfrtn_1_33/a_1547_508# sky130_fd_sc_hs__dfrtn_1_33/a_922_127# sky130_fd_sc_hs__dfrtn_1_33/a_33_74#
+ sky130_fd_sc_hs__dfrtn_1_33/a_714_127# sky130_fd_sc_hs__dfrtn_1_33/a_1934_94# sky130_fd_sc_hs__dfrtn_1_33/a_1550_119#
+ sky130_fd_sc_hs__dfrtn_1_33/a_1598_93# sky130_fd_sc_hs__dfrtn_1_33/a_300_74# sky130_fd_sc_hs__dfrtn_1_33/a_507_368#
+ sky130_fd_sc_hs__dfrtn_1_33/a_856_304# sky130_fd_sc_hs__dfrtn_1_33/a_850_127# sky130_fd_sc_hs__dfrtn_1
Xsky130_fd_sc_hs__nand2_1_106 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__o21a_1_69/A2 sky130_fd_sc_hs__xnor2_1_9/B
+ sky130_fd_sc_hs__inv_4_127/A sky130_fd_sc_hs__nand2_1_107/a_117_74# sky130_fd_sc_hs__nand2_1
Xsky130_fd_sc_hs__dfrtn_1_44 DVSS DVDD sky130_fd_sc_hs__clkbuf_8_1/X DVDD DVSS ref_clk
+ sky130_fd_sc_hs__inv_4_133/A sky130_fd_sc_hs__o21a_1_67/X sky130_fd_sc_hs__dfrtn_1_45/a_1266_119#
+ sky130_fd_sc_hs__dfrtn_1_45/a_1736_119# sky130_fd_sc_hs__dfrtn_1_45/a_817_508# sky130_fd_sc_hs__dfrtn_1_45/a_120_74#
+ sky130_fd_sc_hs__dfrtn_1_45/a_1547_508# sky130_fd_sc_hs__dfrtn_1_45/a_922_127# sky130_fd_sc_hs__dfrtn_1_45/a_33_74#
+ sky130_fd_sc_hs__dfrtn_1_45/a_714_127# sky130_fd_sc_hs__dfrtn_1_45/a_1934_94# sky130_fd_sc_hs__dfrtn_1_45/a_1550_119#
+ sky130_fd_sc_hs__dfrtn_1_45/a_1598_93# sky130_fd_sc_hs__dfrtn_1_45/a_300_74# sky130_fd_sc_hs__dfrtn_1_45/a_507_368#
+ sky130_fd_sc_hs__dfrtn_1_45/a_856_304# sky130_fd_sc_hs__dfrtn_1_45/a_850_127# sky130_fd_sc_hs__dfrtn_1
Xsky130_fd_sc_hs__nand2_1_117 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_2_7/Y sky130_fd_sc_hs__nand3_1_1/B
+ sky130_fd_sc_hs__inv_2_7/A sky130_fd_sc_hs__nand2_1_117/a_117_74# sky130_fd_sc_hs__nand2_1
Xsky130_fd_sc_hs__dfrtn_1_22 DVSS DVDD sky130_fd_sc_hs__clkbuf_8_1/X DVDD DVSS sky130_fd_sc_hs__clkbuf_2_1/X
+ sky130_fd_sc_hs__inv_4_81/A sky130_fd_sc_hs__dfrtn_1_23/D sky130_fd_sc_hs__dfrtn_1_23/a_1266_119#
+ sky130_fd_sc_hs__dfrtn_1_23/a_1736_119# sky130_fd_sc_hs__dfrtn_1_23/a_817_508# sky130_fd_sc_hs__dfrtn_1_23/a_120_74#
+ sky130_fd_sc_hs__dfrtn_1_23/a_1547_508# sky130_fd_sc_hs__dfrtn_1_23/a_922_127# sky130_fd_sc_hs__dfrtn_1_23/a_33_74#
+ sky130_fd_sc_hs__dfrtn_1_23/a_714_127# sky130_fd_sc_hs__dfrtn_1_23/a_1934_94# sky130_fd_sc_hs__dfrtn_1_23/a_1550_119#
+ sky130_fd_sc_hs__dfrtn_1_23/a_1598_93# sky130_fd_sc_hs__dfrtn_1_23/a_300_74# sky130_fd_sc_hs__dfrtn_1_23/a_507_368#
+ sky130_fd_sc_hs__dfrtn_1_23/a_856_304# sky130_fd_sc_hs__dfrtn_1_23/a_850_127# sky130_fd_sc_hs__dfrtn_1
Xsky130_fd_sc_hs__dfstp_2_4 DVSS DVDD sky130_fd_sc_hs__inv_4_49/Y DVDD DVSS sky130_fd_sc_hs__o21ai_1_1/Y
+ sky130_fd_sc_hs__nor3_1_3/Y sky130_fd_sc_hs__dfstp_2_5/D sky130_fd_sc_hs__dfstp_2_4/a_1566_92#
+ sky130_fd_sc_hs__dfstp_2_4/a_1521_508# sky130_fd_sc_hs__dfstp_2_4/a_716_456# sky130_fd_sc_hs__dfstp_2_4/a_1266_341#
+ sky130_fd_sc_hs__dfstp_2_4/a_1278_74# sky130_fd_sc_hs__dfstp_2_4/a_398_74# sky130_fd_sc_hs__dfstp_2_4/a_1057_118#
+ sky130_fd_sc_hs__dfstp_2_4/a_1489_118# sky130_fd_sc_hs__dfstp_2_4/a_27_74# sky130_fd_sc_hs__dfstp_2_4/a_1596_118#
+ sky130_fd_sc_hs__dfstp_2_4/a_225_74# sky130_fd_sc_hs__dfstp_2_4/a_1356_74# sky130_fd_sc_hs__dfstp_2_4/a_612_74#
+ sky130_fd_sc_hs__dfstp_2_4/a_781_74# sky130_fd_sc_hs__dfstp_2_4/a_767_384# sky130_fd_sc_hs__dfstp_2_4/a_2022_94#
+ sky130_fd_sc_hs__dfstp_2
Xsky130_fd_sc_hs__dfrtp_4_6 DVSS DVDD sky130_fd_sc_hs__clkbuf_8_1/A DVDD DVSS sky130_fd_sc_hs__dfrtp_4_7/D
+ sky130_fd_sc_hs__nand2_1_47/B sky130_fd_sc_hs__inv_4_9/A sky130_fd_sc_hs__dfrtp_4_7/a_37_78#
+ sky130_fd_sc_hs__dfrtp_4_7/a_494_366# sky130_fd_sc_hs__dfrtp_4_7/a_699_463# sky130_fd_sc_hs__dfrtp_4_7/a_313_74#
+ sky130_fd_sc_hs__dfrtp_4_7/a_1627_493# sky130_fd_sc_hs__dfrtp_4_7/a_1678_395# sky130_fd_sc_hs__dfrtp_4_7/a_1827_81#
+ sky130_fd_sc_hs__dfrtp_4_7/a_789_463# sky130_fd_sc_hs__dfrtp_4_7/a_1350_392# sky130_fd_sc_hs__dfrtp_4_7/a_834_355#
+ sky130_fd_sc_hs__dfrtp_4_7/a_812_138# sky130_fd_sc_hs__dfrtp_4_7/a_124_78# sky130_fd_sc_hs__dfrtp_4_7/a_1647_81#
+ sky130_fd_sc_hs__dfrtp_4_7/a_2010_409# sky130_fd_sc_hs__dfrtp_4_7/a_890_138# sky130_fd_sc_hs__dfrtp_4
Xsky130_fd_sc_hs__inv_4_11 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nor2_1_7/A sky130_fd_sc_hs__inv_4_11/A
+ sky130_fd_sc_hs__inv_4
Xsky130_fd_sc_hs__inv_4_44 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_45/Y sky130_fd_sc_hs__inv_4_45/A
+ sky130_fd_sc_hs__inv_4
Xsky130_fd_sc_hs__inv_4_33 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_33/Y fine_control_avg_window_select[0]
+ sky130_fd_sc_hs__inv_4
Xsky130_fd_sc_hs__inv_4_22 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nor2_4_1/B sky130_fd_sc_hs__inv_4_23/A
+ sky130_fd_sc_hs__inv_4
Xsky130_fd_sc_hs__inv_4_77 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_77/Y sky130_fd_sc_hs__nor3_1_1/B
+ sky130_fd_sc_hs__inv_4
Xsky130_fd_sc_hs__inv_4_66 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_67/Y sky130_fd_sc_hs__inv_4_67/A
+ sky130_fd_sc_hs__inv_4
Xsky130_fd_sc_hs__inv_4_55 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_55/Y sky130_fd_sc_hs__inv_4_55/A
+ sky130_fd_sc_hs__inv_4
Xsky130_fd_sc_hs__inv_4_99 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_99/Y sky130_fd_sc_hs__inv_4_99/A
+ sky130_fd_sc_hs__inv_4
Xsky130_fd_sc_hs__inv_4_88 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_89/Y sky130_fd_sc_hs__inv_4_89/A
+ sky130_fd_sc_hs__inv_4
Xsky130_fd_sc_hs__nor3_1_3 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nor3_1_3/Y sky130_fd_sc_hs__nor3_1_3/C
+ sky130_fd_sc_hs__nor3_1_3/B sky130_fd_sc_hs__nor3_1_3/A sky130_fd_sc_hs__nor3_1_3/a_198_368#
+ sky130_fd_sc_hs__nor3_1_3/a_114_368# sky130_fd_sc_hs__nor3_1
Xsky130_fd_sc_hs__xnor2_1_11 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__o21ai_1_9/Y sky130_fd_sc_hs__xnor2_1_11/Y
+ sky130_fd_sc_hs__nand2_2_5/B sky130_fd_sc_hs__xnor2_1_11/a_376_368# sky130_fd_sc_hs__xnor2_1_11/a_112_119#
+ sky130_fd_sc_hs__xnor2_1_11/a_138_385# sky130_fd_sc_hs__xnor2_1_11/a_293_74# sky130_fd_sc_hs__xnor2_1
Xsky130_fd_sc_hs__a211oi_1_2 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand4_1_1/Y sky130_fd_sc_hs__nand4_1_5/C
+ sky130_fd_sc_hs__o211ai_1_5/Y sky130_fd_sc_hs__inv_4_75/Y sky130_fd_sc_hs__inv_4_85/A
+ sky130_fd_sc_hs__a211oi_1_3/a_354_368# sky130_fd_sc_hs__a211oi_1_3/a_71_368# sky130_fd_sc_hs__a211oi_1_3/a_159_74#
+ sky130_fd_sc_hs__a211oi_1
Xsky130_fd_sc_hs__a22oi_1_3 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nor2b_1_25/Y sky130_fd_sc_hs__nand2_2_1/A
+ sky130_fd_sc_hs__nand2_1_9/A sky130_fd_sc_hs__nor2b_1_23/Y sky130_fd_sc_hs__o21a_1_1/A1
+ sky130_fd_sc_hs__a22oi_1_3/a_71_368# sky130_fd_sc_hs__a22oi_1_3/a_159_74# sky130_fd_sc_hs__a22oi_1_3/a_339_74#
+ sky130_fd_sc_hs__a22oi_1
Xsky130_fd_sc_hs__sdlclkp_4_0 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__conb_1_1/LO sky130_fd_sc_hs__nand2_1_23/Y
+ sky130_fd_sc_hs__o21ai_1_1/Y sky130_fd_sc_hs__dfstp_2_1/CLK sky130_fd_sc_hs__sdlclkp_4_1/a_1289_368#
+ sky130_fd_sc_hs__sdlclkp_4_1/a_744_74# sky130_fd_sc_hs__sdlclkp_4_1/a_785_455# sky130_fd_sc_hs__sdlclkp_4_1/a_634_74#
+ sky130_fd_sc_hs__sdlclkp_4_1/a_1292_74# sky130_fd_sc_hs__sdlclkp_4_1/a_792_48# sky130_fd_sc_hs__sdlclkp_4_1/a_324_79#
+ sky130_fd_sc_hs__sdlclkp_4_1/a_116_395# sky130_fd_sc_hs__sdlclkp_4_1/a_354_105#
+ sky130_fd_sc_hs__sdlclkp_4_1/a_119_143# sky130_fd_sc_hs__sdlclkp_4
Xsky130_fd_sc_hs__dfrbp_1_11 DVSS DVDD sky130_fd_sc_hs__clkbuf_8_1/X DVDD DVSS sky130_fd_sc_hs__inv_4_79/A
+ sky130_fd_sc_hs__clkbuf_2_1/X sky130_fd_sc_hs__dfrbp_1_11/D sky130_fd_sc_hs__dfrbp_1_11/Q_N
+ sky130_fd_sc_hs__dfrbp_1_11/a_498_360# sky130_fd_sc_hs__dfrbp_1_11/a_1224_74# sky130_fd_sc_hs__dfrbp_1_11/a_2026_424#
+ sky130_fd_sc_hs__dfrbp_1_11/a_1482_48# sky130_fd_sc_hs__dfrbp_1_11/a_125_78# sky130_fd_sc_hs__dfrbp_1_11/a_796_463#
+ sky130_fd_sc_hs__dfrbp_1_11/a_910_118# sky130_fd_sc_hs__dfrbp_1_11/a_1465_471# sky130_fd_sc_hs__dfrbp_1_11/a_832_118#
+ sky130_fd_sc_hs__dfrbp_1_11/a_841_401# sky130_fd_sc_hs__dfrbp_1_11/a_38_78# sky130_fd_sc_hs__dfrbp_1_11/a_1434_74#
+ sky130_fd_sc_hs__dfrbp_1_11/a_706_463# sky130_fd_sc_hs__dfrbp_1_11/a_319_360# sky130_fd_sc_hs__dfrbp_1_11/a_1624_74#
+ sky130_fd_sc_hs__dfrbp_1
Xsky130_fd_sc_hs__dfrbp_1_33 DVSS DVDD sky130_fd_sc_hs__clkbuf_8_1/X DVDD DVSS sky130_fd_sc_hs__maj3_1_3/A
+ ref_clk sky130_fd_sc_hs__o21a_1_61/X sky130_fd_sc_hs__dfrbp_1_33/Q_N sky130_fd_sc_hs__dfrbp_1_33/a_498_360#
+ sky130_fd_sc_hs__dfrbp_1_33/a_1224_74# sky130_fd_sc_hs__dfrbp_1_33/a_2026_424# sky130_fd_sc_hs__dfrbp_1_33/a_1482_48#
+ sky130_fd_sc_hs__dfrbp_1_33/a_125_78# sky130_fd_sc_hs__dfrbp_1_33/a_796_463# sky130_fd_sc_hs__dfrbp_1_33/a_910_118#
+ sky130_fd_sc_hs__dfrbp_1_33/a_1465_471# sky130_fd_sc_hs__dfrbp_1_33/a_832_118# sky130_fd_sc_hs__dfrbp_1_33/a_841_401#
+ sky130_fd_sc_hs__dfrbp_1_33/a_38_78# sky130_fd_sc_hs__dfrbp_1_33/a_1434_74# sky130_fd_sc_hs__dfrbp_1_33/a_706_463#
+ sky130_fd_sc_hs__dfrbp_1_33/a_319_360# sky130_fd_sc_hs__dfrbp_1_33/a_1624_74# sky130_fd_sc_hs__dfrbp_1
Xsky130_fd_sc_hs__dfrbp_1_44 DVSS DVDD sky130_fd_sc_hs__clkbuf_8_1/X DVDD DVSS sky130_fd_sc_hs__inv_4_113/A
+ ref_clk sky130_fd_sc_hs__o21a_1_77/X sky130_fd_sc_hs__dfrbp_1_45/Q_N sky130_fd_sc_hs__dfrbp_1_45/a_498_360#
+ sky130_fd_sc_hs__dfrbp_1_45/a_1224_74# sky130_fd_sc_hs__dfrbp_1_45/a_2026_424# sky130_fd_sc_hs__dfrbp_1_45/a_1482_48#
+ sky130_fd_sc_hs__dfrbp_1_45/a_125_78# sky130_fd_sc_hs__dfrbp_1_45/a_796_463# sky130_fd_sc_hs__dfrbp_1_45/a_910_118#
+ sky130_fd_sc_hs__dfrbp_1_45/a_1465_471# sky130_fd_sc_hs__dfrbp_1_45/a_832_118# sky130_fd_sc_hs__dfrbp_1_45/a_841_401#
+ sky130_fd_sc_hs__dfrbp_1_45/a_38_78# sky130_fd_sc_hs__dfrbp_1_45/a_1434_74# sky130_fd_sc_hs__dfrbp_1_45/a_706_463#
+ sky130_fd_sc_hs__dfrbp_1_45/a_319_360# sky130_fd_sc_hs__dfrbp_1_45/a_1624_74# sky130_fd_sc_hs__dfrbp_1
Xsky130_fd_sc_hs__dfrbp_1_22 DVSS DVDD sky130_fd_sc_hs__clkbuf_8_1/X DVDD DVSS sky130_fd_sc_hs__maj3_1_1/A
+ sky130_fd_sc_hs__clkbuf_2_1/X sky130_fd_sc_hs__o21a_1_51/X sky130_fd_sc_hs__dfrbp_1_23/Q_N
+ sky130_fd_sc_hs__dfrbp_1_23/a_498_360# sky130_fd_sc_hs__dfrbp_1_23/a_1224_74# sky130_fd_sc_hs__dfrbp_1_23/a_2026_424#
+ sky130_fd_sc_hs__dfrbp_1_23/a_1482_48# sky130_fd_sc_hs__dfrbp_1_23/a_125_78# sky130_fd_sc_hs__dfrbp_1_23/a_796_463#
+ sky130_fd_sc_hs__dfrbp_1_23/a_910_118# sky130_fd_sc_hs__dfrbp_1_23/a_1465_471# sky130_fd_sc_hs__dfrbp_1_23/a_832_118#
+ sky130_fd_sc_hs__dfrbp_1_23/a_841_401# sky130_fd_sc_hs__dfrbp_1_23/a_38_78# sky130_fd_sc_hs__dfrbp_1_23/a_1434_74#
+ sky130_fd_sc_hs__dfrbp_1_23/a_706_463# sky130_fd_sc_hs__dfrbp_1_23/a_319_360# sky130_fd_sc_hs__dfrbp_1_23/a_1624_74#
+ sky130_fd_sc_hs__dfrbp_1
Xsky130_fd_sc_hs__nand2_2_12 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_2_13/Y div_ratio_half[3]
+ sky130_fd_sc_hs__xnor2_1_3/A sky130_fd_sc_hs__nand2_2_13/a_27_74# sky130_fd_sc_hs__nand2_2
Xsky130_fd_sc_hs__xor2_1_0 DVSS DVDD DVDD DVSS fine_con_step_size[0] sky130_fd_sc_hs__fa_2_9/B
+ sky130_fd_sc_hs__xor2_1_1/X sky130_fd_sc_hs__xor2_1_1/a_194_125# sky130_fd_sc_hs__xor2_1_1/a_355_368#
+ sky130_fd_sc_hs__xor2_1_1/a_455_87# sky130_fd_sc_hs__xor2_1_1/a_158_392# sky130_fd_sc_hs__xor2_1
Xsky130_fd_sc_hs__o31ai_1_5 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_59/Y sky130_fd_sc_hs__nor3_1_1/B
+ sky130_fd_sc_hs__nand4_1_1/D sky130_fd_sc_hs__inv_4_79/A sky130_fd_sc_hs__o31ai_1_5/Y
+ sky130_fd_sc_hs__o31ai_1_5/a_114_74# sky130_fd_sc_hs__o31ai_1_5/a_119_368# sky130_fd_sc_hs__o31ai_1_5/a_203_368#
+ sky130_fd_sc_hs__o31ai_1
Xsky130_fd_sc_hs__a21oi_1_2 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nor2_1_3/Y sky130_fd_sc_hs__dfrtp_4_3/D
+ sky130_fd_sc_hs__nor2_1_3/B sky130_fd_sc_hs__inv_4_3/Y sky130_fd_sc_hs__a21oi_1_3/a_117_74#
+ sky130_fd_sc_hs__a21oi_1_3/a_29_368# sky130_fd_sc_hs__a21oi_1
Xsky130_fd_sc_hs__dfrtn_1_34 DVSS DVDD sky130_fd_sc_hs__clkbuf_8_1/X DVDD DVSS ref_clk
+ sky130_fd_sc_hs__xnor2_1_9/A sky130_fd_sc_hs__xnor2_1_9/Y sky130_fd_sc_hs__dfrtn_1_35/a_1266_119#
+ sky130_fd_sc_hs__dfrtn_1_35/a_1736_119# sky130_fd_sc_hs__dfrtn_1_35/a_817_508# sky130_fd_sc_hs__dfrtn_1_35/a_120_74#
+ sky130_fd_sc_hs__dfrtn_1_35/a_1547_508# sky130_fd_sc_hs__dfrtn_1_35/a_922_127# sky130_fd_sc_hs__dfrtn_1_35/a_33_74#
+ sky130_fd_sc_hs__dfrtn_1_35/a_714_127# sky130_fd_sc_hs__dfrtn_1_35/a_1934_94# sky130_fd_sc_hs__dfrtn_1_35/a_1550_119#
+ sky130_fd_sc_hs__dfrtn_1_35/a_1598_93# sky130_fd_sc_hs__dfrtn_1_35/a_300_74# sky130_fd_sc_hs__dfrtn_1_35/a_507_368#
+ sky130_fd_sc_hs__dfrtn_1_35/a_856_304# sky130_fd_sc_hs__dfrtn_1_35/a_850_127# sky130_fd_sc_hs__dfrtn_1
Xsky130_fd_sc_hs__nand2_1_107 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__o21a_1_69/A2 sky130_fd_sc_hs__xnor2_1_9/B
+ sky130_fd_sc_hs__inv_4_127/A sky130_fd_sc_hs__nand2_1_107/a_117_74# sky130_fd_sc_hs__nand2_1
Xsky130_fd_sc_hs__dfrtn_1_45 DVSS DVDD sky130_fd_sc_hs__clkbuf_8_1/X DVDD DVSS ref_clk
+ sky130_fd_sc_hs__inv_4_133/A sky130_fd_sc_hs__o21a_1_67/X sky130_fd_sc_hs__dfrtn_1_45/a_1266_119#
+ sky130_fd_sc_hs__dfrtn_1_45/a_1736_119# sky130_fd_sc_hs__dfrtn_1_45/a_817_508# sky130_fd_sc_hs__dfrtn_1_45/a_120_74#
+ sky130_fd_sc_hs__dfrtn_1_45/a_1547_508# sky130_fd_sc_hs__dfrtn_1_45/a_922_127# sky130_fd_sc_hs__dfrtn_1_45/a_33_74#
+ sky130_fd_sc_hs__dfrtn_1_45/a_714_127# sky130_fd_sc_hs__dfrtn_1_45/a_1934_94# sky130_fd_sc_hs__dfrtn_1_45/a_1550_119#
+ sky130_fd_sc_hs__dfrtn_1_45/a_1598_93# sky130_fd_sc_hs__dfrtn_1_45/a_300_74# sky130_fd_sc_hs__dfrtn_1_45/a_507_368#
+ sky130_fd_sc_hs__dfrtn_1_45/a_856_304# sky130_fd_sc_hs__dfrtn_1_45/a_850_127# sky130_fd_sc_hs__dfrtn_1
Xsky130_fd_sc_hs__dfrtn_1_23 DVSS DVDD sky130_fd_sc_hs__clkbuf_8_1/X DVDD DVSS sky130_fd_sc_hs__clkbuf_2_1/X
+ sky130_fd_sc_hs__inv_4_81/A sky130_fd_sc_hs__dfrtn_1_23/D sky130_fd_sc_hs__dfrtn_1_23/a_1266_119#
+ sky130_fd_sc_hs__dfrtn_1_23/a_1736_119# sky130_fd_sc_hs__dfrtn_1_23/a_817_508# sky130_fd_sc_hs__dfrtn_1_23/a_120_74#
+ sky130_fd_sc_hs__dfrtn_1_23/a_1547_508# sky130_fd_sc_hs__dfrtn_1_23/a_922_127# sky130_fd_sc_hs__dfrtn_1_23/a_33_74#
+ sky130_fd_sc_hs__dfrtn_1_23/a_714_127# sky130_fd_sc_hs__dfrtn_1_23/a_1934_94# sky130_fd_sc_hs__dfrtn_1_23/a_1550_119#
+ sky130_fd_sc_hs__dfrtn_1_23/a_1598_93# sky130_fd_sc_hs__dfrtn_1_23/a_300_74# sky130_fd_sc_hs__dfrtn_1_23/a_507_368#
+ sky130_fd_sc_hs__dfrtn_1_23/a_856_304# sky130_fd_sc_hs__dfrtn_1_23/a_850_127# sky130_fd_sc_hs__dfrtn_1
Xsky130_fd_sc_hs__dfrtn_1_12 DVSS DVDD sky130_fd_sc_hs__clkbuf_8_1/X DVDD DVSS sky130_fd_sc_hs__clkbuf_2_1/X
+ sky130_fd_sc_hs__inv_4_59/A sky130_fd_sc_hs__dfrtn_1_13/D sky130_fd_sc_hs__dfrtn_1_13/a_1266_119#
+ sky130_fd_sc_hs__dfrtn_1_13/a_1736_119# sky130_fd_sc_hs__dfrtn_1_13/a_817_508# sky130_fd_sc_hs__dfrtn_1_13/a_120_74#
+ sky130_fd_sc_hs__dfrtn_1_13/a_1547_508# sky130_fd_sc_hs__dfrtn_1_13/a_922_127# sky130_fd_sc_hs__dfrtn_1_13/a_33_74#
+ sky130_fd_sc_hs__dfrtn_1_13/a_714_127# sky130_fd_sc_hs__dfrtn_1_13/a_1934_94# sky130_fd_sc_hs__dfrtn_1_13/a_1550_119#
+ sky130_fd_sc_hs__dfrtn_1_13/a_1598_93# sky130_fd_sc_hs__dfrtn_1_13/a_300_74# sky130_fd_sc_hs__dfrtn_1_13/a_507_368#
+ sky130_fd_sc_hs__dfrtn_1_13/a_856_304# sky130_fd_sc_hs__dfrtn_1_13/a_850_127# sky130_fd_sc_hs__dfrtn_1
Xsky130_fd_sc_hs__nand2_1_118 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__o21a_1_75/A2 sky130_fd_sc_hs__o21a_1_75/B1
+ sky130_fd_sc_hs__o21a_1_75/A1 sky130_fd_sc_hs__nand2_1_119/a_117_74# sky130_fd_sc_hs__nand2_1
Xsky130_fd_sc_hs__dfrbp_1_0 DVSS DVDD sky130_fd_sc_hs__clkbuf_8_1/X DVDD DVSS sky130_fd_sc_hs__dfrbp_1_1/Q
+ sky130_fd_sc_hs__clkbuf_2_1/X sky130_fd_sc_hs__o21a_1_35/X sky130_fd_sc_hs__dfrbp_1_1/Q_N
+ sky130_fd_sc_hs__dfrbp_1_1/a_498_360# sky130_fd_sc_hs__dfrbp_1_1/a_1224_74# sky130_fd_sc_hs__dfrbp_1_1/a_2026_424#
+ sky130_fd_sc_hs__dfrbp_1_1/a_1482_48# sky130_fd_sc_hs__dfrbp_1_1/a_125_78# sky130_fd_sc_hs__dfrbp_1_1/a_796_463#
+ sky130_fd_sc_hs__dfrbp_1_1/a_910_118# sky130_fd_sc_hs__dfrbp_1_1/a_1465_471# sky130_fd_sc_hs__dfrbp_1_1/a_832_118#
+ sky130_fd_sc_hs__dfrbp_1_1/a_841_401# sky130_fd_sc_hs__dfrbp_1_1/a_38_78# sky130_fd_sc_hs__dfrbp_1_1/a_1434_74#
+ sky130_fd_sc_hs__dfrbp_1_1/a_706_463# sky130_fd_sc_hs__dfrbp_1_1/a_319_360# sky130_fd_sc_hs__dfrbp_1_1/a_1624_74#
+ sky130_fd_sc_hs__dfrbp_1
Xsky130_fd_sc_hs__dfstp_2_5 DVSS DVDD sky130_fd_sc_hs__inv_4_49/Y DVDD DVSS sky130_fd_sc_hs__o21ai_1_1/Y
+ sky130_fd_sc_hs__dfstp_2_5/D sky130_fd_sc_hs__or2_1_1/A sky130_fd_sc_hs__dfstp_2_5/a_1566_92#
+ sky130_fd_sc_hs__dfstp_2_5/a_1521_508# sky130_fd_sc_hs__dfstp_2_5/a_716_456# sky130_fd_sc_hs__dfstp_2_5/a_1266_341#
+ sky130_fd_sc_hs__dfstp_2_5/a_1278_74# sky130_fd_sc_hs__dfstp_2_5/a_398_74# sky130_fd_sc_hs__dfstp_2_5/a_1057_118#
+ sky130_fd_sc_hs__dfstp_2_5/a_1489_118# sky130_fd_sc_hs__dfstp_2_5/a_27_74# sky130_fd_sc_hs__dfstp_2_5/a_1596_118#
+ sky130_fd_sc_hs__dfstp_2_5/a_225_74# sky130_fd_sc_hs__dfstp_2_5/a_1356_74# sky130_fd_sc_hs__dfstp_2_5/a_612_74#
+ sky130_fd_sc_hs__dfstp_2_5/a_781_74# sky130_fd_sc_hs__dfstp_2_5/a_767_384# sky130_fd_sc_hs__dfstp_2_5/a_2022_94#
+ sky130_fd_sc_hs__dfstp_2
Xsky130_fd_sc_hs__dfrtp_4_7 DVSS DVDD sky130_fd_sc_hs__clkbuf_8_1/A DVDD DVSS sky130_fd_sc_hs__dfrtp_4_7/D
+ sky130_fd_sc_hs__nand2_1_47/B sky130_fd_sc_hs__inv_4_9/A sky130_fd_sc_hs__dfrtp_4_7/a_37_78#
+ sky130_fd_sc_hs__dfrtp_4_7/a_494_366# sky130_fd_sc_hs__dfrtp_4_7/a_699_463# sky130_fd_sc_hs__dfrtp_4_7/a_313_74#
+ sky130_fd_sc_hs__dfrtp_4_7/a_1627_493# sky130_fd_sc_hs__dfrtp_4_7/a_1678_395# sky130_fd_sc_hs__dfrtp_4_7/a_1827_81#
+ sky130_fd_sc_hs__dfrtp_4_7/a_789_463# sky130_fd_sc_hs__dfrtp_4_7/a_1350_392# sky130_fd_sc_hs__dfrtp_4_7/a_834_355#
+ sky130_fd_sc_hs__dfrtp_4_7/a_812_138# sky130_fd_sc_hs__dfrtp_4_7/a_124_78# sky130_fd_sc_hs__dfrtp_4_7/a_1647_81#
+ sky130_fd_sc_hs__dfrtp_4_7/a_2010_409# sky130_fd_sc_hs__dfrtp_4_7/a_890_138# sky130_fd_sc_hs__dfrtp_4
Xsky130_fd_sc_hs__inv_4_45 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_45/Y sky130_fd_sc_hs__inv_4_45/A
+ sky130_fd_sc_hs__inv_4
Xsky130_fd_sc_hs__inv_4_34 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_35/Y sky130_fd_sc_hs__inv_4_35/A
+ sky130_fd_sc_hs__inv_4
Xsky130_fd_sc_hs__inv_4_23 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nor2_4_1/B sky130_fd_sc_hs__inv_4_23/A
+ sky130_fd_sc_hs__inv_4
Xsky130_fd_sc_hs__inv_4_12 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_13/Y sky130_fd_sc_hs__inv_4_13/A
+ sky130_fd_sc_hs__inv_4
Xsky130_fd_sc_hs__inv_4_78 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_79/Y sky130_fd_sc_hs__inv_4_79/A
+ sky130_fd_sc_hs__inv_4
Xsky130_fd_sc_hs__inv_4_67 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_67/Y sky130_fd_sc_hs__inv_4_67/A
+ sky130_fd_sc_hs__inv_4
Xsky130_fd_sc_hs__inv_4_56 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_57/Y out_star
+ sky130_fd_sc_hs__inv_4
Xsky130_fd_sc_hs__inv_4_89 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_89/Y sky130_fd_sc_hs__inv_4_89/A
+ sky130_fd_sc_hs__inv_4
Xsky130_fd_sc_hs__fa_2_0 DVSS DVDD sky130_fd_sc_hs__fa_2_1/A DVDD DVSS sky130_fd_sc_hs__fa_2_1/CIN
+ sky130_fd_sc_hs__fa_2_1/B sky130_fd_sc_hs__fa_2_7/CIN sky130_fd_sc_hs__fa_2_1/SUM
+ sky130_fd_sc_hs__fa_2_1/a_27_378# sky130_fd_sc_hs__fa_2_1/a_701_79# sky130_fd_sc_hs__fa_2_1/a_484_347#
+ sky130_fd_sc_hs__fa_2_1/a_1094_347# sky130_fd_sc_hs__fa_2_1/a_1205_79# sky130_fd_sc_hs__fa_2_1/a_27_79#
+ sky130_fd_sc_hs__fa_2_1/a_1202_368# sky130_fd_sc_hs__fa_2_1/a_336_347# sky130_fd_sc_hs__fa_2_1/a_992_347#
+ sky130_fd_sc_hs__fa_2_1/a_1119_79# sky130_fd_sc_hs__fa_2_1/a_487_79# sky130_fd_sc_hs__fa_2_1/a_683_347#
+ sky130_fd_sc_hs__fa_2
Xsky130_fd_sc_hs__nor3_1_4 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nor3_1_5/Y sky130_fd_sc_hs__nor3_1_5/C
+ sky130_fd_sc_hs__nor3_1_5/B sky130_fd_sc_hs__nor3_1_5/A sky130_fd_sc_hs__nor3_1_5/a_198_368#
+ sky130_fd_sc_hs__nor3_1_5/a_114_368# sky130_fd_sc_hs__nor3_1
Xsky130_fd_sc_hs__xnor2_1_12 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__xnor2_1_13/A sky130_fd_sc_hs__nand4_2_1/C
+ sky130_fd_sc_hs__xnor2_1_15/Y sky130_fd_sc_hs__xnor2_1_13/a_376_368# sky130_fd_sc_hs__xnor2_1_13/a_112_119#
+ sky130_fd_sc_hs__xnor2_1_13/a_138_385# sky130_fd_sc_hs__xnor2_1_13/a_293_74# sky130_fd_sc_hs__xnor2_1
Xsky130_fd_sc_hs__a211oi_1_3 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand4_1_1/Y sky130_fd_sc_hs__nand4_1_5/C
+ sky130_fd_sc_hs__o211ai_1_5/Y sky130_fd_sc_hs__inv_4_75/Y sky130_fd_sc_hs__inv_4_85/A
+ sky130_fd_sc_hs__a211oi_1_3/a_354_368# sky130_fd_sc_hs__a211oi_1_3/a_71_368# sky130_fd_sc_hs__a211oi_1_3/a_159_74#
+ sky130_fd_sc_hs__a211oi_1
Xsky130_fd_sc_hs__a22oi_1_4 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nor2b_1_25/Y sky130_fd_sc_hs__a22oi_1_5/Y
+ sky130_fd_sc_hs__inv_4_19/A sky130_fd_sc_hs__nor2b_1_23/Y sky130_fd_sc_hs__inv_4_7/A
+ sky130_fd_sc_hs__a22oi_1_5/a_71_368# sky130_fd_sc_hs__a22oi_1_5/a_159_74# sky130_fd_sc_hs__a22oi_1_5/a_339_74#
+ sky130_fd_sc_hs__a22oi_1
Xsky130_fd_sc_hs__sdlclkp_4_1 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__conb_1_1/LO sky130_fd_sc_hs__nand2_1_23/Y
+ sky130_fd_sc_hs__o21ai_1_1/Y sky130_fd_sc_hs__dfstp_2_1/CLK sky130_fd_sc_hs__sdlclkp_4_1/a_1289_368#
+ sky130_fd_sc_hs__sdlclkp_4_1/a_744_74# sky130_fd_sc_hs__sdlclkp_4_1/a_785_455# sky130_fd_sc_hs__sdlclkp_4_1/a_634_74#
+ sky130_fd_sc_hs__sdlclkp_4_1/a_1292_74# sky130_fd_sc_hs__sdlclkp_4_1/a_792_48# sky130_fd_sc_hs__sdlclkp_4_1/a_324_79#
+ sky130_fd_sc_hs__sdlclkp_4_1/a_116_395# sky130_fd_sc_hs__sdlclkp_4_1/a_354_105#
+ sky130_fd_sc_hs__sdlclkp_4_1/a_119_143# sky130_fd_sc_hs__sdlclkp_4
Xsky130_fd_sc_hs__dfrbp_1_12 DVSS DVDD sky130_fd_sc_hs__clkbuf_8_1/X DVDD DVSS sky130_fd_sc_hs__nor2_1_59/A
+ sky130_fd_sc_hs__clkbuf_2_1/X sky130_fd_sc_hs__o21a_1_47/X sky130_fd_sc_hs__dfrbp_1_13/Q_N
+ sky130_fd_sc_hs__dfrbp_1_13/a_498_360# sky130_fd_sc_hs__dfrbp_1_13/a_1224_74# sky130_fd_sc_hs__dfrbp_1_13/a_2026_424#
+ sky130_fd_sc_hs__dfrbp_1_13/a_1482_48# sky130_fd_sc_hs__dfrbp_1_13/a_125_78# sky130_fd_sc_hs__dfrbp_1_13/a_796_463#
+ sky130_fd_sc_hs__dfrbp_1_13/a_910_118# sky130_fd_sc_hs__dfrbp_1_13/a_1465_471# sky130_fd_sc_hs__dfrbp_1_13/a_832_118#
+ sky130_fd_sc_hs__dfrbp_1_13/a_841_401# sky130_fd_sc_hs__dfrbp_1_13/a_38_78# sky130_fd_sc_hs__dfrbp_1_13/a_1434_74#
+ sky130_fd_sc_hs__dfrbp_1_13/a_706_463# sky130_fd_sc_hs__dfrbp_1_13/a_319_360# sky130_fd_sc_hs__dfrbp_1_13/a_1624_74#
+ sky130_fd_sc_hs__dfrbp_1
Xsky130_fd_sc_hs__dfrbp_1_34 DVSS DVDD sky130_fd_sc_hs__clkbuf_8_1/X DVDD DVSS sky130_fd_sc_hs__o21a_1_63/A1
+ ref_clk sky130_fd_sc_hs__o21a_1_63/X sky130_fd_sc_hs__dfrbp_1_35/Q_N sky130_fd_sc_hs__dfrbp_1_35/a_498_360#
+ sky130_fd_sc_hs__dfrbp_1_35/a_1224_74# sky130_fd_sc_hs__dfrbp_1_35/a_2026_424# sky130_fd_sc_hs__dfrbp_1_35/a_1482_48#
+ sky130_fd_sc_hs__dfrbp_1_35/a_125_78# sky130_fd_sc_hs__dfrbp_1_35/a_796_463# sky130_fd_sc_hs__dfrbp_1_35/a_910_118#
+ sky130_fd_sc_hs__dfrbp_1_35/a_1465_471# sky130_fd_sc_hs__dfrbp_1_35/a_832_118# sky130_fd_sc_hs__dfrbp_1_35/a_841_401#
+ sky130_fd_sc_hs__dfrbp_1_35/a_38_78# sky130_fd_sc_hs__dfrbp_1_35/a_1434_74# sky130_fd_sc_hs__dfrbp_1_35/a_706_463#
+ sky130_fd_sc_hs__dfrbp_1_35/a_319_360# sky130_fd_sc_hs__dfrbp_1_35/a_1624_74# sky130_fd_sc_hs__dfrbp_1
Xsky130_fd_sc_hs__dfrbp_1_45 DVSS DVDD sky130_fd_sc_hs__clkbuf_8_1/X DVDD DVSS sky130_fd_sc_hs__inv_4_113/A
+ ref_clk sky130_fd_sc_hs__o21a_1_77/X sky130_fd_sc_hs__dfrbp_1_45/Q_N sky130_fd_sc_hs__dfrbp_1_45/a_498_360#
+ sky130_fd_sc_hs__dfrbp_1_45/a_1224_74# sky130_fd_sc_hs__dfrbp_1_45/a_2026_424# sky130_fd_sc_hs__dfrbp_1_45/a_1482_48#
+ sky130_fd_sc_hs__dfrbp_1_45/a_125_78# sky130_fd_sc_hs__dfrbp_1_45/a_796_463# sky130_fd_sc_hs__dfrbp_1_45/a_910_118#
+ sky130_fd_sc_hs__dfrbp_1_45/a_1465_471# sky130_fd_sc_hs__dfrbp_1_45/a_832_118# sky130_fd_sc_hs__dfrbp_1_45/a_841_401#
+ sky130_fd_sc_hs__dfrbp_1_45/a_38_78# sky130_fd_sc_hs__dfrbp_1_45/a_1434_74# sky130_fd_sc_hs__dfrbp_1_45/a_706_463#
+ sky130_fd_sc_hs__dfrbp_1_45/a_319_360# sky130_fd_sc_hs__dfrbp_1_45/a_1624_74# sky130_fd_sc_hs__dfrbp_1
Xsky130_fd_sc_hs__dfrbp_1_23 DVSS DVDD sky130_fd_sc_hs__clkbuf_8_1/X DVDD DVSS sky130_fd_sc_hs__maj3_1_1/A
+ sky130_fd_sc_hs__clkbuf_2_1/X sky130_fd_sc_hs__o21a_1_51/X sky130_fd_sc_hs__dfrbp_1_23/Q_N
+ sky130_fd_sc_hs__dfrbp_1_23/a_498_360# sky130_fd_sc_hs__dfrbp_1_23/a_1224_74# sky130_fd_sc_hs__dfrbp_1_23/a_2026_424#
+ sky130_fd_sc_hs__dfrbp_1_23/a_1482_48# sky130_fd_sc_hs__dfrbp_1_23/a_125_78# sky130_fd_sc_hs__dfrbp_1_23/a_796_463#
+ sky130_fd_sc_hs__dfrbp_1_23/a_910_118# sky130_fd_sc_hs__dfrbp_1_23/a_1465_471# sky130_fd_sc_hs__dfrbp_1_23/a_832_118#
+ sky130_fd_sc_hs__dfrbp_1_23/a_841_401# sky130_fd_sc_hs__dfrbp_1_23/a_38_78# sky130_fd_sc_hs__dfrbp_1_23/a_1434_74#
+ sky130_fd_sc_hs__dfrbp_1_23/a_706_463# sky130_fd_sc_hs__dfrbp_1_23/a_319_360# sky130_fd_sc_hs__dfrbp_1_23/a_1624_74#
+ sky130_fd_sc_hs__dfrbp_1
Xsky130_fd_sc_hs__nand2_2_13 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_2_13/Y div_ratio_half[3]
+ sky130_fd_sc_hs__xnor2_1_3/A sky130_fd_sc_hs__nand2_2_13/a_27_74# sky130_fd_sc_hs__nand2_2
Xsky130_fd_sc_hs__xor2_1_1 DVSS DVDD DVDD DVSS fine_con_step_size[0] sky130_fd_sc_hs__fa_2_9/B
+ sky130_fd_sc_hs__xor2_1_1/X sky130_fd_sc_hs__xor2_1_1/a_194_125# sky130_fd_sc_hs__xor2_1_1/a_355_368#
+ sky130_fd_sc_hs__xor2_1_1/a_455_87# sky130_fd_sc_hs__xor2_1_1/a_158_392# sky130_fd_sc_hs__xor2_1
Xsky130_fd_sc_hs__o31ai_1_6 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nor3_1_15/Y sky130_fd_sc_hs__nor3_1_13/A
+ sky130_fd_sc_hs__nand4_1_5/D sky130_fd_sc_hs__o31ai_1_7/A1 sky130_fd_sc_hs__o31ai_1_7/Y
+ sky130_fd_sc_hs__o31ai_1_7/a_114_74# sky130_fd_sc_hs__o31ai_1_7/a_119_368# sky130_fd_sc_hs__o31ai_1_7/a_203_368#
+ sky130_fd_sc_hs__o31ai_1
Xsky130_fd_sc_hs__a21oi_1_3 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nor2_1_3/Y sky130_fd_sc_hs__dfrtp_4_3/D
+ sky130_fd_sc_hs__nor2_1_3/B sky130_fd_sc_hs__inv_4_3/Y sky130_fd_sc_hs__a21oi_1_3/a_117_74#
+ sky130_fd_sc_hs__a21oi_1_3/a_29_368# sky130_fd_sc_hs__a21oi_1
Xsky130_fd_sc_hs__dfrtn_1_35 DVSS DVDD sky130_fd_sc_hs__clkbuf_8_1/X DVDD DVSS ref_clk
+ sky130_fd_sc_hs__xnor2_1_9/A sky130_fd_sc_hs__xnor2_1_9/Y sky130_fd_sc_hs__dfrtn_1_35/a_1266_119#
+ sky130_fd_sc_hs__dfrtn_1_35/a_1736_119# sky130_fd_sc_hs__dfrtn_1_35/a_817_508# sky130_fd_sc_hs__dfrtn_1_35/a_120_74#
+ sky130_fd_sc_hs__dfrtn_1_35/a_1547_508# sky130_fd_sc_hs__dfrtn_1_35/a_922_127# sky130_fd_sc_hs__dfrtn_1_35/a_33_74#
+ sky130_fd_sc_hs__dfrtn_1_35/a_714_127# sky130_fd_sc_hs__dfrtn_1_35/a_1934_94# sky130_fd_sc_hs__dfrtn_1_35/a_1550_119#
+ sky130_fd_sc_hs__dfrtn_1_35/a_1598_93# sky130_fd_sc_hs__dfrtn_1_35/a_300_74# sky130_fd_sc_hs__dfrtn_1_35/a_507_368#
+ sky130_fd_sc_hs__dfrtn_1_35/a_856_304# sky130_fd_sc_hs__dfrtn_1_35/a_850_127# sky130_fd_sc_hs__dfrtn_1
Xsky130_fd_sc_hs__nand2_1_108 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_137/Y sky130_fd_sc_hs__nand4_1_1/C
+ sky130_fd_sc_hs__inv_4_129/A sky130_fd_sc_hs__nand2_1_109/a_117_74# sky130_fd_sc_hs__nand2_1
Xsky130_fd_sc_hs__dfrtn_1_24 DVSS DVDD sky130_fd_sc_hs__clkbuf_8_1/X DVDD DVSS ref_clk
+ sky130_fd_sc_hs__inv_4_97/A sky130_fd_sc_hs__o21a_1_55/X sky130_fd_sc_hs__dfrtn_1_25/a_1266_119#
+ sky130_fd_sc_hs__dfrtn_1_25/a_1736_119# sky130_fd_sc_hs__dfrtn_1_25/a_817_508# sky130_fd_sc_hs__dfrtn_1_25/a_120_74#
+ sky130_fd_sc_hs__dfrtn_1_25/a_1547_508# sky130_fd_sc_hs__dfrtn_1_25/a_922_127# sky130_fd_sc_hs__dfrtn_1_25/a_33_74#
+ sky130_fd_sc_hs__dfrtn_1_25/a_714_127# sky130_fd_sc_hs__dfrtn_1_25/a_1934_94# sky130_fd_sc_hs__dfrtn_1_25/a_1550_119#
+ sky130_fd_sc_hs__dfrtn_1_25/a_1598_93# sky130_fd_sc_hs__dfrtn_1_25/a_300_74# sky130_fd_sc_hs__dfrtn_1_25/a_507_368#
+ sky130_fd_sc_hs__dfrtn_1_25/a_856_304# sky130_fd_sc_hs__dfrtn_1_25/a_850_127# sky130_fd_sc_hs__dfrtn_1
Xsky130_fd_sc_hs__dfrtn_1_13 DVSS DVDD sky130_fd_sc_hs__clkbuf_8_1/X DVDD DVSS sky130_fd_sc_hs__clkbuf_2_1/X
+ sky130_fd_sc_hs__inv_4_59/A sky130_fd_sc_hs__dfrtn_1_13/D sky130_fd_sc_hs__dfrtn_1_13/a_1266_119#
+ sky130_fd_sc_hs__dfrtn_1_13/a_1736_119# sky130_fd_sc_hs__dfrtn_1_13/a_817_508# sky130_fd_sc_hs__dfrtn_1_13/a_120_74#
+ sky130_fd_sc_hs__dfrtn_1_13/a_1547_508# sky130_fd_sc_hs__dfrtn_1_13/a_922_127# sky130_fd_sc_hs__dfrtn_1_13/a_33_74#
+ sky130_fd_sc_hs__dfrtn_1_13/a_714_127# sky130_fd_sc_hs__dfrtn_1_13/a_1934_94# sky130_fd_sc_hs__dfrtn_1_13/a_1550_119#
+ sky130_fd_sc_hs__dfrtn_1_13/a_1598_93# sky130_fd_sc_hs__dfrtn_1_13/a_300_74# sky130_fd_sc_hs__dfrtn_1_13/a_507_368#
+ sky130_fd_sc_hs__dfrtn_1_13/a_856_304# sky130_fd_sc_hs__dfrtn_1_13/a_850_127# sky130_fd_sc_hs__dfrtn_1
Xsky130_fd_sc_hs__dfrtn_1_46 DVSS DVDD sky130_fd_sc_hs__clkbuf_8_1/X DVDD DVSS ref_clk
+ sky130_fd_sc_hs__inv_4_127/A sky130_fd_sc_hs__o21a_1_69/X sky130_fd_sc_hs__dfrtn_1_47/a_1266_119#
+ sky130_fd_sc_hs__dfrtn_1_47/a_1736_119# sky130_fd_sc_hs__dfrtn_1_47/a_817_508# sky130_fd_sc_hs__dfrtn_1_47/a_120_74#
+ sky130_fd_sc_hs__dfrtn_1_47/a_1547_508# sky130_fd_sc_hs__dfrtn_1_47/a_922_127# sky130_fd_sc_hs__dfrtn_1_47/a_33_74#
+ sky130_fd_sc_hs__dfrtn_1_47/a_714_127# sky130_fd_sc_hs__dfrtn_1_47/a_1934_94# sky130_fd_sc_hs__dfrtn_1_47/a_1550_119#
+ sky130_fd_sc_hs__dfrtn_1_47/a_1598_93# sky130_fd_sc_hs__dfrtn_1_47/a_300_74# sky130_fd_sc_hs__dfrtn_1_47/a_507_368#
+ sky130_fd_sc_hs__dfrtn_1_47/a_856_304# sky130_fd_sc_hs__dfrtn_1_47/a_850_127# sky130_fd_sc_hs__dfrtn_1
Xsky130_fd_sc_hs__nand2_1_119 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__o21a_1_75/A2 sky130_fd_sc_hs__o21a_1_75/B1
+ sky130_fd_sc_hs__o21a_1_75/A1 sky130_fd_sc_hs__nand2_1_119/a_117_74# sky130_fd_sc_hs__nand2_1
Xsky130_fd_sc_hs__dfrbp_1_1 DVSS DVDD sky130_fd_sc_hs__clkbuf_8_1/X DVDD DVSS sky130_fd_sc_hs__dfrbp_1_1/Q
+ sky130_fd_sc_hs__clkbuf_2_1/X sky130_fd_sc_hs__o21a_1_35/X sky130_fd_sc_hs__dfrbp_1_1/Q_N
+ sky130_fd_sc_hs__dfrbp_1_1/a_498_360# sky130_fd_sc_hs__dfrbp_1_1/a_1224_74# sky130_fd_sc_hs__dfrbp_1_1/a_2026_424#
+ sky130_fd_sc_hs__dfrbp_1_1/a_1482_48# sky130_fd_sc_hs__dfrbp_1_1/a_125_78# sky130_fd_sc_hs__dfrbp_1_1/a_796_463#
+ sky130_fd_sc_hs__dfrbp_1_1/a_910_118# sky130_fd_sc_hs__dfrbp_1_1/a_1465_471# sky130_fd_sc_hs__dfrbp_1_1/a_832_118#
+ sky130_fd_sc_hs__dfrbp_1_1/a_841_401# sky130_fd_sc_hs__dfrbp_1_1/a_38_78# sky130_fd_sc_hs__dfrbp_1_1/a_1434_74#
+ sky130_fd_sc_hs__dfrbp_1_1/a_706_463# sky130_fd_sc_hs__dfrbp_1_1/a_319_360# sky130_fd_sc_hs__dfrbp_1_1/a_1624_74#
+ sky130_fd_sc_hs__dfrbp_1
Xsky130_fd_sc_hs__dfstp_2_6 DVSS DVDD sky130_fd_sc_hs__inv_4_49/Y DVDD DVSS sky130_fd_sc_hs__o21ai_1_1/Y
+ sky130_fd_sc_hs__dfstp_2_7/D sky130_fd_sc_hs__dfstp_2_7/Q sky130_fd_sc_hs__dfstp_2_7/a_1566_92#
+ sky130_fd_sc_hs__dfstp_2_7/a_1521_508# sky130_fd_sc_hs__dfstp_2_7/a_716_456# sky130_fd_sc_hs__dfstp_2_7/a_1266_341#
+ sky130_fd_sc_hs__dfstp_2_7/a_1278_74# sky130_fd_sc_hs__dfstp_2_7/a_398_74# sky130_fd_sc_hs__dfstp_2_7/a_1057_118#
+ sky130_fd_sc_hs__dfstp_2_7/a_1489_118# sky130_fd_sc_hs__dfstp_2_7/a_27_74# sky130_fd_sc_hs__dfstp_2_7/a_1596_118#
+ sky130_fd_sc_hs__dfstp_2_7/a_225_74# sky130_fd_sc_hs__dfstp_2_7/a_1356_74# sky130_fd_sc_hs__dfstp_2_7/a_612_74#
+ sky130_fd_sc_hs__dfstp_2_7/a_781_74# sky130_fd_sc_hs__dfstp_2_7/a_767_384# sky130_fd_sc_hs__dfstp_2_7/a_2022_94#
+ sky130_fd_sc_hs__dfstp_2
Xsky130_fd_sc_hs__dfrtp_4_8 DVSS DVDD sky130_fd_sc_hs__clkbuf_8_1/X DVDD DVSS sky130_fd_sc_hs__o21a_1_1/X
+ sky130_fd_sc_hs__nand2_1_47/B sky130_fd_sc_hs__o21a_1_1/A1 sky130_fd_sc_hs__dfrtp_4_9/a_37_78#
+ sky130_fd_sc_hs__dfrtp_4_9/a_494_366# sky130_fd_sc_hs__dfrtp_4_9/a_699_463# sky130_fd_sc_hs__dfrtp_4_9/a_313_74#
+ sky130_fd_sc_hs__dfrtp_4_9/a_1627_493# sky130_fd_sc_hs__dfrtp_4_9/a_1678_395# sky130_fd_sc_hs__dfrtp_4_9/a_1827_81#
+ sky130_fd_sc_hs__dfrtp_4_9/a_789_463# sky130_fd_sc_hs__dfrtp_4_9/a_1350_392# sky130_fd_sc_hs__dfrtp_4_9/a_834_355#
+ sky130_fd_sc_hs__dfrtp_4_9/a_812_138# sky130_fd_sc_hs__dfrtp_4_9/a_124_78# sky130_fd_sc_hs__dfrtp_4_9/a_1647_81#
+ sky130_fd_sc_hs__dfrtp_4_9/a_2010_409# sky130_fd_sc_hs__dfrtp_4_9/a_890_138# sky130_fd_sc_hs__dfrtp_4
Xsky130_fd_sc_hs__inv_4_35 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_35/Y sky130_fd_sc_hs__inv_4_35/A
+ sky130_fd_sc_hs__inv_4
Xsky130_fd_sc_hs__inv_4_24 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_25/Y sky130_fd_sc_hs__inv_4_25/A
+ sky130_fd_sc_hs__inv_4
Xsky130_fd_sc_hs__inv_4_13 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_13/Y sky130_fd_sc_hs__inv_4_13/A
+ sky130_fd_sc_hs__inv_4
Xsky130_fd_sc_hs__inv_4_68 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_69/Y sky130_fd_sc_hs__inv_4_69/A
+ sky130_fd_sc_hs__inv_4
Xsky130_fd_sc_hs__inv_4_57 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_57/Y out_star
+ sky130_fd_sc_hs__inv_4
Xsky130_fd_sc_hs__inv_4_46 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_47/Y sky130_fd_sc_hs__inv_4_47/A
+ sky130_fd_sc_hs__inv_4
Xsky130_fd_sc_hs__inv_4_79 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_79/Y sky130_fd_sc_hs__inv_4_79/A
+ sky130_fd_sc_hs__inv_4
Xsky130_fd_sc_hs__fa_2_1 DVSS DVDD sky130_fd_sc_hs__fa_2_1/A DVDD DVSS sky130_fd_sc_hs__fa_2_1/CIN
+ sky130_fd_sc_hs__fa_2_1/B sky130_fd_sc_hs__fa_2_7/CIN sky130_fd_sc_hs__fa_2_1/SUM
+ sky130_fd_sc_hs__fa_2_1/a_27_378# sky130_fd_sc_hs__fa_2_1/a_701_79# sky130_fd_sc_hs__fa_2_1/a_484_347#
+ sky130_fd_sc_hs__fa_2_1/a_1094_347# sky130_fd_sc_hs__fa_2_1/a_1205_79# sky130_fd_sc_hs__fa_2_1/a_27_79#
+ sky130_fd_sc_hs__fa_2_1/a_1202_368# sky130_fd_sc_hs__fa_2_1/a_336_347# sky130_fd_sc_hs__fa_2_1/a_992_347#
+ sky130_fd_sc_hs__fa_2_1/a_1119_79# sky130_fd_sc_hs__fa_2_1/a_487_79# sky130_fd_sc_hs__fa_2_1/a_683_347#
+ sky130_fd_sc_hs__fa_2
Xsky130_fd_sc_hs__nor3_1_5 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nor3_1_5/Y sky130_fd_sc_hs__nor3_1_5/C
+ sky130_fd_sc_hs__nor3_1_5/B sky130_fd_sc_hs__nor3_1_5/A sky130_fd_sc_hs__nor3_1_5/a_198_368#
+ sky130_fd_sc_hs__nor3_1_5/a_114_368# sky130_fd_sc_hs__nor3_1
Xsky130_fd_sc_hs__xnor2_1_13 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__xnor2_1_13/A sky130_fd_sc_hs__nand4_2_1/C
+ sky130_fd_sc_hs__xnor2_1_15/Y sky130_fd_sc_hs__xnor2_1_13/a_376_368# sky130_fd_sc_hs__xnor2_1_13/a_112_119#
+ sky130_fd_sc_hs__xnor2_1_13/a_138_385# sky130_fd_sc_hs__xnor2_1_13/a_293_74# sky130_fd_sc_hs__xnor2_1
Xsky130_fd_sc_hs__a22oi_1_5 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nor2b_1_25/Y sky130_fd_sc_hs__a22oi_1_5/Y
+ sky130_fd_sc_hs__inv_4_19/A sky130_fd_sc_hs__nor2b_1_23/Y sky130_fd_sc_hs__inv_4_7/A
+ sky130_fd_sc_hs__a22oi_1_5/a_71_368# sky130_fd_sc_hs__a22oi_1_5/a_159_74# sky130_fd_sc_hs__a22oi_1_5/a_339_74#
+ sky130_fd_sc_hs__a22oi_1
Xsky130_fd_sc_hs__a21oi_1_90 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__o22ai_1_9/B1 sky130_fd_sc_hs__a21oi_1_91/Y
+ sky130_fd_sc_hs__maj3_1_1/C sky130_fd_sc_hs__maj3_1_1/A sky130_fd_sc_hs__a21oi_1_91/a_117_74#
+ sky130_fd_sc_hs__a21oi_1_91/a_29_368# sky130_fd_sc_hs__a21oi_1
Xsky130_fd_sc_hs__dfrbp_1_35 DVSS DVDD sky130_fd_sc_hs__clkbuf_8_1/X DVDD DVSS sky130_fd_sc_hs__o21a_1_63/A1
+ ref_clk sky130_fd_sc_hs__o21a_1_63/X sky130_fd_sc_hs__dfrbp_1_35/Q_N sky130_fd_sc_hs__dfrbp_1_35/a_498_360#
+ sky130_fd_sc_hs__dfrbp_1_35/a_1224_74# sky130_fd_sc_hs__dfrbp_1_35/a_2026_424# sky130_fd_sc_hs__dfrbp_1_35/a_1482_48#
+ sky130_fd_sc_hs__dfrbp_1_35/a_125_78# sky130_fd_sc_hs__dfrbp_1_35/a_796_463# sky130_fd_sc_hs__dfrbp_1_35/a_910_118#
+ sky130_fd_sc_hs__dfrbp_1_35/a_1465_471# sky130_fd_sc_hs__dfrbp_1_35/a_832_118# sky130_fd_sc_hs__dfrbp_1_35/a_841_401#
+ sky130_fd_sc_hs__dfrbp_1_35/a_38_78# sky130_fd_sc_hs__dfrbp_1_35/a_1434_74# sky130_fd_sc_hs__dfrbp_1_35/a_706_463#
+ sky130_fd_sc_hs__dfrbp_1_35/a_319_360# sky130_fd_sc_hs__dfrbp_1_35/a_1624_74# sky130_fd_sc_hs__dfrbp_1
Xsky130_fd_sc_hs__dfrbp_1_46 DVSS DVDD sky130_fd_sc_hs__clkbuf_8_1/X DVDD DVSS sky130_fd_sc_hs__or2_1_3/A
+ ref_clk sky130_fd_sc_hs__o21a_1_73/X sky130_fd_sc_hs__dfrbp_1_47/Q_N sky130_fd_sc_hs__dfrbp_1_47/a_498_360#
+ sky130_fd_sc_hs__dfrbp_1_47/a_1224_74# sky130_fd_sc_hs__dfrbp_1_47/a_2026_424# sky130_fd_sc_hs__dfrbp_1_47/a_1482_48#
+ sky130_fd_sc_hs__dfrbp_1_47/a_125_78# sky130_fd_sc_hs__dfrbp_1_47/a_796_463# sky130_fd_sc_hs__dfrbp_1_47/a_910_118#
+ sky130_fd_sc_hs__dfrbp_1_47/a_1465_471# sky130_fd_sc_hs__dfrbp_1_47/a_832_118# sky130_fd_sc_hs__dfrbp_1_47/a_841_401#
+ sky130_fd_sc_hs__dfrbp_1_47/a_38_78# sky130_fd_sc_hs__dfrbp_1_47/a_1434_74# sky130_fd_sc_hs__dfrbp_1_47/a_706_463#
+ sky130_fd_sc_hs__dfrbp_1_47/a_319_360# sky130_fd_sc_hs__dfrbp_1_47/a_1624_74# sky130_fd_sc_hs__dfrbp_1
Xsky130_fd_sc_hs__dfrbp_1_24 DVSS DVDD sky130_fd_sc_hs__clkbuf_8_1/X DVDD DVSS sky130_fd_sc_hs__o22ai_1_7/A1
+ sky130_fd_sc_hs__clkbuf_2_1/X sky130_fd_sc_hs__o21a_1_53/X sky130_fd_sc_hs__dfrbp_1_25/Q_N
+ sky130_fd_sc_hs__dfrbp_1_25/a_498_360# sky130_fd_sc_hs__dfrbp_1_25/a_1224_74# sky130_fd_sc_hs__dfrbp_1_25/a_2026_424#
+ sky130_fd_sc_hs__dfrbp_1_25/a_1482_48# sky130_fd_sc_hs__dfrbp_1_25/a_125_78# sky130_fd_sc_hs__dfrbp_1_25/a_796_463#
+ sky130_fd_sc_hs__dfrbp_1_25/a_910_118# sky130_fd_sc_hs__dfrbp_1_25/a_1465_471# sky130_fd_sc_hs__dfrbp_1_25/a_832_118#
+ sky130_fd_sc_hs__dfrbp_1_25/a_841_401# sky130_fd_sc_hs__dfrbp_1_25/a_38_78# sky130_fd_sc_hs__dfrbp_1_25/a_1434_74#
+ sky130_fd_sc_hs__dfrbp_1_25/a_706_463# sky130_fd_sc_hs__dfrbp_1_25/a_319_360# sky130_fd_sc_hs__dfrbp_1_25/a_1624_74#
+ sky130_fd_sc_hs__dfrbp_1
Xsky130_fd_sc_hs__dfrbp_1_13 DVSS DVDD sky130_fd_sc_hs__clkbuf_8_1/X DVDD DVSS sky130_fd_sc_hs__nor2_1_59/A
+ sky130_fd_sc_hs__clkbuf_2_1/X sky130_fd_sc_hs__o21a_1_47/X sky130_fd_sc_hs__dfrbp_1_13/Q_N
+ sky130_fd_sc_hs__dfrbp_1_13/a_498_360# sky130_fd_sc_hs__dfrbp_1_13/a_1224_74# sky130_fd_sc_hs__dfrbp_1_13/a_2026_424#
+ sky130_fd_sc_hs__dfrbp_1_13/a_1482_48# sky130_fd_sc_hs__dfrbp_1_13/a_125_78# sky130_fd_sc_hs__dfrbp_1_13/a_796_463#
+ sky130_fd_sc_hs__dfrbp_1_13/a_910_118# sky130_fd_sc_hs__dfrbp_1_13/a_1465_471# sky130_fd_sc_hs__dfrbp_1_13/a_832_118#
+ sky130_fd_sc_hs__dfrbp_1_13/a_841_401# sky130_fd_sc_hs__dfrbp_1_13/a_38_78# sky130_fd_sc_hs__dfrbp_1_13/a_1434_74#
+ sky130_fd_sc_hs__dfrbp_1_13/a_706_463# sky130_fd_sc_hs__dfrbp_1_13/a_319_360# sky130_fd_sc_hs__dfrbp_1_13/a_1624_74#
+ sky130_fd_sc_hs__dfrbp_1
Xsky130_fd_sc_hs__nand2_2_14 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand3_1_1/C div_ratio_half[3]
+ sky130_fd_sc_hs__xnor2_1_3/A sky130_fd_sc_hs__nand2_2_15/a_27_74# sky130_fd_sc_hs__nand2_2
Xsky130_fd_sc_hs__xor2_1_2 DVSS DVDD DVDD DVSS fine_con_step_size[1] sky130_fd_sc_hs__fa_2_9/B
+ sky130_fd_sc_hs__fa_2_5/A sky130_fd_sc_hs__xor2_1_3/a_194_125# sky130_fd_sc_hs__xor2_1_3/a_355_368#
+ sky130_fd_sc_hs__xor2_1_3/a_455_87# sky130_fd_sc_hs__xor2_1_3/a_158_392# sky130_fd_sc_hs__xor2_1
Xsky130_fd_sc_hs__o31ai_1_7 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nor3_1_15/Y sky130_fd_sc_hs__nor3_1_13/A
+ sky130_fd_sc_hs__nand4_1_5/D sky130_fd_sc_hs__o31ai_1_7/A1 sky130_fd_sc_hs__o31ai_1_7/Y
+ sky130_fd_sc_hs__o31ai_1_7/a_114_74# sky130_fd_sc_hs__o31ai_1_7/a_119_368# sky130_fd_sc_hs__o31ai_1_7/a_203_368#
+ sky130_fd_sc_hs__o31ai_1
Xsky130_fd_sc_hs__a21oi_1_4 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nor2_1_5/Y sky130_fd_sc_hs__dfrtp_4_5/D
+ sky130_fd_sc_hs__nor2_1_5/B sky130_fd_sc_hs__inv_4_7/Y sky130_fd_sc_hs__a21oi_1_5/a_117_74#
+ sky130_fd_sc_hs__a21oi_1_5/a_29_368# sky130_fd_sc_hs__a21oi_1
Xsky130_fd_sc_hs__dfrtn_1_36 DVSS DVDD sky130_fd_sc_hs__clkbuf_8_1/X DVDD DVSS ref_clk
+ sky130_fd_sc_hs__inv_4_111/A sky130_fd_sc_hs__dfrtn_1_37/D sky130_fd_sc_hs__dfrtn_1_37/a_1266_119#
+ sky130_fd_sc_hs__dfrtn_1_37/a_1736_119# sky130_fd_sc_hs__dfrtn_1_37/a_817_508# sky130_fd_sc_hs__dfrtn_1_37/a_120_74#
+ sky130_fd_sc_hs__dfrtn_1_37/a_1547_508# sky130_fd_sc_hs__dfrtn_1_37/a_922_127# sky130_fd_sc_hs__dfrtn_1_37/a_33_74#
+ sky130_fd_sc_hs__dfrtn_1_37/a_714_127# sky130_fd_sc_hs__dfrtn_1_37/a_1934_94# sky130_fd_sc_hs__dfrtn_1_37/a_1550_119#
+ sky130_fd_sc_hs__dfrtn_1_37/a_1598_93# sky130_fd_sc_hs__dfrtn_1_37/a_300_74# sky130_fd_sc_hs__dfrtn_1_37/a_507_368#
+ sky130_fd_sc_hs__dfrtn_1_37/a_856_304# sky130_fd_sc_hs__dfrtn_1_37/a_850_127# sky130_fd_sc_hs__dfrtn_1
Xsky130_fd_sc_hs__dfrtn_1_25 DVSS DVDD sky130_fd_sc_hs__clkbuf_8_1/X DVDD DVSS ref_clk
+ sky130_fd_sc_hs__inv_4_97/A sky130_fd_sc_hs__o21a_1_55/X sky130_fd_sc_hs__dfrtn_1_25/a_1266_119#
+ sky130_fd_sc_hs__dfrtn_1_25/a_1736_119# sky130_fd_sc_hs__dfrtn_1_25/a_817_508# sky130_fd_sc_hs__dfrtn_1_25/a_120_74#
+ sky130_fd_sc_hs__dfrtn_1_25/a_1547_508# sky130_fd_sc_hs__dfrtn_1_25/a_922_127# sky130_fd_sc_hs__dfrtn_1_25/a_33_74#
+ sky130_fd_sc_hs__dfrtn_1_25/a_714_127# sky130_fd_sc_hs__dfrtn_1_25/a_1934_94# sky130_fd_sc_hs__dfrtn_1_25/a_1550_119#
+ sky130_fd_sc_hs__dfrtn_1_25/a_1598_93# sky130_fd_sc_hs__dfrtn_1_25/a_300_74# sky130_fd_sc_hs__dfrtn_1_25/a_507_368#
+ sky130_fd_sc_hs__dfrtn_1_25/a_856_304# sky130_fd_sc_hs__dfrtn_1_25/a_850_127# sky130_fd_sc_hs__dfrtn_1
Xsky130_fd_sc_hs__dfrtn_1_14 DVSS DVDD sky130_fd_sc_hs__clkbuf_8_1/X DVDD DVSS sky130_fd_sc_hs__clkbuf_2_1/X
+ sky130_fd_sc_hs__inv_4_65/A sky130_fd_sc_hs__dfrtn_1_15/D sky130_fd_sc_hs__dfrtn_1_15/a_1266_119#
+ sky130_fd_sc_hs__dfrtn_1_15/a_1736_119# sky130_fd_sc_hs__dfrtn_1_15/a_817_508# sky130_fd_sc_hs__dfrtn_1_15/a_120_74#
+ sky130_fd_sc_hs__dfrtn_1_15/a_1547_508# sky130_fd_sc_hs__dfrtn_1_15/a_922_127# sky130_fd_sc_hs__dfrtn_1_15/a_33_74#
+ sky130_fd_sc_hs__dfrtn_1_15/a_714_127# sky130_fd_sc_hs__dfrtn_1_15/a_1934_94# sky130_fd_sc_hs__dfrtn_1_15/a_1550_119#
+ sky130_fd_sc_hs__dfrtn_1_15/a_1598_93# sky130_fd_sc_hs__dfrtn_1_15/a_300_74# sky130_fd_sc_hs__dfrtn_1_15/a_507_368#
+ sky130_fd_sc_hs__dfrtn_1_15/a_856_304# sky130_fd_sc_hs__dfrtn_1_15/a_850_127# sky130_fd_sc_hs__dfrtn_1
Xsky130_fd_sc_hs__nand2_1_109 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_137/Y sky130_fd_sc_hs__nand4_1_1/C
+ sky130_fd_sc_hs__inv_4_129/A sky130_fd_sc_hs__nand2_1_109/a_117_74# sky130_fd_sc_hs__nand2_1
Xsky130_fd_sc_hs__dfrtn_1_47 DVSS DVDD sky130_fd_sc_hs__clkbuf_8_1/X DVDD DVSS ref_clk
+ sky130_fd_sc_hs__inv_4_127/A sky130_fd_sc_hs__o21a_1_69/X sky130_fd_sc_hs__dfrtn_1_47/a_1266_119#
+ sky130_fd_sc_hs__dfrtn_1_47/a_1736_119# sky130_fd_sc_hs__dfrtn_1_47/a_817_508# sky130_fd_sc_hs__dfrtn_1_47/a_120_74#
+ sky130_fd_sc_hs__dfrtn_1_47/a_1547_508# sky130_fd_sc_hs__dfrtn_1_47/a_922_127# sky130_fd_sc_hs__dfrtn_1_47/a_33_74#
+ sky130_fd_sc_hs__dfrtn_1_47/a_714_127# sky130_fd_sc_hs__dfrtn_1_47/a_1934_94# sky130_fd_sc_hs__dfrtn_1_47/a_1550_119#
+ sky130_fd_sc_hs__dfrtn_1_47/a_1598_93# sky130_fd_sc_hs__dfrtn_1_47/a_300_74# sky130_fd_sc_hs__dfrtn_1_47/a_507_368#
+ sky130_fd_sc_hs__dfrtn_1_47/a_856_304# sky130_fd_sc_hs__dfrtn_1_47/a_850_127# sky130_fd_sc_hs__dfrtn_1
Xsky130_fd_sc_hs__nand2b_1_0 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_1_47/B sky130_fd_sc_hs__nor2b_1_33/Y
+ sky130_fd_sc_hs__nor2_1_73/B sky130_fd_sc_hs__nand2b_1_1/a_269_74# sky130_fd_sc_hs__nand2b_1_1/a_27_112#
+ sky130_fd_sc_hs__nand2b_1
Xsky130_fd_sc_hs__dfrbp_1_2 DVSS DVDD sky130_fd_sc_hs__clkbuf_8_1/X DVDD DVSS sky130_fd_sc_hs__inv_4_61/A
+ sky130_fd_sc_hs__clkbuf_2_1/X sky130_fd_sc_hs__dfrbp_1_3/D sky130_fd_sc_hs__dfrbp_1_3/Q_N
+ sky130_fd_sc_hs__dfrbp_1_3/a_498_360# sky130_fd_sc_hs__dfrbp_1_3/a_1224_74# sky130_fd_sc_hs__dfrbp_1_3/a_2026_424#
+ sky130_fd_sc_hs__dfrbp_1_3/a_1482_48# sky130_fd_sc_hs__dfrbp_1_3/a_125_78# sky130_fd_sc_hs__dfrbp_1_3/a_796_463#
+ sky130_fd_sc_hs__dfrbp_1_3/a_910_118# sky130_fd_sc_hs__dfrbp_1_3/a_1465_471# sky130_fd_sc_hs__dfrbp_1_3/a_832_118#
+ sky130_fd_sc_hs__dfrbp_1_3/a_841_401# sky130_fd_sc_hs__dfrbp_1_3/a_38_78# sky130_fd_sc_hs__dfrbp_1_3/a_1434_74#
+ sky130_fd_sc_hs__dfrbp_1_3/a_706_463# sky130_fd_sc_hs__dfrbp_1_3/a_319_360# sky130_fd_sc_hs__dfrbp_1_3/a_1624_74#
+ sky130_fd_sc_hs__dfrbp_1
Xsky130_fd_sc_hs__dfrtn_1_0 DVSS DVDD sky130_fd_sc_hs__clkbuf_8_1/X DVDD DVSS sky130_fd_sc_hs__clkbuf_2_1/X
+ sky130_fd_sc_hs__inv_4_39/A sky130_fd_sc_hs__o21a_1_29/X sky130_fd_sc_hs__dfrtn_1_1/a_1266_119#
+ sky130_fd_sc_hs__dfrtn_1_1/a_1736_119# sky130_fd_sc_hs__dfrtn_1_1/a_817_508# sky130_fd_sc_hs__dfrtn_1_1/a_120_74#
+ sky130_fd_sc_hs__dfrtn_1_1/a_1547_508# sky130_fd_sc_hs__dfrtn_1_1/a_922_127# sky130_fd_sc_hs__dfrtn_1_1/a_33_74#
+ sky130_fd_sc_hs__dfrtn_1_1/a_714_127# sky130_fd_sc_hs__dfrtn_1_1/a_1934_94# sky130_fd_sc_hs__dfrtn_1_1/a_1550_119#
+ sky130_fd_sc_hs__dfrtn_1_1/a_1598_93# sky130_fd_sc_hs__dfrtn_1_1/a_300_74# sky130_fd_sc_hs__dfrtn_1_1/a_507_368#
+ sky130_fd_sc_hs__dfrtn_1_1/a_856_304# sky130_fd_sc_hs__dfrtn_1_1/a_850_127# sky130_fd_sc_hs__dfrtn_1
Xsky130_fd_sc_hs__dfstp_2_7 DVSS DVDD sky130_fd_sc_hs__inv_4_49/Y DVDD DVSS sky130_fd_sc_hs__o21ai_1_1/Y
+ sky130_fd_sc_hs__dfstp_2_7/D sky130_fd_sc_hs__dfstp_2_7/Q sky130_fd_sc_hs__dfstp_2_7/a_1566_92#
+ sky130_fd_sc_hs__dfstp_2_7/a_1521_508# sky130_fd_sc_hs__dfstp_2_7/a_716_456# sky130_fd_sc_hs__dfstp_2_7/a_1266_341#
+ sky130_fd_sc_hs__dfstp_2_7/a_1278_74# sky130_fd_sc_hs__dfstp_2_7/a_398_74# sky130_fd_sc_hs__dfstp_2_7/a_1057_118#
+ sky130_fd_sc_hs__dfstp_2_7/a_1489_118# sky130_fd_sc_hs__dfstp_2_7/a_27_74# sky130_fd_sc_hs__dfstp_2_7/a_1596_118#
+ sky130_fd_sc_hs__dfstp_2_7/a_225_74# sky130_fd_sc_hs__dfstp_2_7/a_1356_74# sky130_fd_sc_hs__dfstp_2_7/a_612_74#
+ sky130_fd_sc_hs__dfstp_2_7/a_781_74# sky130_fd_sc_hs__dfstp_2_7/a_767_384# sky130_fd_sc_hs__dfstp_2_7/a_2022_94#
+ sky130_fd_sc_hs__dfstp_2
Xsky130_fd_sc_hs__dfrtp_4_9 DVSS DVDD sky130_fd_sc_hs__clkbuf_8_1/X DVDD DVSS sky130_fd_sc_hs__o21a_1_1/X
+ sky130_fd_sc_hs__nand2_1_47/B sky130_fd_sc_hs__o21a_1_1/A1 sky130_fd_sc_hs__dfrtp_4_9/a_37_78#
+ sky130_fd_sc_hs__dfrtp_4_9/a_494_366# sky130_fd_sc_hs__dfrtp_4_9/a_699_463# sky130_fd_sc_hs__dfrtp_4_9/a_313_74#
+ sky130_fd_sc_hs__dfrtp_4_9/a_1627_493# sky130_fd_sc_hs__dfrtp_4_9/a_1678_395# sky130_fd_sc_hs__dfrtp_4_9/a_1827_81#
+ sky130_fd_sc_hs__dfrtp_4_9/a_789_463# sky130_fd_sc_hs__dfrtp_4_9/a_1350_392# sky130_fd_sc_hs__dfrtp_4_9/a_834_355#
+ sky130_fd_sc_hs__dfrtp_4_9/a_812_138# sky130_fd_sc_hs__dfrtp_4_9/a_124_78# sky130_fd_sc_hs__dfrtp_4_9/a_1647_81#
+ sky130_fd_sc_hs__dfrtp_4_9/a_2010_409# sky130_fd_sc_hs__dfrtp_4_9/a_890_138# sky130_fd_sc_hs__dfrtp_4
Xsky130_fd_sc_hs__o211ai_1_0 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__a21oi_1_91/Y sky130_fd_sc_hs__nor2_1_61/B
+ sky130_fd_sc_hs__nand2_1_67/Y sky130_fd_sc_hs__inv_4_79/Y sky130_fd_sc_hs__inv_4_59/A
+ sky130_fd_sc_hs__o211ai_1_1/a_31_74# sky130_fd_sc_hs__o211ai_1_1/a_311_74# sky130_fd_sc_hs__o211ai_1_1/a_116_368#
+ sky130_fd_sc_hs__o211ai_1
Xsky130_fd_sc_hs__inv_4_36 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_37/Y sky130_fd_sc_hs__inv_4_37/A
+ sky130_fd_sc_hs__inv_4
Xsky130_fd_sc_hs__inv_4_25 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_25/Y sky130_fd_sc_hs__inv_4_25/A
+ sky130_fd_sc_hs__inv_4
Xsky130_fd_sc_hs__inv_4_14 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_15/Y sky130_fd_sc_hs__inv_4_15/A
+ sky130_fd_sc_hs__inv_4
Xsky130_fd_sc_hs__inv_4_69 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_69/Y sky130_fd_sc_hs__inv_4_69/A
+ sky130_fd_sc_hs__inv_4
Xsky130_fd_sc_hs__inv_4_58 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_59/Y sky130_fd_sc_hs__inv_4_59/A
+ sky130_fd_sc_hs__inv_4
Xsky130_fd_sc_hs__inv_4_47 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_47/Y sky130_fd_sc_hs__inv_4_47/A
+ sky130_fd_sc_hs__inv_4
Xsky130_fd_sc_hs__fa_2_2 DVSS DVDD sky130_fd_sc_hs__fa_2_3/A DVDD DVSS sky130_fd_sc_hs__fa_2_3/CIN
+ sky130_fd_sc_hs__fa_2_3/B sky130_fd_sc_hs__fa_2_1/CIN sky130_fd_sc_hs__fa_2_3/SUM
+ sky130_fd_sc_hs__fa_2_3/a_27_378# sky130_fd_sc_hs__fa_2_3/a_701_79# sky130_fd_sc_hs__fa_2_3/a_484_347#
+ sky130_fd_sc_hs__fa_2_3/a_1094_347# sky130_fd_sc_hs__fa_2_3/a_1205_79# sky130_fd_sc_hs__fa_2_3/a_27_79#
+ sky130_fd_sc_hs__fa_2_3/a_1202_368# sky130_fd_sc_hs__fa_2_3/a_336_347# sky130_fd_sc_hs__fa_2_3/a_992_347#
+ sky130_fd_sc_hs__fa_2_3/a_1119_79# sky130_fd_sc_hs__fa_2_3/a_487_79# sky130_fd_sc_hs__fa_2_3/a_683_347#
+ sky130_fd_sc_hs__fa_2
Xsky130_fd_sc_hs__nor3_1_6 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nor3_1_7/Y sky130_fd_sc_hs__or3b_2_1/B
+ rst sky130_fd_sc_hs__nor3_1_7/A sky130_fd_sc_hs__nor3_1_7/a_198_368# sky130_fd_sc_hs__nor3_1_7/a_114_368#
+ sky130_fd_sc_hs__nor3_1
Xsky130_fd_sc_hs__xnor2_1_14 DVSS DVDD DVDD DVSS div_ratio_half[5] sky130_fd_sc_hs__xnor2_1_15/Y
+ sky130_fd_sc_hs__xnor2_1_7/A sky130_fd_sc_hs__xnor2_1_15/a_376_368# sky130_fd_sc_hs__xnor2_1_15/a_112_119#
+ sky130_fd_sc_hs__xnor2_1_15/a_138_385# sky130_fd_sc_hs__xnor2_1_15/a_293_74# sky130_fd_sc_hs__xnor2_1
Xsky130_fd_sc_hs__a22oi_1_6 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nor2_1_33/Y sky130_fd_sc_hs__nand2_2_1/B
+ sky130_fd_sc_hs__o21a_1_5/A1 sky130_fd_sc_hs__and2_2_1/X sky130_fd_sc_hs__o21a_1_9/A1
+ sky130_fd_sc_hs__a22oi_1_7/a_71_368# sky130_fd_sc_hs__a22oi_1_7/a_159_74# sky130_fd_sc_hs__a22oi_1_7/a_339_74#
+ sky130_fd_sc_hs__a22oi_1
Xsky130_fd_sc_hs__a21oi_1_91 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__o22ai_1_9/B1 sky130_fd_sc_hs__a21oi_1_91/Y
+ sky130_fd_sc_hs__maj3_1_1/C sky130_fd_sc_hs__maj3_1_1/A sky130_fd_sc_hs__a21oi_1_91/a_117_74#
+ sky130_fd_sc_hs__a21oi_1_91/a_29_368# sky130_fd_sc_hs__a21oi_1
Xsky130_fd_sc_hs__a21oi_1_80 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nor4_1_3/B sky130_fd_sc_hs__a21oi_1_82/Y
+ sky130_fd_sc_hs__inv_4_63/Y sky130_fd_sc_hs__inv_4_67/A sky130_fd_sc_hs__a21oi_1_82/a_117_74#
+ sky130_fd_sc_hs__a21oi_1_82/a_29_368# sky130_fd_sc_hs__a21oi_1
Xsky130_fd_sc_hs__dfrbp_1_36 DVSS DVDD sky130_fd_sc_hs__clkbuf_8_1/X DVDD DVSS sky130_fd_sc_hs__nor3_1_15/A
+ ref_clk sky130_fd_sc_hs__dfrbp_1_37/D sky130_fd_sc_hs__dfrbp_1_37/Q_N sky130_fd_sc_hs__dfrbp_1_37/a_498_360#
+ sky130_fd_sc_hs__dfrbp_1_37/a_1224_74# sky130_fd_sc_hs__dfrbp_1_37/a_2026_424# sky130_fd_sc_hs__dfrbp_1_37/a_1482_48#
+ sky130_fd_sc_hs__dfrbp_1_37/a_125_78# sky130_fd_sc_hs__dfrbp_1_37/a_796_463# sky130_fd_sc_hs__dfrbp_1_37/a_910_118#
+ sky130_fd_sc_hs__dfrbp_1_37/a_1465_471# sky130_fd_sc_hs__dfrbp_1_37/a_832_118# sky130_fd_sc_hs__dfrbp_1_37/a_841_401#
+ sky130_fd_sc_hs__dfrbp_1_37/a_38_78# sky130_fd_sc_hs__dfrbp_1_37/a_1434_74# sky130_fd_sc_hs__dfrbp_1_37/a_706_463#
+ sky130_fd_sc_hs__dfrbp_1_37/a_319_360# sky130_fd_sc_hs__dfrbp_1_37/a_1624_74# sky130_fd_sc_hs__dfrbp_1
Xsky130_fd_sc_hs__dfrbp_1_25 DVSS DVDD sky130_fd_sc_hs__clkbuf_8_1/X DVDD DVSS sky130_fd_sc_hs__o22ai_1_7/A1
+ sky130_fd_sc_hs__clkbuf_2_1/X sky130_fd_sc_hs__o21a_1_53/X sky130_fd_sc_hs__dfrbp_1_25/Q_N
+ sky130_fd_sc_hs__dfrbp_1_25/a_498_360# sky130_fd_sc_hs__dfrbp_1_25/a_1224_74# sky130_fd_sc_hs__dfrbp_1_25/a_2026_424#
+ sky130_fd_sc_hs__dfrbp_1_25/a_1482_48# sky130_fd_sc_hs__dfrbp_1_25/a_125_78# sky130_fd_sc_hs__dfrbp_1_25/a_796_463#
+ sky130_fd_sc_hs__dfrbp_1_25/a_910_118# sky130_fd_sc_hs__dfrbp_1_25/a_1465_471# sky130_fd_sc_hs__dfrbp_1_25/a_832_118#
+ sky130_fd_sc_hs__dfrbp_1_25/a_841_401# sky130_fd_sc_hs__dfrbp_1_25/a_38_78# sky130_fd_sc_hs__dfrbp_1_25/a_1434_74#
+ sky130_fd_sc_hs__dfrbp_1_25/a_706_463# sky130_fd_sc_hs__dfrbp_1_25/a_319_360# sky130_fd_sc_hs__dfrbp_1_25/a_1624_74#
+ sky130_fd_sc_hs__dfrbp_1
Xsky130_fd_sc_hs__dfrbp_1_14 DVSS DVDD sky130_fd_sc_hs__clkbuf_8_1/X DVDD DVSS sky130_fd_sc_hs__inv_4_67/A
+ sky130_fd_sc_hs__clkbuf_2_1/X sky130_fd_sc_hs__dfrbp_1_15/D sky130_fd_sc_hs__dfrbp_1_15/Q_N
+ sky130_fd_sc_hs__dfrbp_1_15/a_498_360# sky130_fd_sc_hs__dfrbp_1_15/a_1224_74# sky130_fd_sc_hs__dfrbp_1_15/a_2026_424#
+ sky130_fd_sc_hs__dfrbp_1_15/a_1482_48# sky130_fd_sc_hs__dfrbp_1_15/a_125_78# sky130_fd_sc_hs__dfrbp_1_15/a_796_463#
+ sky130_fd_sc_hs__dfrbp_1_15/a_910_118# sky130_fd_sc_hs__dfrbp_1_15/a_1465_471# sky130_fd_sc_hs__dfrbp_1_15/a_832_118#
+ sky130_fd_sc_hs__dfrbp_1_15/a_841_401# sky130_fd_sc_hs__dfrbp_1_15/a_38_78# sky130_fd_sc_hs__dfrbp_1_15/a_1434_74#
+ sky130_fd_sc_hs__dfrbp_1_15/a_706_463# sky130_fd_sc_hs__dfrbp_1_15/a_319_360# sky130_fd_sc_hs__dfrbp_1_15/a_1624_74#
+ sky130_fd_sc_hs__dfrbp_1
Xsky130_fd_sc_hs__a222oi_1_0 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nor2_1_33/Y sky130_fd_sc_hs__o21a_1_27/A1
+ sky130_fd_sc_hs__o21a_1_25/A1 sky130_fd_sc_hs__nor2b_1_23/Y sky130_fd_sc_hs__o21ai_1_3/B1
+ sky130_fd_sc_hs__a222oi_1_1/Y sky130_fd_sc_hs__nor2b_1_25/Y sky130_fd_sc_hs__a222oi_1_1/a_461_74#
+ sky130_fd_sc_hs__a222oi_1_1/a_697_74# sky130_fd_sc_hs__a222oi_1_1/a_119_74# sky130_fd_sc_hs__a222oi_1_1/a_116_392#
+ sky130_fd_sc_hs__a222oi_1_1/a_369_392# sky130_fd_sc_hs__a222oi_1
Xsky130_fd_sc_hs__dfrbp_1_47 DVSS DVDD sky130_fd_sc_hs__clkbuf_8_1/X DVDD DVSS sky130_fd_sc_hs__or2_1_3/A
+ ref_clk sky130_fd_sc_hs__o21a_1_73/X sky130_fd_sc_hs__dfrbp_1_47/Q_N sky130_fd_sc_hs__dfrbp_1_47/a_498_360#
+ sky130_fd_sc_hs__dfrbp_1_47/a_1224_74# sky130_fd_sc_hs__dfrbp_1_47/a_2026_424# sky130_fd_sc_hs__dfrbp_1_47/a_1482_48#
+ sky130_fd_sc_hs__dfrbp_1_47/a_125_78# sky130_fd_sc_hs__dfrbp_1_47/a_796_463# sky130_fd_sc_hs__dfrbp_1_47/a_910_118#
+ sky130_fd_sc_hs__dfrbp_1_47/a_1465_471# sky130_fd_sc_hs__dfrbp_1_47/a_832_118# sky130_fd_sc_hs__dfrbp_1_47/a_841_401#
+ sky130_fd_sc_hs__dfrbp_1_47/a_38_78# sky130_fd_sc_hs__dfrbp_1_47/a_1434_74# sky130_fd_sc_hs__dfrbp_1_47/a_706_463#
+ sky130_fd_sc_hs__dfrbp_1_47/a_319_360# sky130_fd_sc_hs__dfrbp_1_47/a_1624_74# sky130_fd_sc_hs__dfrbp_1
Xsky130_fd_sc_hs__nand2_2_15 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand3_1_1/C div_ratio_half[3]
+ sky130_fd_sc_hs__xnor2_1_3/A sky130_fd_sc_hs__nand2_2_15/a_27_74# sky130_fd_sc_hs__nand2_2
Xsky130_fd_sc_hs__xor2_1_3 DVSS DVDD DVDD DVSS fine_con_step_size[1] sky130_fd_sc_hs__fa_2_9/B
+ sky130_fd_sc_hs__fa_2_5/A sky130_fd_sc_hs__xor2_1_3/a_194_125# sky130_fd_sc_hs__xor2_1_3/a_355_368#
+ sky130_fd_sc_hs__xor2_1_3/a_455_87# sky130_fd_sc_hs__xor2_1_3/a_158_392# sky130_fd_sc_hs__xor2_1
Xsky130_fd_sc_hs__a21oi_1_5 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nor2_1_5/Y sky130_fd_sc_hs__dfrtp_4_5/D
+ sky130_fd_sc_hs__nor2_1_5/B sky130_fd_sc_hs__inv_4_7/Y sky130_fd_sc_hs__a21oi_1_5/a_117_74#
+ sky130_fd_sc_hs__a21oi_1_5/a_29_368# sky130_fd_sc_hs__a21oi_1
Xsky130_fd_sc_hs__dfrtn_1_26 DVSS DVDD sky130_fd_sc_hs__clkbuf_8_1/X DVDD DVSS ref_clk
+ sky130_fd_sc_hs__inv_4_93/A sky130_fd_sc_hs__o21a_1_57/X sky130_fd_sc_hs__dfrtn_1_27/a_1266_119#
+ sky130_fd_sc_hs__dfrtn_1_27/a_1736_119# sky130_fd_sc_hs__dfrtn_1_27/a_817_508# sky130_fd_sc_hs__dfrtn_1_27/a_120_74#
+ sky130_fd_sc_hs__dfrtn_1_27/a_1547_508# sky130_fd_sc_hs__dfrtn_1_27/a_922_127# sky130_fd_sc_hs__dfrtn_1_27/a_33_74#
+ sky130_fd_sc_hs__dfrtn_1_27/a_714_127# sky130_fd_sc_hs__dfrtn_1_27/a_1934_94# sky130_fd_sc_hs__dfrtn_1_27/a_1550_119#
+ sky130_fd_sc_hs__dfrtn_1_27/a_1598_93# sky130_fd_sc_hs__dfrtn_1_27/a_300_74# sky130_fd_sc_hs__dfrtn_1_27/a_507_368#
+ sky130_fd_sc_hs__dfrtn_1_27/a_856_304# sky130_fd_sc_hs__dfrtn_1_27/a_850_127# sky130_fd_sc_hs__dfrtn_1
Xsky130_fd_sc_hs__dfrtn_1_15 DVSS DVDD sky130_fd_sc_hs__clkbuf_8_1/X DVDD DVSS sky130_fd_sc_hs__clkbuf_2_1/X
+ sky130_fd_sc_hs__inv_4_65/A sky130_fd_sc_hs__dfrtn_1_15/D sky130_fd_sc_hs__dfrtn_1_15/a_1266_119#
+ sky130_fd_sc_hs__dfrtn_1_15/a_1736_119# sky130_fd_sc_hs__dfrtn_1_15/a_817_508# sky130_fd_sc_hs__dfrtn_1_15/a_120_74#
+ sky130_fd_sc_hs__dfrtn_1_15/a_1547_508# sky130_fd_sc_hs__dfrtn_1_15/a_922_127# sky130_fd_sc_hs__dfrtn_1_15/a_33_74#
+ sky130_fd_sc_hs__dfrtn_1_15/a_714_127# sky130_fd_sc_hs__dfrtn_1_15/a_1934_94# sky130_fd_sc_hs__dfrtn_1_15/a_1550_119#
+ sky130_fd_sc_hs__dfrtn_1_15/a_1598_93# sky130_fd_sc_hs__dfrtn_1_15/a_300_74# sky130_fd_sc_hs__dfrtn_1_15/a_507_368#
+ sky130_fd_sc_hs__dfrtn_1_15/a_856_304# sky130_fd_sc_hs__dfrtn_1_15/a_850_127# sky130_fd_sc_hs__dfrtn_1
Xsky130_fd_sc_hs__dfrtn_1_37 DVSS DVDD sky130_fd_sc_hs__clkbuf_8_1/X DVDD DVSS ref_clk
+ sky130_fd_sc_hs__inv_4_111/A sky130_fd_sc_hs__dfrtn_1_37/D sky130_fd_sc_hs__dfrtn_1_37/a_1266_119#
+ sky130_fd_sc_hs__dfrtn_1_37/a_1736_119# sky130_fd_sc_hs__dfrtn_1_37/a_817_508# sky130_fd_sc_hs__dfrtn_1_37/a_120_74#
+ sky130_fd_sc_hs__dfrtn_1_37/a_1547_508# sky130_fd_sc_hs__dfrtn_1_37/a_922_127# sky130_fd_sc_hs__dfrtn_1_37/a_33_74#
+ sky130_fd_sc_hs__dfrtn_1_37/a_714_127# sky130_fd_sc_hs__dfrtn_1_37/a_1934_94# sky130_fd_sc_hs__dfrtn_1_37/a_1550_119#
+ sky130_fd_sc_hs__dfrtn_1_37/a_1598_93# sky130_fd_sc_hs__dfrtn_1_37/a_300_74# sky130_fd_sc_hs__dfrtn_1_37/a_507_368#
+ sky130_fd_sc_hs__dfrtn_1_37/a_856_304# sky130_fd_sc_hs__dfrtn_1_37/a_850_127# sky130_fd_sc_hs__dfrtn_1
Xsky130_fd_sc_hs__dfrtn_1_48 DVSS DVDD sky130_fd_sc_hs__clkbuf_8_1/X DVDD DVSS ref_clk
+ sky130_fd_sc_hs__o21a_1_71/A1 sky130_fd_sc_hs__o21a_1_71/X sky130_fd_sc_hs__dfrtn_1_49/a_1266_119#
+ sky130_fd_sc_hs__dfrtn_1_49/a_1736_119# sky130_fd_sc_hs__dfrtn_1_49/a_817_508# sky130_fd_sc_hs__dfrtn_1_49/a_120_74#
+ sky130_fd_sc_hs__dfrtn_1_49/a_1547_508# sky130_fd_sc_hs__dfrtn_1_49/a_922_127# sky130_fd_sc_hs__dfrtn_1_49/a_33_74#
+ sky130_fd_sc_hs__dfrtn_1_49/a_714_127# sky130_fd_sc_hs__dfrtn_1_49/a_1934_94# sky130_fd_sc_hs__dfrtn_1_49/a_1550_119#
+ sky130_fd_sc_hs__dfrtn_1_49/a_1598_93# sky130_fd_sc_hs__dfrtn_1_49/a_300_74# sky130_fd_sc_hs__dfrtn_1_49/a_507_368#
+ sky130_fd_sc_hs__dfrtn_1_49/a_856_304# sky130_fd_sc_hs__dfrtn_1_49/a_850_127# sky130_fd_sc_hs__dfrtn_1
Xsky130_fd_sc_hs__nand2b_1_1 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_1_47/B sky130_fd_sc_hs__nor2b_1_33/Y
+ sky130_fd_sc_hs__nor2_1_73/B sky130_fd_sc_hs__nand2b_1_1/a_269_74# sky130_fd_sc_hs__nand2b_1_1/a_27_112#
+ sky130_fd_sc_hs__nand2b_1
Xsky130_fd_sc_hs__dfrbp_1_3 DVSS DVDD sky130_fd_sc_hs__clkbuf_8_1/X DVDD DVSS sky130_fd_sc_hs__inv_4_61/A
+ sky130_fd_sc_hs__clkbuf_2_1/X sky130_fd_sc_hs__dfrbp_1_3/D sky130_fd_sc_hs__dfrbp_1_3/Q_N
+ sky130_fd_sc_hs__dfrbp_1_3/a_498_360# sky130_fd_sc_hs__dfrbp_1_3/a_1224_74# sky130_fd_sc_hs__dfrbp_1_3/a_2026_424#
+ sky130_fd_sc_hs__dfrbp_1_3/a_1482_48# sky130_fd_sc_hs__dfrbp_1_3/a_125_78# sky130_fd_sc_hs__dfrbp_1_3/a_796_463#
+ sky130_fd_sc_hs__dfrbp_1_3/a_910_118# sky130_fd_sc_hs__dfrbp_1_3/a_1465_471# sky130_fd_sc_hs__dfrbp_1_3/a_832_118#
+ sky130_fd_sc_hs__dfrbp_1_3/a_841_401# sky130_fd_sc_hs__dfrbp_1_3/a_38_78# sky130_fd_sc_hs__dfrbp_1_3/a_1434_74#
+ sky130_fd_sc_hs__dfrbp_1_3/a_706_463# sky130_fd_sc_hs__dfrbp_1_3/a_319_360# sky130_fd_sc_hs__dfrbp_1_3/a_1624_74#
+ sky130_fd_sc_hs__dfrbp_1
Xsky130_fd_sc_hs__a32oi_1_0 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_2_1/Y fine_control_avg_window_select[1]
+ sky130_fd_sc_hs__a32oi_1_3/B1 sky130_fd_sc_hs__inv_4_21/Y sky130_fd_sc_hs__a32oi_1_1/Y
+ fine_control_avg_window_select[2] sky130_fd_sc_hs__a32oi_1_1/a_391_74# sky130_fd_sc_hs__a32oi_1_1/a_27_368#
+ sky130_fd_sc_hs__a32oi_1_1/a_119_74# sky130_fd_sc_hs__a32oi_1_1/a_469_74# sky130_fd_sc_hs__a32oi_1
Xsky130_fd_sc_hs__dfrtn_1_1 DVSS DVDD sky130_fd_sc_hs__clkbuf_8_1/X DVDD DVSS sky130_fd_sc_hs__clkbuf_2_1/X
+ sky130_fd_sc_hs__inv_4_39/A sky130_fd_sc_hs__o21a_1_29/X sky130_fd_sc_hs__dfrtn_1_1/a_1266_119#
+ sky130_fd_sc_hs__dfrtn_1_1/a_1736_119# sky130_fd_sc_hs__dfrtn_1_1/a_817_508# sky130_fd_sc_hs__dfrtn_1_1/a_120_74#
+ sky130_fd_sc_hs__dfrtn_1_1/a_1547_508# sky130_fd_sc_hs__dfrtn_1_1/a_922_127# sky130_fd_sc_hs__dfrtn_1_1/a_33_74#
+ sky130_fd_sc_hs__dfrtn_1_1/a_714_127# sky130_fd_sc_hs__dfrtn_1_1/a_1934_94# sky130_fd_sc_hs__dfrtn_1_1/a_1550_119#
+ sky130_fd_sc_hs__dfrtn_1_1/a_1598_93# sky130_fd_sc_hs__dfrtn_1_1/a_300_74# sky130_fd_sc_hs__dfrtn_1_1/a_507_368#
+ sky130_fd_sc_hs__dfrtn_1_1/a_856_304# sky130_fd_sc_hs__dfrtn_1_1/a_850_127# sky130_fd_sc_hs__dfrtn_1
Xsky130_fd_sc_hs__o211ai_1_1 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__a21oi_1_91/Y sky130_fd_sc_hs__nor2_1_61/B
+ sky130_fd_sc_hs__nand2_1_67/Y sky130_fd_sc_hs__inv_4_79/Y sky130_fd_sc_hs__inv_4_59/A
+ sky130_fd_sc_hs__o211ai_1_1/a_31_74# sky130_fd_sc_hs__o211ai_1_1/a_311_74# sky130_fd_sc_hs__o211ai_1_1/a_116_368#
+ sky130_fd_sc_hs__o211ai_1
Xsky130_fd_sc_hs__inv_4_26 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_27/Y fine_control_avg_window_select[2]
+ sky130_fd_sc_hs__inv_4
Xsky130_fd_sc_hs__inv_4_15 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_15/Y sky130_fd_sc_hs__inv_4_15/A
+ sky130_fd_sc_hs__inv_4
Xsky130_fd_sc_hs__inv_4_59 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_59/Y sky130_fd_sc_hs__inv_4_59/A
+ sky130_fd_sc_hs__inv_4
Xsky130_fd_sc_hs__inv_4_48 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_49/Y rst sky130_fd_sc_hs__inv_4
Xsky130_fd_sc_hs__inv_4_37 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_37/Y sky130_fd_sc_hs__inv_4_37/A
+ sky130_fd_sc_hs__inv_4
Xsky130_fd_sc_hs__a22o_1_0 DVSS DVDD DVDD DVSS osc_fine_con_final[3] manual_control_osc[3]
+ sky130_fd_sc_hs__inv_4_43/Y sky130_fd_sc_hs__fa_2_1/B fftl_en sky130_fd_sc_hs__a22o_1_1/a_222_392#
+ sky130_fd_sc_hs__a22o_1_1/a_230_79# sky130_fd_sc_hs__a22o_1_1/a_52_123# sky130_fd_sc_hs__a22o_1_1/a_132_392#
+ sky130_fd_sc_hs__a22o_1
Xsky130_fd_sc_hs__fa_2_3 DVSS DVDD sky130_fd_sc_hs__fa_2_3/A DVDD DVSS sky130_fd_sc_hs__fa_2_3/CIN
+ sky130_fd_sc_hs__fa_2_3/B sky130_fd_sc_hs__fa_2_1/CIN sky130_fd_sc_hs__fa_2_3/SUM
+ sky130_fd_sc_hs__fa_2_3/a_27_378# sky130_fd_sc_hs__fa_2_3/a_701_79# sky130_fd_sc_hs__fa_2_3/a_484_347#
+ sky130_fd_sc_hs__fa_2_3/a_1094_347# sky130_fd_sc_hs__fa_2_3/a_1205_79# sky130_fd_sc_hs__fa_2_3/a_27_79#
+ sky130_fd_sc_hs__fa_2_3/a_1202_368# sky130_fd_sc_hs__fa_2_3/a_336_347# sky130_fd_sc_hs__fa_2_3/a_992_347#
+ sky130_fd_sc_hs__fa_2_3/a_1119_79# sky130_fd_sc_hs__fa_2_3/a_487_79# sky130_fd_sc_hs__fa_2_3/a_683_347#
+ sky130_fd_sc_hs__fa_2
Xsky130_fd_sc_hs__nor3_1_7 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nor3_1_7/Y sky130_fd_sc_hs__or3b_2_1/B
+ rst sky130_fd_sc_hs__nor3_1_7/A sky130_fd_sc_hs__nor3_1_7/a_198_368# sky130_fd_sc_hs__nor3_1_7/a_114_368#
+ sky130_fd_sc_hs__nor3_1
Xsky130_fd_sc_hs__xnor2_1_15 DVSS DVDD DVDD DVSS div_ratio_half[5] sky130_fd_sc_hs__xnor2_1_15/Y
+ sky130_fd_sc_hs__xnor2_1_7/A sky130_fd_sc_hs__xnor2_1_15/a_376_368# sky130_fd_sc_hs__xnor2_1_15/a_112_119#
+ sky130_fd_sc_hs__xnor2_1_15/a_138_385# sky130_fd_sc_hs__xnor2_1_15/a_293_74# sky130_fd_sc_hs__xnor2_1
Xsky130_fd_sc_hs__nand2_1_0 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nor2_1_1/Y sky130_fd_sc_hs__nor2_1_3/B
+ sky130_fd_sc_hs__o21a_1_3/A1 sky130_fd_sc_hs__nand2_1_1/a_117_74# sky130_fd_sc_hs__nand2_1
Xsky130_fd_sc_hs__a22oi_1_7 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nor2_1_33/Y sky130_fd_sc_hs__nand2_2_1/B
+ sky130_fd_sc_hs__o21a_1_5/A1 sky130_fd_sc_hs__and2_2_1/X sky130_fd_sc_hs__o21a_1_9/A1
+ sky130_fd_sc_hs__a22oi_1_7/a_71_368# sky130_fd_sc_hs__a22oi_1_7/a_159_74# sky130_fd_sc_hs__a22oi_1_7/a_339_74#
+ sky130_fd_sc_hs__a22oi_1
Xsky130_fd_sc_hs__a21oi_1_92 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nor3_1_13/C sky130_fd_sc_hs__a21oi_1_93/Y
+ sky130_fd_sc_hs__nand4_1_1/C sky130_fd_sc_hs__o31ai_1_7/Y sky130_fd_sc_hs__a21oi_1_93/a_117_74#
+ sky130_fd_sc_hs__a21oi_1_93/a_29_368# sky130_fd_sc_hs__a21oi_1
Xsky130_fd_sc_hs__a21oi_1_81 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nor3_1_5/B sky130_fd_sc_hs__o31ai_1_3/B1
+ sky130_fd_sc_hs__nor4_1_3/A sky130_fd_sc_hs__a21oi_1_82/Y sky130_fd_sc_hs__a21oi_1_83/a_117_74#
+ sky130_fd_sc_hs__a21oi_1_83/a_29_368# sky130_fd_sc_hs__a21oi_1
Xsky130_fd_sc_hs__a21oi_1_70 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nor2_1_73/Y sky130_fd_sc_hs__dfrbp_1_21/D
+ sky130_fd_sc_hs__nor2_1_73/B sky130_fd_sc_hs__inv_4_85/Y sky130_fd_sc_hs__a21oi_1_71/a_117_74#
+ sky130_fd_sc_hs__a21oi_1_71/a_29_368# sky130_fd_sc_hs__a21oi_1
Xsky130_fd_sc_hs__dfrbp_1_26 DVSS DVDD sky130_fd_sc_hs__clkbuf_8_1/X DVDD DVSS sky130_fd_sc_hs__inv_4_95/A
+ ref_clk sky130_fd_sc_hs__xnor2_1_5/Y sky130_fd_sc_hs__dfrbp_1_27/Q_N sky130_fd_sc_hs__dfrbp_1_27/a_498_360#
+ sky130_fd_sc_hs__dfrbp_1_27/a_1224_74# sky130_fd_sc_hs__dfrbp_1_27/a_2026_424# sky130_fd_sc_hs__dfrbp_1_27/a_1482_48#
+ sky130_fd_sc_hs__dfrbp_1_27/a_125_78# sky130_fd_sc_hs__dfrbp_1_27/a_796_463# sky130_fd_sc_hs__dfrbp_1_27/a_910_118#
+ sky130_fd_sc_hs__dfrbp_1_27/a_1465_471# sky130_fd_sc_hs__dfrbp_1_27/a_832_118# sky130_fd_sc_hs__dfrbp_1_27/a_841_401#
+ sky130_fd_sc_hs__dfrbp_1_27/a_38_78# sky130_fd_sc_hs__dfrbp_1_27/a_1434_74# sky130_fd_sc_hs__dfrbp_1_27/a_706_463#
+ sky130_fd_sc_hs__dfrbp_1_27/a_319_360# sky130_fd_sc_hs__dfrbp_1_27/a_1624_74# sky130_fd_sc_hs__dfrbp_1
Xsky130_fd_sc_hs__dfrbp_1_37 DVSS DVDD sky130_fd_sc_hs__clkbuf_8_1/X DVDD DVSS sky130_fd_sc_hs__nor3_1_15/A
+ ref_clk sky130_fd_sc_hs__dfrbp_1_37/D sky130_fd_sc_hs__dfrbp_1_37/Q_N sky130_fd_sc_hs__dfrbp_1_37/a_498_360#
+ sky130_fd_sc_hs__dfrbp_1_37/a_1224_74# sky130_fd_sc_hs__dfrbp_1_37/a_2026_424# sky130_fd_sc_hs__dfrbp_1_37/a_1482_48#
+ sky130_fd_sc_hs__dfrbp_1_37/a_125_78# sky130_fd_sc_hs__dfrbp_1_37/a_796_463# sky130_fd_sc_hs__dfrbp_1_37/a_910_118#
+ sky130_fd_sc_hs__dfrbp_1_37/a_1465_471# sky130_fd_sc_hs__dfrbp_1_37/a_832_118# sky130_fd_sc_hs__dfrbp_1_37/a_841_401#
+ sky130_fd_sc_hs__dfrbp_1_37/a_38_78# sky130_fd_sc_hs__dfrbp_1_37/a_1434_74# sky130_fd_sc_hs__dfrbp_1_37/a_706_463#
+ sky130_fd_sc_hs__dfrbp_1_37/a_319_360# sky130_fd_sc_hs__dfrbp_1_37/a_1624_74# sky130_fd_sc_hs__dfrbp_1
Xsky130_fd_sc_hs__dfrbp_1_15 DVSS DVDD sky130_fd_sc_hs__clkbuf_8_1/X DVDD DVSS sky130_fd_sc_hs__inv_4_67/A
+ sky130_fd_sc_hs__clkbuf_2_1/X sky130_fd_sc_hs__dfrbp_1_15/D sky130_fd_sc_hs__dfrbp_1_15/Q_N
+ sky130_fd_sc_hs__dfrbp_1_15/a_498_360# sky130_fd_sc_hs__dfrbp_1_15/a_1224_74# sky130_fd_sc_hs__dfrbp_1_15/a_2026_424#
+ sky130_fd_sc_hs__dfrbp_1_15/a_1482_48# sky130_fd_sc_hs__dfrbp_1_15/a_125_78# sky130_fd_sc_hs__dfrbp_1_15/a_796_463#
+ sky130_fd_sc_hs__dfrbp_1_15/a_910_118# sky130_fd_sc_hs__dfrbp_1_15/a_1465_471# sky130_fd_sc_hs__dfrbp_1_15/a_832_118#
+ sky130_fd_sc_hs__dfrbp_1_15/a_841_401# sky130_fd_sc_hs__dfrbp_1_15/a_38_78# sky130_fd_sc_hs__dfrbp_1_15/a_1434_74#
+ sky130_fd_sc_hs__dfrbp_1_15/a_706_463# sky130_fd_sc_hs__dfrbp_1_15/a_319_360# sky130_fd_sc_hs__dfrbp_1_15/a_1624_74#
+ sky130_fd_sc_hs__dfrbp_1
Xsky130_fd_sc_hs__a222oi_1_1 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nor2_1_33/Y sky130_fd_sc_hs__o21a_1_27/A1
+ sky130_fd_sc_hs__o21a_1_25/A1 sky130_fd_sc_hs__nor2b_1_23/Y sky130_fd_sc_hs__o21ai_1_3/B1
+ sky130_fd_sc_hs__a222oi_1_1/Y sky130_fd_sc_hs__nor2b_1_25/Y sky130_fd_sc_hs__a222oi_1_1/a_461_74#
+ sky130_fd_sc_hs__a222oi_1_1/a_697_74# sky130_fd_sc_hs__a222oi_1_1/a_119_74# sky130_fd_sc_hs__a222oi_1_1/a_116_392#
+ sky130_fd_sc_hs__a222oi_1_1/a_369_392# sky130_fd_sc_hs__a222oi_1
Xsky130_fd_sc_hs__xor2_1_4 DVSS DVDD DVDD DVSS fine_con_step_size[2] sky130_fd_sc_hs__fa_2_9/B
+ sky130_fd_sc_hs__fa_2_3/A sky130_fd_sc_hs__xor2_1_5/a_194_125# sky130_fd_sc_hs__xor2_1_5/a_355_368#
+ sky130_fd_sc_hs__xor2_1_5/a_455_87# sky130_fd_sc_hs__xor2_1_5/a_158_392# sky130_fd_sc_hs__xor2_1
Xsky130_fd_sc_hs__a21oi_1_6 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nor2_1_9/Y sky130_fd_sc_hs__dfrtp_4_7/D
+ sky130_fd_sc_hs__nor2_1_9/B sky130_fd_sc_hs__inv_4_9/Y sky130_fd_sc_hs__a21oi_1_7/a_117_74#
+ sky130_fd_sc_hs__a21oi_1_7/a_29_368# sky130_fd_sc_hs__a21oi_1
Xsky130_fd_sc_hs__dfrtn_1_27 DVSS DVDD sky130_fd_sc_hs__clkbuf_8_1/X DVDD DVSS ref_clk
+ sky130_fd_sc_hs__inv_4_93/A sky130_fd_sc_hs__o21a_1_57/X sky130_fd_sc_hs__dfrtn_1_27/a_1266_119#
+ sky130_fd_sc_hs__dfrtn_1_27/a_1736_119# sky130_fd_sc_hs__dfrtn_1_27/a_817_508# sky130_fd_sc_hs__dfrtn_1_27/a_120_74#
+ sky130_fd_sc_hs__dfrtn_1_27/a_1547_508# sky130_fd_sc_hs__dfrtn_1_27/a_922_127# sky130_fd_sc_hs__dfrtn_1_27/a_33_74#
+ sky130_fd_sc_hs__dfrtn_1_27/a_714_127# sky130_fd_sc_hs__dfrtn_1_27/a_1934_94# sky130_fd_sc_hs__dfrtn_1_27/a_1550_119#
+ sky130_fd_sc_hs__dfrtn_1_27/a_1598_93# sky130_fd_sc_hs__dfrtn_1_27/a_300_74# sky130_fd_sc_hs__dfrtn_1_27/a_507_368#
+ sky130_fd_sc_hs__dfrtn_1_27/a_856_304# sky130_fd_sc_hs__dfrtn_1_27/a_850_127# sky130_fd_sc_hs__dfrtn_1
Xsky130_fd_sc_hs__dfrtn_1_16 DVSS DVDD sky130_fd_sc_hs__clkbuf_8_1/X DVDD DVSS sky130_fd_sc_hs__clkbuf_2_1/X
+ sky130_fd_sc_hs__inv_4_63/A sky130_fd_sc_hs__dfrtn_1_17/D sky130_fd_sc_hs__dfrtn_1_17/a_1266_119#
+ sky130_fd_sc_hs__dfrtn_1_17/a_1736_119# sky130_fd_sc_hs__dfrtn_1_17/a_817_508# sky130_fd_sc_hs__dfrtn_1_17/a_120_74#
+ sky130_fd_sc_hs__dfrtn_1_17/a_1547_508# sky130_fd_sc_hs__dfrtn_1_17/a_922_127# sky130_fd_sc_hs__dfrtn_1_17/a_33_74#
+ sky130_fd_sc_hs__dfrtn_1_17/a_714_127# sky130_fd_sc_hs__dfrtn_1_17/a_1934_94# sky130_fd_sc_hs__dfrtn_1_17/a_1550_119#
+ sky130_fd_sc_hs__dfrtn_1_17/a_1598_93# sky130_fd_sc_hs__dfrtn_1_17/a_300_74# sky130_fd_sc_hs__dfrtn_1_17/a_507_368#
+ sky130_fd_sc_hs__dfrtn_1_17/a_856_304# sky130_fd_sc_hs__dfrtn_1_17/a_850_127# sky130_fd_sc_hs__dfrtn_1
Xsky130_fd_sc_hs__dfrtn_1_38 DVSS DVDD sky130_fd_sc_hs__clkbuf_8_1/X DVDD DVSS ref_clk
+ sky130_fd_sc_hs__inv_4_125/A sky130_fd_sc_hs__dfrtn_1_39/D sky130_fd_sc_hs__dfrtn_1_39/a_1266_119#
+ sky130_fd_sc_hs__dfrtn_1_39/a_1736_119# sky130_fd_sc_hs__dfrtn_1_39/a_817_508# sky130_fd_sc_hs__dfrtn_1_39/a_120_74#
+ sky130_fd_sc_hs__dfrtn_1_39/a_1547_508# sky130_fd_sc_hs__dfrtn_1_39/a_922_127# sky130_fd_sc_hs__dfrtn_1_39/a_33_74#
+ sky130_fd_sc_hs__dfrtn_1_39/a_714_127# sky130_fd_sc_hs__dfrtn_1_39/a_1934_94# sky130_fd_sc_hs__dfrtn_1_39/a_1550_119#
+ sky130_fd_sc_hs__dfrtn_1_39/a_1598_93# sky130_fd_sc_hs__dfrtn_1_39/a_300_74# sky130_fd_sc_hs__dfrtn_1_39/a_507_368#
+ sky130_fd_sc_hs__dfrtn_1_39/a_856_304# sky130_fd_sc_hs__dfrtn_1_39/a_850_127# sky130_fd_sc_hs__dfrtn_1
Xsky130_fd_sc_hs__dfrtn_1_49 DVSS DVDD sky130_fd_sc_hs__clkbuf_8_1/X DVDD DVSS ref_clk
+ sky130_fd_sc_hs__o21a_1_71/A1 sky130_fd_sc_hs__o21a_1_71/X sky130_fd_sc_hs__dfrtn_1_49/a_1266_119#
+ sky130_fd_sc_hs__dfrtn_1_49/a_1736_119# sky130_fd_sc_hs__dfrtn_1_49/a_817_508# sky130_fd_sc_hs__dfrtn_1_49/a_120_74#
+ sky130_fd_sc_hs__dfrtn_1_49/a_1547_508# sky130_fd_sc_hs__dfrtn_1_49/a_922_127# sky130_fd_sc_hs__dfrtn_1_49/a_33_74#
+ sky130_fd_sc_hs__dfrtn_1_49/a_714_127# sky130_fd_sc_hs__dfrtn_1_49/a_1934_94# sky130_fd_sc_hs__dfrtn_1_49/a_1550_119#
+ sky130_fd_sc_hs__dfrtn_1_49/a_1598_93# sky130_fd_sc_hs__dfrtn_1_49/a_300_74# sky130_fd_sc_hs__dfrtn_1_49/a_507_368#
+ sky130_fd_sc_hs__dfrtn_1_49/a_856_304# sky130_fd_sc_hs__dfrtn_1_49/a_850_127# sky130_fd_sc_hs__dfrtn_1
Xsky130_fd_sc_hs__nand2b_1_2 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_87/A sky130_fd_sc_hs__nor2_1_53/Y
+ sky130_fd_sc_hs__nand2b_1_3/Y sky130_fd_sc_hs__nand2b_1_3/a_269_74# sky130_fd_sc_hs__nand2b_1_3/a_27_112#
+ sky130_fd_sc_hs__nand2b_1
Xsky130_fd_sc_hs__dfrbp_1_4 DVSS DVDD sky130_fd_sc_hs__clkbuf_8_1/X DVDD DVSS sky130_fd_sc_hs__inv_4_51/A
+ sky130_fd_sc_hs__clkbuf_2_1/X sky130_fd_sc_hs__dfrbp_1_5/D sky130_fd_sc_hs__dfrbp_1_5/Q_N
+ sky130_fd_sc_hs__dfrbp_1_5/a_498_360# sky130_fd_sc_hs__dfrbp_1_5/a_1224_74# sky130_fd_sc_hs__dfrbp_1_5/a_2026_424#
+ sky130_fd_sc_hs__dfrbp_1_5/a_1482_48# sky130_fd_sc_hs__dfrbp_1_5/a_125_78# sky130_fd_sc_hs__dfrbp_1_5/a_796_463#
+ sky130_fd_sc_hs__dfrbp_1_5/a_910_118# sky130_fd_sc_hs__dfrbp_1_5/a_1465_471# sky130_fd_sc_hs__dfrbp_1_5/a_832_118#
+ sky130_fd_sc_hs__dfrbp_1_5/a_841_401# sky130_fd_sc_hs__dfrbp_1_5/a_38_78# sky130_fd_sc_hs__dfrbp_1_5/a_1434_74#
+ sky130_fd_sc_hs__dfrbp_1_5/a_706_463# sky130_fd_sc_hs__dfrbp_1_5/a_319_360# sky130_fd_sc_hs__dfrbp_1_5/a_1624_74#
+ sky130_fd_sc_hs__dfrbp_1
Xsky130_fd_sc_hs__a32oi_1_1 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_2_1/Y fine_control_avg_window_select[1]
+ sky130_fd_sc_hs__a32oi_1_3/B1 sky130_fd_sc_hs__inv_4_21/Y sky130_fd_sc_hs__a32oi_1_1/Y
+ fine_control_avg_window_select[2] sky130_fd_sc_hs__a32oi_1_1/a_391_74# sky130_fd_sc_hs__a32oi_1_1/a_27_368#
+ sky130_fd_sc_hs__a32oi_1_1/a_119_74# sky130_fd_sc_hs__a32oi_1_1/a_469_74# sky130_fd_sc_hs__a32oi_1
Xsky130_fd_sc_hs__dfrtn_1_2 DVSS DVDD sky130_fd_sc_hs__clkbuf_8_1/X DVDD DVSS sky130_fd_sc_hs__clkbuf_2_1/X
+ sky130_fd_sc_hs__inv_4_37/A sky130_fd_sc_hs__dfrtn_1_3/D sky130_fd_sc_hs__dfrtn_1_3/a_1266_119#
+ sky130_fd_sc_hs__dfrtn_1_3/a_1736_119# sky130_fd_sc_hs__dfrtn_1_3/a_817_508# sky130_fd_sc_hs__dfrtn_1_3/a_120_74#
+ sky130_fd_sc_hs__dfrtn_1_3/a_1547_508# sky130_fd_sc_hs__dfrtn_1_3/a_922_127# sky130_fd_sc_hs__dfrtn_1_3/a_33_74#
+ sky130_fd_sc_hs__dfrtn_1_3/a_714_127# sky130_fd_sc_hs__dfrtn_1_3/a_1934_94# sky130_fd_sc_hs__dfrtn_1_3/a_1550_119#
+ sky130_fd_sc_hs__dfrtn_1_3/a_1598_93# sky130_fd_sc_hs__dfrtn_1_3/a_300_74# sky130_fd_sc_hs__dfrtn_1_3/a_507_368#
+ sky130_fd_sc_hs__dfrtn_1_3/a_856_304# sky130_fd_sc_hs__dfrtn_1_3/a_850_127# sky130_fd_sc_hs__dfrtn_1
Xsky130_fd_sc_hs__o211ai_1_2 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__a21oi_1_82/Y sky130_fd_sc_hs__o211ai_1_3/Y
+ sky130_fd_sc_hs__nand4_1_5/A sky130_fd_sc_hs__a21oi_1_93/Y sky130_fd_sc_hs__nor3_1_1/A
+ sky130_fd_sc_hs__o211ai_1_3/a_31_74# sky130_fd_sc_hs__o211ai_1_3/a_311_74# sky130_fd_sc_hs__o211ai_1_3/a_116_368#
+ sky130_fd_sc_hs__o211ai_1
Xsky130_fd_sc_hs__a31oi_1_0 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__dfstp_2_7/D sky130_fd_sc_hs__nand2_1_71/Y
+ sky130_fd_sc_hs__nor4_1_1/A sky130_fd_sc_hs__a31oi_1_1/A2 sky130_fd_sc_hs__maj3_1_3/X
+ sky130_fd_sc_hs__a31oi_1_1/a_136_368# sky130_fd_sc_hs__a31oi_1_1/a_223_74# sky130_fd_sc_hs__a31oi_1_1/a_145_74#
+ sky130_fd_sc_hs__a31oi_1
Xsky130_fd_sc_hs__inv_4_16 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_17/Y sky130_fd_sc_hs__inv_4_17/A
+ sky130_fd_sc_hs__inv_4
Xsky130_fd_sc_hs__inv_4_49 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_49/Y rst sky130_fd_sc_hs__inv_4
Xsky130_fd_sc_hs__inv_4_38 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_39/Y sky130_fd_sc_hs__inv_4_39/A
+ sky130_fd_sc_hs__inv_4
Xsky130_fd_sc_hs__inv_4_27 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_27/Y fine_control_avg_window_select[2]
+ sky130_fd_sc_hs__inv_4
Xsky130_fd_sc_hs__a22o_1_1 DVSS DVDD DVDD DVSS osc_fine_con_final[3] manual_control_osc[3]
+ sky130_fd_sc_hs__inv_4_43/Y sky130_fd_sc_hs__fa_2_1/B fftl_en sky130_fd_sc_hs__a22o_1_1/a_222_392#
+ sky130_fd_sc_hs__a22o_1_1/a_230_79# sky130_fd_sc_hs__a22o_1_1/a_52_123# sky130_fd_sc_hs__a22o_1_1/a_132_392#
+ sky130_fd_sc_hs__a22o_1
Xsky130_fd_sc_hs__dfrtp_4_90 DVSS DVDD sky130_fd_sc_hs__inv_4_49/Y DVDD DVSS sky130_fd_sc_hs__nor2b_1_27/Y
+ sky130_fd_sc_hs__dfstp_2_1/CLK sky130_fd_sc_hs__fa_2_19/B sky130_fd_sc_hs__dfrtp_4_91/a_37_78#
+ sky130_fd_sc_hs__dfrtp_4_91/a_494_366# sky130_fd_sc_hs__dfrtp_4_91/a_699_463# sky130_fd_sc_hs__dfrtp_4_91/a_313_74#
+ sky130_fd_sc_hs__dfrtp_4_91/a_1627_493# sky130_fd_sc_hs__dfrtp_4_91/a_1678_395#
+ sky130_fd_sc_hs__dfrtp_4_91/a_1827_81# sky130_fd_sc_hs__dfrtp_4_91/a_789_463# sky130_fd_sc_hs__dfrtp_4_91/a_1350_392#
+ sky130_fd_sc_hs__dfrtp_4_91/a_834_355# sky130_fd_sc_hs__dfrtp_4_91/a_812_138# sky130_fd_sc_hs__dfrtp_4_91/a_124_78#
+ sky130_fd_sc_hs__dfrtp_4_91/a_1647_81# sky130_fd_sc_hs__dfrtp_4_91/a_2010_409# sky130_fd_sc_hs__dfrtp_4_91/a_890_138#
+ sky130_fd_sc_hs__dfrtp_4
Xsky130_fd_sc_hs__fa_2_4 DVSS DVDD sky130_fd_sc_hs__fa_2_5/A DVDD DVSS sky130_fd_sc_hs__fa_2_5/CIN
+ sky130_fd_sc_hs__fa_2_5/B sky130_fd_sc_hs__fa_2_3/CIN sky130_fd_sc_hs__fa_2_5/SUM
+ sky130_fd_sc_hs__fa_2_5/a_27_378# sky130_fd_sc_hs__fa_2_5/a_701_79# sky130_fd_sc_hs__fa_2_5/a_484_347#
+ sky130_fd_sc_hs__fa_2_5/a_1094_347# sky130_fd_sc_hs__fa_2_5/a_1205_79# sky130_fd_sc_hs__fa_2_5/a_27_79#
+ sky130_fd_sc_hs__fa_2_5/a_1202_368# sky130_fd_sc_hs__fa_2_5/a_336_347# sky130_fd_sc_hs__fa_2_5/a_992_347#
+ sky130_fd_sc_hs__fa_2_5/a_1119_79# sky130_fd_sc_hs__fa_2_5/a_487_79# sky130_fd_sc_hs__fa_2_5/a_683_347#
+ sky130_fd_sc_hs__fa_2
Xsky130_fd_sc_hs__nor3_1_8 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nor3_1_9/Y sky130_fd_sc_hs__nor3_1_9/C
+ sky130_fd_sc_hs__nor3_1_9/B sky130_fd_sc_hs__nor3_1_9/A sky130_fd_sc_hs__nor3_1_9/a_198_368#
+ sky130_fd_sc_hs__nor3_1_9/a_114_368# sky130_fd_sc_hs__nor3_1
Xsky130_fd_sc_hs__nand2_1_1 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nor2_1_1/Y sky130_fd_sc_hs__nor2_1_3/B
+ sky130_fd_sc_hs__o21a_1_3/A1 sky130_fd_sc_hs__nand2_1_1/a_117_74# sky130_fd_sc_hs__nand2_1
Xsky130_fd_sc_hs__a22oi_1_8 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nor2b_1_25/Y sky130_fd_sc_hs__nand2_2_3/A
+ sky130_fd_sc_hs__o21a_1_17/A1 sky130_fd_sc_hs__nor2b_1_23/Y sky130_fd_sc_hs__o21a_1_7/A1
+ sky130_fd_sc_hs__a22oi_1_9/a_71_368# sky130_fd_sc_hs__a22oi_1_9/a_159_74# sky130_fd_sc_hs__a22oi_1_9/a_339_74#
+ sky130_fd_sc_hs__a22oi_1
Xsky130_fd_sc_hs__a21oi_1_82 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nor4_1_3/B sky130_fd_sc_hs__a21oi_1_82/Y
+ sky130_fd_sc_hs__inv_4_63/Y sky130_fd_sc_hs__inv_4_67/A sky130_fd_sc_hs__a21oi_1_82/a_117_74#
+ sky130_fd_sc_hs__a21oi_1_82/a_29_368# sky130_fd_sc_hs__a21oi_1
Xsky130_fd_sc_hs__a21oi_1_71 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nor2_1_73/Y sky130_fd_sc_hs__dfrbp_1_21/D
+ sky130_fd_sc_hs__nor2_1_73/B sky130_fd_sc_hs__inv_4_85/Y sky130_fd_sc_hs__a21oi_1_71/a_117_74#
+ sky130_fd_sc_hs__a21oi_1_71/a_29_368# sky130_fd_sc_hs__a21oi_1
Xsky130_fd_sc_hs__a21oi_1_60 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__a22o_1_27/X sky130_fd_sc_hs__o21ai_1_5/B1
+ sky130_fd_sc_hs__inv_4_55/Y sky130_fd_sc_hs__nor2_1_59/A sky130_fd_sc_hs__a21oi_1_61/a_117_74#
+ sky130_fd_sc_hs__a21oi_1_61/a_29_368# sky130_fd_sc_hs__a21oi_1
Xsky130_fd_sc_hs__a21oi_1_93 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nor3_1_13/C sky130_fd_sc_hs__a21oi_1_93/Y
+ sky130_fd_sc_hs__nand4_1_1/C sky130_fd_sc_hs__o31ai_1_7/Y sky130_fd_sc_hs__a21oi_1_93/a_117_74#
+ sky130_fd_sc_hs__a21oi_1_93/a_29_368# sky130_fd_sc_hs__a21oi_1
Xsky130_fd_sc_hs__dfrbp_1_27 DVSS DVDD sky130_fd_sc_hs__clkbuf_8_1/X DVDD DVSS sky130_fd_sc_hs__inv_4_95/A
+ ref_clk sky130_fd_sc_hs__xnor2_1_5/Y sky130_fd_sc_hs__dfrbp_1_27/Q_N sky130_fd_sc_hs__dfrbp_1_27/a_498_360#
+ sky130_fd_sc_hs__dfrbp_1_27/a_1224_74# sky130_fd_sc_hs__dfrbp_1_27/a_2026_424# sky130_fd_sc_hs__dfrbp_1_27/a_1482_48#
+ sky130_fd_sc_hs__dfrbp_1_27/a_125_78# sky130_fd_sc_hs__dfrbp_1_27/a_796_463# sky130_fd_sc_hs__dfrbp_1_27/a_910_118#
+ sky130_fd_sc_hs__dfrbp_1_27/a_1465_471# sky130_fd_sc_hs__dfrbp_1_27/a_832_118# sky130_fd_sc_hs__dfrbp_1_27/a_841_401#
+ sky130_fd_sc_hs__dfrbp_1_27/a_38_78# sky130_fd_sc_hs__dfrbp_1_27/a_1434_74# sky130_fd_sc_hs__dfrbp_1_27/a_706_463#
+ sky130_fd_sc_hs__dfrbp_1_27/a_319_360# sky130_fd_sc_hs__dfrbp_1_27/a_1624_74# sky130_fd_sc_hs__dfrbp_1
Xsky130_fd_sc_hs__dfrbp_1_16 DVSS DVDD sky130_fd_sc_hs__clkbuf_8_1/X DVDD DVSS sky130_fd_sc_hs__inv_4_71/A
+ sky130_fd_sc_hs__clkbuf_2_1/X sky130_fd_sc_hs__dfrbp_1_17/D sky130_fd_sc_hs__dfrbp_1_17/Q_N
+ sky130_fd_sc_hs__dfrbp_1_17/a_498_360# sky130_fd_sc_hs__dfrbp_1_17/a_1224_74# sky130_fd_sc_hs__dfrbp_1_17/a_2026_424#
+ sky130_fd_sc_hs__dfrbp_1_17/a_1482_48# sky130_fd_sc_hs__dfrbp_1_17/a_125_78# sky130_fd_sc_hs__dfrbp_1_17/a_796_463#
+ sky130_fd_sc_hs__dfrbp_1_17/a_910_118# sky130_fd_sc_hs__dfrbp_1_17/a_1465_471# sky130_fd_sc_hs__dfrbp_1_17/a_832_118#
+ sky130_fd_sc_hs__dfrbp_1_17/a_841_401# sky130_fd_sc_hs__dfrbp_1_17/a_38_78# sky130_fd_sc_hs__dfrbp_1_17/a_1434_74#
+ sky130_fd_sc_hs__dfrbp_1_17/a_706_463# sky130_fd_sc_hs__dfrbp_1_17/a_319_360# sky130_fd_sc_hs__dfrbp_1_17/a_1624_74#
+ sky130_fd_sc_hs__dfrbp_1
Xsky130_fd_sc_hs__a222oi_1_2 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nor2_1_33/Y sky130_fd_sc_hs__inv_4_45/A
+ sky130_fd_sc_hs__inv_4_41/A sky130_fd_sc_hs__nor2b_1_23/Y sky130_fd_sc_hs__inv_4_47/A
+ sky130_fd_sc_hs__a32oi_1_5/A1 sky130_fd_sc_hs__nor2b_1_25/Y sky130_fd_sc_hs__a222oi_1_3/a_461_74#
+ sky130_fd_sc_hs__a222oi_1_3/a_697_74# sky130_fd_sc_hs__a222oi_1_3/a_119_74# sky130_fd_sc_hs__a222oi_1_3/a_116_392#
+ sky130_fd_sc_hs__a222oi_1_3/a_369_392# sky130_fd_sc_hs__a222oi_1
Xsky130_fd_sc_hs__dfrbp_1_38 DVSS DVDD sky130_fd_sc_hs__clkbuf_8_1/X DVDD DVSS sky130_fd_sc_hs__o21a_1_75/A1
+ ref_clk sky130_fd_sc_hs__o21a_1_75/X sky130_fd_sc_hs__dfrbp_1_39/Q_N sky130_fd_sc_hs__dfrbp_1_39/a_498_360#
+ sky130_fd_sc_hs__dfrbp_1_39/a_1224_74# sky130_fd_sc_hs__dfrbp_1_39/a_2026_424# sky130_fd_sc_hs__dfrbp_1_39/a_1482_48#
+ sky130_fd_sc_hs__dfrbp_1_39/a_125_78# sky130_fd_sc_hs__dfrbp_1_39/a_796_463# sky130_fd_sc_hs__dfrbp_1_39/a_910_118#
+ sky130_fd_sc_hs__dfrbp_1_39/a_1465_471# sky130_fd_sc_hs__dfrbp_1_39/a_832_118# sky130_fd_sc_hs__dfrbp_1_39/a_841_401#
+ sky130_fd_sc_hs__dfrbp_1_39/a_38_78# sky130_fd_sc_hs__dfrbp_1_39/a_1434_74# sky130_fd_sc_hs__dfrbp_1_39/a_706_463#
+ sky130_fd_sc_hs__dfrbp_1_39/a_319_360# sky130_fd_sc_hs__dfrbp_1_39/a_1624_74# sky130_fd_sc_hs__dfrbp_1
Xsky130_fd_sc_hs__xor2_1_5 DVSS DVDD DVDD DVSS fine_con_step_size[2] sky130_fd_sc_hs__fa_2_9/B
+ sky130_fd_sc_hs__fa_2_3/A sky130_fd_sc_hs__xor2_1_5/a_194_125# sky130_fd_sc_hs__xor2_1_5/a_355_368#
+ sky130_fd_sc_hs__xor2_1_5/a_455_87# sky130_fd_sc_hs__xor2_1_5/a_158_392# sky130_fd_sc_hs__xor2_1
Xsky130_fd_sc_hs__o21ai_2_0 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__o21ai_2_1/B1 sky130_fd_sc_hs__inv_4_103/A
+ div_ratio_half[4] sky130_fd_sc_hs__inv_2_7/A sky130_fd_sc_hs__o21ai_2_1/a_116_368#
+ sky130_fd_sc_hs__o21ai_2_1/a_27_74# sky130_fd_sc_hs__o21ai_2
Xsky130_fd_sc_hs__a21oi_1_7 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nor2_1_9/Y sky130_fd_sc_hs__dfrtp_4_7/D
+ sky130_fd_sc_hs__nor2_1_9/B sky130_fd_sc_hs__inv_4_9/Y sky130_fd_sc_hs__a21oi_1_7/a_117_74#
+ sky130_fd_sc_hs__a21oi_1_7/a_29_368# sky130_fd_sc_hs__a21oi_1
Xsky130_fd_sc_hs__dfrtn_1_17 DVSS DVDD sky130_fd_sc_hs__clkbuf_8_1/X DVDD DVSS sky130_fd_sc_hs__clkbuf_2_1/X
+ sky130_fd_sc_hs__inv_4_63/A sky130_fd_sc_hs__dfrtn_1_17/D sky130_fd_sc_hs__dfrtn_1_17/a_1266_119#
+ sky130_fd_sc_hs__dfrtn_1_17/a_1736_119# sky130_fd_sc_hs__dfrtn_1_17/a_817_508# sky130_fd_sc_hs__dfrtn_1_17/a_120_74#
+ sky130_fd_sc_hs__dfrtn_1_17/a_1547_508# sky130_fd_sc_hs__dfrtn_1_17/a_922_127# sky130_fd_sc_hs__dfrtn_1_17/a_33_74#
+ sky130_fd_sc_hs__dfrtn_1_17/a_714_127# sky130_fd_sc_hs__dfrtn_1_17/a_1934_94# sky130_fd_sc_hs__dfrtn_1_17/a_1550_119#
+ sky130_fd_sc_hs__dfrtn_1_17/a_1598_93# sky130_fd_sc_hs__dfrtn_1_17/a_300_74# sky130_fd_sc_hs__dfrtn_1_17/a_507_368#
+ sky130_fd_sc_hs__dfrtn_1_17/a_856_304# sky130_fd_sc_hs__dfrtn_1_17/a_850_127# sky130_fd_sc_hs__dfrtn_1
Xsky130_fd_sc_hs__dfrtn_1_28 DVSS DVDD sky130_fd_sc_hs__clkbuf_8_1/X DVDD DVSS ref_clk
+ sky130_fd_sc_hs__o21a_1_59/A1 sky130_fd_sc_hs__o21a_1_59/X sky130_fd_sc_hs__dfrtn_1_29/a_1266_119#
+ sky130_fd_sc_hs__dfrtn_1_29/a_1736_119# sky130_fd_sc_hs__dfrtn_1_29/a_817_508# sky130_fd_sc_hs__dfrtn_1_29/a_120_74#
+ sky130_fd_sc_hs__dfrtn_1_29/a_1547_508# sky130_fd_sc_hs__dfrtn_1_29/a_922_127# sky130_fd_sc_hs__dfrtn_1_29/a_33_74#
+ sky130_fd_sc_hs__dfrtn_1_29/a_714_127# sky130_fd_sc_hs__dfrtn_1_29/a_1934_94# sky130_fd_sc_hs__dfrtn_1_29/a_1550_119#
+ sky130_fd_sc_hs__dfrtn_1_29/a_1598_93# sky130_fd_sc_hs__dfrtn_1_29/a_300_74# sky130_fd_sc_hs__dfrtn_1_29/a_507_368#
+ sky130_fd_sc_hs__dfrtn_1_29/a_856_304# sky130_fd_sc_hs__dfrtn_1_29/a_850_127# sky130_fd_sc_hs__dfrtn_1
Xsky130_fd_sc_hs__dfrtn_1_39 DVSS DVDD sky130_fd_sc_hs__clkbuf_8_1/X DVDD DVSS ref_clk
+ sky130_fd_sc_hs__inv_4_125/A sky130_fd_sc_hs__dfrtn_1_39/D sky130_fd_sc_hs__dfrtn_1_39/a_1266_119#
+ sky130_fd_sc_hs__dfrtn_1_39/a_1736_119# sky130_fd_sc_hs__dfrtn_1_39/a_817_508# sky130_fd_sc_hs__dfrtn_1_39/a_120_74#
+ sky130_fd_sc_hs__dfrtn_1_39/a_1547_508# sky130_fd_sc_hs__dfrtn_1_39/a_922_127# sky130_fd_sc_hs__dfrtn_1_39/a_33_74#
+ sky130_fd_sc_hs__dfrtn_1_39/a_714_127# sky130_fd_sc_hs__dfrtn_1_39/a_1934_94# sky130_fd_sc_hs__dfrtn_1_39/a_1550_119#
+ sky130_fd_sc_hs__dfrtn_1_39/a_1598_93# sky130_fd_sc_hs__dfrtn_1_39/a_300_74# sky130_fd_sc_hs__dfrtn_1_39/a_507_368#
+ sky130_fd_sc_hs__dfrtn_1_39/a_856_304# sky130_fd_sc_hs__dfrtn_1_39/a_850_127# sky130_fd_sc_hs__dfrtn_1
Xsky130_fd_sc_hs__xor2_1_10 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__xor2_1_9/X sky130_fd_sc_hs__xor2_1_11/B
+ sky130_fd_sc_hs__or2_1_1/B sky130_fd_sc_hs__xor2_1_11/a_194_125# sky130_fd_sc_hs__xor2_1_11/a_355_368#
+ sky130_fd_sc_hs__xor2_1_11/a_455_87# sky130_fd_sc_hs__xor2_1_11/a_158_392# sky130_fd_sc_hs__xor2_1
Xsky130_fd_sc_hs__nand2b_1_3 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_87/A sky130_fd_sc_hs__nor2_1_53/Y
+ sky130_fd_sc_hs__nand2b_1_3/Y sky130_fd_sc_hs__nand2b_1_3/a_269_74# sky130_fd_sc_hs__nand2b_1_3/a_27_112#
+ sky130_fd_sc_hs__nand2b_1
Xsky130_fd_sc_hs__dfrbp_1_5 DVSS DVDD sky130_fd_sc_hs__clkbuf_8_1/X DVDD DVSS sky130_fd_sc_hs__inv_4_51/A
+ sky130_fd_sc_hs__clkbuf_2_1/X sky130_fd_sc_hs__dfrbp_1_5/D sky130_fd_sc_hs__dfrbp_1_5/Q_N
+ sky130_fd_sc_hs__dfrbp_1_5/a_498_360# sky130_fd_sc_hs__dfrbp_1_5/a_1224_74# sky130_fd_sc_hs__dfrbp_1_5/a_2026_424#
+ sky130_fd_sc_hs__dfrbp_1_5/a_1482_48# sky130_fd_sc_hs__dfrbp_1_5/a_125_78# sky130_fd_sc_hs__dfrbp_1_5/a_796_463#
+ sky130_fd_sc_hs__dfrbp_1_5/a_910_118# sky130_fd_sc_hs__dfrbp_1_5/a_1465_471# sky130_fd_sc_hs__dfrbp_1_5/a_832_118#
+ sky130_fd_sc_hs__dfrbp_1_5/a_841_401# sky130_fd_sc_hs__dfrbp_1_5/a_38_78# sky130_fd_sc_hs__dfrbp_1_5/a_1434_74#
+ sky130_fd_sc_hs__dfrbp_1_5/a_706_463# sky130_fd_sc_hs__dfrbp_1_5/a_319_360# sky130_fd_sc_hs__dfrbp_1_5/a_1624_74#
+ sky130_fd_sc_hs__dfrbp_1
Xsky130_fd_sc_hs__a32oi_1_2 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_2_1/Y sky130_fd_sc_hs__inv_4_21/Y
+ sky130_fd_sc_hs__a32oi_1_3/B1 fine_control_avg_window_select[1] sky130_fd_sc_hs__a32oi_1_3/Y
+ sky130_fd_sc_hs__inv_4_27/Y sky130_fd_sc_hs__a32oi_1_3/a_391_74# sky130_fd_sc_hs__a32oi_1_3/a_27_368#
+ sky130_fd_sc_hs__a32oi_1_3/a_119_74# sky130_fd_sc_hs__a32oi_1_3/a_469_74# sky130_fd_sc_hs__a32oi_1
Xsky130_fd_sc_hs__dfrtn_1_3 DVSS DVDD sky130_fd_sc_hs__clkbuf_8_1/X DVDD DVSS sky130_fd_sc_hs__clkbuf_2_1/X
+ sky130_fd_sc_hs__inv_4_37/A sky130_fd_sc_hs__dfrtn_1_3/D sky130_fd_sc_hs__dfrtn_1_3/a_1266_119#
+ sky130_fd_sc_hs__dfrtn_1_3/a_1736_119# sky130_fd_sc_hs__dfrtn_1_3/a_817_508# sky130_fd_sc_hs__dfrtn_1_3/a_120_74#
+ sky130_fd_sc_hs__dfrtn_1_3/a_1547_508# sky130_fd_sc_hs__dfrtn_1_3/a_922_127# sky130_fd_sc_hs__dfrtn_1_3/a_33_74#
+ sky130_fd_sc_hs__dfrtn_1_3/a_714_127# sky130_fd_sc_hs__dfrtn_1_3/a_1934_94# sky130_fd_sc_hs__dfrtn_1_3/a_1550_119#
+ sky130_fd_sc_hs__dfrtn_1_3/a_1598_93# sky130_fd_sc_hs__dfrtn_1_3/a_300_74# sky130_fd_sc_hs__dfrtn_1_3/a_507_368#
+ sky130_fd_sc_hs__dfrtn_1_3/a_856_304# sky130_fd_sc_hs__dfrtn_1_3/a_850_127# sky130_fd_sc_hs__dfrtn_1
Xsky130_fd_sc_hs__o211ai_1_3 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__a21oi_1_82/Y sky130_fd_sc_hs__o211ai_1_3/Y
+ sky130_fd_sc_hs__nand4_1_5/A sky130_fd_sc_hs__a21oi_1_93/Y sky130_fd_sc_hs__nor3_1_1/A
+ sky130_fd_sc_hs__o211ai_1_3/a_31_74# sky130_fd_sc_hs__o211ai_1_3/a_311_74# sky130_fd_sc_hs__o211ai_1_3/a_116_368#
+ sky130_fd_sc_hs__o211ai_1
Xsky130_fd_sc_hs__inv_4_17 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_17/Y sky130_fd_sc_hs__inv_4_17/A
+ sky130_fd_sc_hs__inv_4
Xsky130_fd_sc_hs__a31oi_1_1 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__dfstp_2_7/D sky130_fd_sc_hs__nand2_1_71/Y
+ sky130_fd_sc_hs__nor4_1_1/A sky130_fd_sc_hs__a31oi_1_1/A2 sky130_fd_sc_hs__maj3_1_3/X
+ sky130_fd_sc_hs__a31oi_1_1/a_136_368# sky130_fd_sc_hs__a31oi_1_1/a_223_74# sky130_fd_sc_hs__a31oi_1_1/a_145_74#
+ sky130_fd_sc_hs__a31oi_1
Xsky130_fd_sc_hs__inv_4_39 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_39/Y sky130_fd_sc_hs__inv_4_39/A
+ sky130_fd_sc_hs__inv_4
Xsky130_fd_sc_hs__inv_4_28 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_29/Y sky130_fd_sc_hs__inv_4_29/A
+ sky130_fd_sc_hs__inv_4
Xsky130_fd_sc_hs__dfrtp_4_80 DVSS DVDD sky130_fd_sc_hs__clkbuf_8_1/X DVDD DVSS sky130_fd_sc_hs__o21a_1_43/X
+ sky130_fd_sc_hs__clkbuf_2_1/X sky130_fd_sc_hs__inv_4_73/A sky130_fd_sc_hs__dfrtp_4_81/a_37_78#
+ sky130_fd_sc_hs__dfrtp_4_81/a_494_366# sky130_fd_sc_hs__dfrtp_4_81/a_699_463# sky130_fd_sc_hs__dfrtp_4_81/a_313_74#
+ sky130_fd_sc_hs__dfrtp_4_81/a_1627_493# sky130_fd_sc_hs__dfrtp_4_81/a_1678_395#
+ sky130_fd_sc_hs__dfrtp_4_81/a_1827_81# sky130_fd_sc_hs__dfrtp_4_81/a_789_463# sky130_fd_sc_hs__dfrtp_4_81/a_1350_392#
+ sky130_fd_sc_hs__dfrtp_4_81/a_834_355# sky130_fd_sc_hs__dfrtp_4_81/a_812_138# sky130_fd_sc_hs__dfrtp_4_81/a_124_78#
+ sky130_fd_sc_hs__dfrtp_4_81/a_1647_81# sky130_fd_sc_hs__dfrtp_4_81/a_2010_409# sky130_fd_sc_hs__dfrtp_4_81/a_890_138#
+ sky130_fd_sc_hs__dfrtp_4
Xsky130_fd_sc_hs__a22o_1_2 DVSS DVDD DVDD DVSS osc_fine_con_final[2] manual_control_osc[2]
+ sky130_fd_sc_hs__inv_4_43/Y sky130_fd_sc_hs__fa_2_3/B fftl_en sky130_fd_sc_hs__a22o_1_3/a_222_392#
+ sky130_fd_sc_hs__a22o_1_3/a_230_79# sky130_fd_sc_hs__a22o_1_3/a_52_123# sky130_fd_sc_hs__a22o_1_3/a_132_392#
+ sky130_fd_sc_hs__a22o_1
Xsky130_fd_sc_hs__dfrtp_4_91 DVSS DVDD sky130_fd_sc_hs__inv_4_49/Y DVDD DVSS sky130_fd_sc_hs__nor2b_1_27/Y
+ sky130_fd_sc_hs__dfstp_2_1/CLK sky130_fd_sc_hs__fa_2_19/B sky130_fd_sc_hs__dfrtp_4_91/a_37_78#
+ sky130_fd_sc_hs__dfrtp_4_91/a_494_366# sky130_fd_sc_hs__dfrtp_4_91/a_699_463# sky130_fd_sc_hs__dfrtp_4_91/a_313_74#
+ sky130_fd_sc_hs__dfrtp_4_91/a_1627_493# sky130_fd_sc_hs__dfrtp_4_91/a_1678_395#
+ sky130_fd_sc_hs__dfrtp_4_91/a_1827_81# sky130_fd_sc_hs__dfrtp_4_91/a_789_463# sky130_fd_sc_hs__dfrtp_4_91/a_1350_392#
+ sky130_fd_sc_hs__dfrtp_4_91/a_834_355# sky130_fd_sc_hs__dfrtp_4_91/a_812_138# sky130_fd_sc_hs__dfrtp_4_91/a_124_78#
+ sky130_fd_sc_hs__dfrtp_4_91/a_1647_81# sky130_fd_sc_hs__dfrtp_4_91/a_2010_409# sky130_fd_sc_hs__dfrtp_4_91/a_890_138#
+ sky130_fd_sc_hs__dfrtp_4
Xsky130_fd_sc_hs__fa_2_5 DVSS DVDD sky130_fd_sc_hs__fa_2_5/A DVDD DVSS sky130_fd_sc_hs__fa_2_5/CIN
+ sky130_fd_sc_hs__fa_2_5/B sky130_fd_sc_hs__fa_2_3/CIN sky130_fd_sc_hs__fa_2_5/SUM
+ sky130_fd_sc_hs__fa_2_5/a_27_378# sky130_fd_sc_hs__fa_2_5/a_701_79# sky130_fd_sc_hs__fa_2_5/a_484_347#
+ sky130_fd_sc_hs__fa_2_5/a_1094_347# sky130_fd_sc_hs__fa_2_5/a_1205_79# sky130_fd_sc_hs__fa_2_5/a_27_79#
+ sky130_fd_sc_hs__fa_2_5/a_1202_368# sky130_fd_sc_hs__fa_2_5/a_336_347# sky130_fd_sc_hs__fa_2_5/a_992_347#
+ sky130_fd_sc_hs__fa_2_5/a_1119_79# sky130_fd_sc_hs__fa_2_5/a_487_79# sky130_fd_sc_hs__fa_2_5/a_683_347#
+ sky130_fd_sc_hs__fa_2
Xsky130_fd_sc_hs__nor3_1_9 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nor3_1_9/Y sky130_fd_sc_hs__nor3_1_9/C
+ sky130_fd_sc_hs__nor3_1_9/B sky130_fd_sc_hs__nor3_1_9/A sky130_fd_sc_hs__nor3_1_9/a_198_368#
+ sky130_fd_sc_hs__nor3_1_9/a_114_368# sky130_fd_sc_hs__nor3_1
Xsky130_fd_sc_hs__nor2b_1_0 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__fa_2_1/SUM sky130_fd_sc_hs__nor2b_1_1/Y
+ sky130_fd_sc_hs__or2_1_1/A sky130_fd_sc_hs__nor2b_1_1/a_278_368# sky130_fd_sc_hs__nor2b_1_1/a_27_112#
+ sky130_fd_sc_hs__nor2b_1
Xsky130_fd_sc_hs__nand2_1_2 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nor2_1_5/Y sky130_fd_sc_hs__nor2_1_7/B
+ sky130_fd_sc_hs__o21a_1_1/A1 sky130_fd_sc_hs__nand2_1_3/a_117_74# sky130_fd_sc_hs__nand2_1
Xsky130_fd_sc_hs__a22oi_1_9 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nor2b_1_25/Y sky130_fd_sc_hs__nand2_2_3/A
+ sky130_fd_sc_hs__o21a_1_17/A1 sky130_fd_sc_hs__nor2b_1_23/Y sky130_fd_sc_hs__o21a_1_7/A1
+ sky130_fd_sc_hs__a22oi_1_9/a_71_368# sky130_fd_sc_hs__a22oi_1_9/a_159_74# sky130_fd_sc_hs__a22oi_1_9/a_339_74#
+ sky130_fd_sc_hs__a22oi_1
Xsky130_fd_sc_hs__a21oi_1_83 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nor3_1_5/B sky130_fd_sc_hs__o31ai_1_3/B1
+ sky130_fd_sc_hs__nor4_1_3/A sky130_fd_sc_hs__a21oi_1_82/Y sky130_fd_sc_hs__a21oi_1_83/a_117_74#
+ sky130_fd_sc_hs__a21oi_1_83/a_29_368# sky130_fd_sc_hs__a21oi_1
Xsky130_fd_sc_hs__a21oi_1_72 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nor2_1_75/Y sky130_fd_sc_hs__dfrtn_1_19/D
+ sky130_fd_sc_hs__nor2_1_75/B sky130_fd_sc_hs__inv_4_75/Y sky130_fd_sc_hs__a21oi_1_73/a_117_74#
+ sky130_fd_sc_hs__a21oi_1_73/a_29_368# sky130_fd_sc_hs__a21oi_1
Xsky130_fd_sc_hs__a21oi_1_61 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__a22o_1_27/X sky130_fd_sc_hs__o21ai_1_5/B1
+ sky130_fd_sc_hs__inv_4_55/Y sky130_fd_sc_hs__nor2_1_59/A sky130_fd_sc_hs__a21oi_1_61/a_117_74#
+ sky130_fd_sc_hs__a21oi_1_61/a_29_368# sky130_fd_sc_hs__a21oi_1
Xsky130_fd_sc_hs__a21oi_1_50 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nor2_1_41/Y sky130_fd_sc_hs__dfrbp_1_5/D
+ sky130_fd_sc_hs__nor2_1_41/B sky130_fd_sc_hs__inv_4_51/Y sky130_fd_sc_hs__a21oi_1_51/a_117_74#
+ sky130_fd_sc_hs__a21oi_1_51/a_29_368# sky130_fd_sc_hs__a21oi_1
Xsky130_fd_sc_hs__a21oi_1_94 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nor4_1_3/D sky130_fd_sc_hs__o31ai_1_7/A1
+ sky130_fd_sc_hs__or2_1_3/X sky130_fd_sc_hs__a22oi_1_23/Y sky130_fd_sc_hs__a21oi_1_95/a_117_74#
+ sky130_fd_sc_hs__a21oi_1_95/a_29_368# sky130_fd_sc_hs__a21oi_1
Xsky130_fd_sc_hs__dfrbp_1_17 DVSS DVDD sky130_fd_sc_hs__clkbuf_8_1/X DVDD DVSS sky130_fd_sc_hs__inv_4_71/A
+ sky130_fd_sc_hs__clkbuf_2_1/X sky130_fd_sc_hs__dfrbp_1_17/D sky130_fd_sc_hs__dfrbp_1_17/Q_N
+ sky130_fd_sc_hs__dfrbp_1_17/a_498_360# sky130_fd_sc_hs__dfrbp_1_17/a_1224_74# sky130_fd_sc_hs__dfrbp_1_17/a_2026_424#
+ sky130_fd_sc_hs__dfrbp_1_17/a_1482_48# sky130_fd_sc_hs__dfrbp_1_17/a_125_78# sky130_fd_sc_hs__dfrbp_1_17/a_796_463#
+ sky130_fd_sc_hs__dfrbp_1_17/a_910_118# sky130_fd_sc_hs__dfrbp_1_17/a_1465_471# sky130_fd_sc_hs__dfrbp_1_17/a_832_118#
+ sky130_fd_sc_hs__dfrbp_1_17/a_841_401# sky130_fd_sc_hs__dfrbp_1_17/a_38_78# sky130_fd_sc_hs__dfrbp_1_17/a_1434_74#
+ sky130_fd_sc_hs__dfrbp_1_17/a_706_463# sky130_fd_sc_hs__dfrbp_1_17/a_319_360# sky130_fd_sc_hs__dfrbp_1_17/a_1624_74#
+ sky130_fd_sc_hs__dfrbp_1
Xsky130_fd_sc_hs__a222oi_1_3 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nor2_1_33/Y sky130_fd_sc_hs__inv_4_45/A
+ sky130_fd_sc_hs__inv_4_41/A sky130_fd_sc_hs__nor2b_1_23/Y sky130_fd_sc_hs__inv_4_47/A
+ sky130_fd_sc_hs__a32oi_1_5/A1 sky130_fd_sc_hs__nor2b_1_25/Y sky130_fd_sc_hs__a222oi_1_3/a_461_74#
+ sky130_fd_sc_hs__a222oi_1_3/a_697_74# sky130_fd_sc_hs__a222oi_1_3/a_119_74# sky130_fd_sc_hs__a222oi_1_3/a_116_392#
+ sky130_fd_sc_hs__a222oi_1_3/a_369_392# sky130_fd_sc_hs__a222oi_1
Xsky130_fd_sc_hs__dfrbp_1_28 DVSS DVDD sky130_fd_sc_hs__clkbuf_8_1/X DVDD DVSS sky130_fd_sc_hs__nor2_1_97/A
+ ref_clk sky130_fd_sc_hs__dfrbp_1_29/D sky130_fd_sc_hs__dfrbp_1_29/Q_N sky130_fd_sc_hs__dfrbp_1_29/a_498_360#
+ sky130_fd_sc_hs__dfrbp_1_29/a_1224_74# sky130_fd_sc_hs__dfrbp_1_29/a_2026_424# sky130_fd_sc_hs__dfrbp_1_29/a_1482_48#
+ sky130_fd_sc_hs__dfrbp_1_29/a_125_78# sky130_fd_sc_hs__dfrbp_1_29/a_796_463# sky130_fd_sc_hs__dfrbp_1_29/a_910_118#
+ sky130_fd_sc_hs__dfrbp_1_29/a_1465_471# sky130_fd_sc_hs__dfrbp_1_29/a_832_118# sky130_fd_sc_hs__dfrbp_1_29/a_841_401#
+ sky130_fd_sc_hs__dfrbp_1_29/a_38_78# sky130_fd_sc_hs__dfrbp_1_29/a_1434_74# sky130_fd_sc_hs__dfrbp_1_29/a_706_463#
+ sky130_fd_sc_hs__dfrbp_1_29/a_319_360# sky130_fd_sc_hs__dfrbp_1_29/a_1624_74# sky130_fd_sc_hs__dfrbp_1
Xsky130_fd_sc_hs__dfrbp_1_39 DVSS DVDD sky130_fd_sc_hs__clkbuf_8_1/X DVDD DVSS sky130_fd_sc_hs__o21a_1_75/A1
+ ref_clk sky130_fd_sc_hs__o21a_1_75/X sky130_fd_sc_hs__dfrbp_1_39/Q_N sky130_fd_sc_hs__dfrbp_1_39/a_498_360#
+ sky130_fd_sc_hs__dfrbp_1_39/a_1224_74# sky130_fd_sc_hs__dfrbp_1_39/a_2026_424# sky130_fd_sc_hs__dfrbp_1_39/a_1482_48#
+ sky130_fd_sc_hs__dfrbp_1_39/a_125_78# sky130_fd_sc_hs__dfrbp_1_39/a_796_463# sky130_fd_sc_hs__dfrbp_1_39/a_910_118#
+ sky130_fd_sc_hs__dfrbp_1_39/a_1465_471# sky130_fd_sc_hs__dfrbp_1_39/a_832_118# sky130_fd_sc_hs__dfrbp_1_39/a_841_401#
+ sky130_fd_sc_hs__dfrbp_1_39/a_38_78# sky130_fd_sc_hs__dfrbp_1_39/a_1434_74# sky130_fd_sc_hs__dfrbp_1_39/a_706_463#
+ sky130_fd_sc_hs__dfrbp_1_39/a_319_360# sky130_fd_sc_hs__dfrbp_1_39/a_1624_74# sky130_fd_sc_hs__dfrbp_1
Xsky130_fd_sc_hs__xor2_1_6 DVSS DVDD DVDD DVSS fine_con_step_size[3] sky130_fd_sc_hs__fa_2_9/B
+ sky130_fd_sc_hs__fa_2_1/A sky130_fd_sc_hs__xor2_1_7/a_194_125# sky130_fd_sc_hs__xor2_1_7/a_355_368#
+ sky130_fd_sc_hs__xor2_1_7/a_455_87# sky130_fd_sc_hs__xor2_1_7/a_158_392# sky130_fd_sc_hs__xor2_1
Xsky130_fd_sc_hs__o21ai_2_1 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__o21ai_2_1/B1 sky130_fd_sc_hs__inv_4_103/A
+ div_ratio_half[4] sky130_fd_sc_hs__inv_2_7/A sky130_fd_sc_hs__o21ai_2_1/a_116_368#
+ sky130_fd_sc_hs__o21ai_2_1/a_27_74# sky130_fd_sc_hs__o21ai_2
Xsky130_fd_sc_hs__a21oi_1_8 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nor2_1_7/Y sky130_fd_sc_hs__a21oi_1_9/Y
+ sky130_fd_sc_hs__nor2_1_7/B sky130_fd_sc_hs__nor2_1_7/A sky130_fd_sc_hs__a21oi_1_9/a_117_74#
+ sky130_fd_sc_hs__a21oi_1_9/a_29_368# sky130_fd_sc_hs__a21oi_1
Xsky130_fd_sc_hs__dfrtn_1_18 DVSS DVDD sky130_fd_sc_hs__clkbuf_8_1/X DVDD DVSS sky130_fd_sc_hs__clkbuf_2_1/X
+ sky130_fd_sc_hs__inv_4_75/A sky130_fd_sc_hs__dfrtn_1_19/D sky130_fd_sc_hs__dfrtn_1_19/a_1266_119#
+ sky130_fd_sc_hs__dfrtn_1_19/a_1736_119# sky130_fd_sc_hs__dfrtn_1_19/a_817_508# sky130_fd_sc_hs__dfrtn_1_19/a_120_74#
+ sky130_fd_sc_hs__dfrtn_1_19/a_1547_508# sky130_fd_sc_hs__dfrtn_1_19/a_922_127# sky130_fd_sc_hs__dfrtn_1_19/a_33_74#
+ sky130_fd_sc_hs__dfrtn_1_19/a_714_127# sky130_fd_sc_hs__dfrtn_1_19/a_1934_94# sky130_fd_sc_hs__dfrtn_1_19/a_1550_119#
+ sky130_fd_sc_hs__dfrtn_1_19/a_1598_93# sky130_fd_sc_hs__dfrtn_1_19/a_300_74# sky130_fd_sc_hs__dfrtn_1_19/a_507_368#
+ sky130_fd_sc_hs__dfrtn_1_19/a_856_304# sky130_fd_sc_hs__dfrtn_1_19/a_850_127# sky130_fd_sc_hs__dfrtn_1
Xsky130_fd_sc_hs__dfrtn_1_29 DVSS DVDD sky130_fd_sc_hs__clkbuf_8_1/X DVDD DVSS ref_clk
+ sky130_fd_sc_hs__o21a_1_59/A1 sky130_fd_sc_hs__o21a_1_59/X sky130_fd_sc_hs__dfrtn_1_29/a_1266_119#
+ sky130_fd_sc_hs__dfrtn_1_29/a_1736_119# sky130_fd_sc_hs__dfrtn_1_29/a_817_508# sky130_fd_sc_hs__dfrtn_1_29/a_120_74#
+ sky130_fd_sc_hs__dfrtn_1_29/a_1547_508# sky130_fd_sc_hs__dfrtn_1_29/a_922_127# sky130_fd_sc_hs__dfrtn_1_29/a_33_74#
+ sky130_fd_sc_hs__dfrtn_1_29/a_714_127# sky130_fd_sc_hs__dfrtn_1_29/a_1934_94# sky130_fd_sc_hs__dfrtn_1_29/a_1550_119#
+ sky130_fd_sc_hs__dfrtn_1_29/a_1598_93# sky130_fd_sc_hs__dfrtn_1_29/a_300_74# sky130_fd_sc_hs__dfrtn_1_29/a_507_368#
+ sky130_fd_sc_hs__dfrtn_1_29/a_856_304# sky130_fd_sc_hs__dfrtn_1_29/a_850_127# sky130_fd_sc_hs__dfrtn_1
Xsky130_fd_sc_hs__xor2_1_11 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__xor2_1_9/X sky130_fd_sc_hs__xor2_1_11/B
+ sky130_fd_sc_hs__or2_1_1/B sky130_fd_sc_hs__xor2_1_11/a_194_125# sky130_fd_sc_hs__xor2_1_11/a_355_368#
+ sky130_fd_sc_hs__xor2_1_11/a_455_87# sky130_fd_sc_hs__xor2_1_11/a_158_392# sky130_fd_sc_hs__xor2_1
Xsky130_fd_sc_hs__nand2b_1_4 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__xnor2_1_3/Y sky130_fd_sc_hs__inv_4_91/A
+ sky130_fd_sc_hs__nor2_2_1/A sky130_fd_sc_hs__nand2b_1_5/a_269_74# sky130_fd_sc_hs__nand2b_1_5/a_27_112#
+ sky130_fd_sc_hs__nand2b_1
Xsky130_fd_sc_hs__dfrbp_1_6 DVSS DVDD sky130_fd_sc_hs__clkbuf_8_1/X DVDD DVSS sky130_fd_sc_hs__dfrbp_1_7/Q
+ sky130_fd_sc_hs__clkbuf_2_1/X sky130_fd_sc_hs__o21a_1_41/X sky130_fd_sc_hs__dfrbp_1_7/Q_N
+ sky130_fd_sc_hs__dfrbp_1_7/a_498_360# sky130_fd_sc_hs__dfrbp_1_7/a_1224_74# sky130_fd_sc_hs__dfrbp_1_7/a_2026_424#
+ sky130_fd_sc_hs__dfrbp_1_7/a_1482_48# sky130_fd_sc_hs__dfrbp_1_7/a_125_78# sky130_fd_sc_hs__dfrbp_1_7/a_796_463#
+ sky130_fd_sc_hs__dfrbp_1_7/a_910_118# sky130_fd_sc_hs__dfrbp_1_7/a_1465_471# sky130_fd_sc_hs__dfrbp_1_7/a_832_118#
+ sky130_fd_sc_hs__dfrbp_1_7/a_841_401# sky130_fd_sc_hs__dfrbp_1_7/a_38_78# sky130_fd_sc_hs__dfrbp_1_7/a_1434_74#
+ sky130_fd_sc_hs__dfrbp_1_7/a_706_463# sky130_fd_sc_hs__dfrbp_1_7/a_319_360# sky130_fd_sc_hs__dfrbp_1_7/a_1624_74#
+ sky130_fd_sc_hs__dfrbp_1
Xsky130_fd_sc_hs__a32oi_1_3 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_2_1/Y sky130_fd_sc_hs__inv_4_21/Y
+ sky130_fd_sc_hs__a32oi_1_3/B1 fine_control_avg_window_select[1] sky130_fd_sc_hs__a32oi_1_3/Y
+ sky130_fd_sc_hs__inv_4_27/Y sky130_fd_sc_hs__a32oi_1_3/a_391_74# sky130_fd_sc_hs__a32oi_1_3/a_27_368#
+ sky130_fd_sc_hs__a32oi_1_3/a_119_74# sky130_fd_sc_hs__a32oi_1_3/a_469_74# sky130_fd_sc_hs__a32oi_1
Xsky130_fd_sc_hs__dfrtn_1_4 DVSS DVDD sky130_fd_sc_hs__clkbuf_8_1/X DVDD DVSS sky130_fd_sc_hs__clkbuf_2_1/X
+ sky130_fd_sc_hs__inv_4_55/A sky130_fd_sc_hs__o21a_1_33/X sky130_fd_sc_hs__dfrtn_1_5/a_1266_119#
+ sky130_fd_sc_hs__dfrtn_1_5/a_1736_119# sky130_fd_sc_hs__dfrtn_1_5/a_817_508# sky130_fd_sc_hs__dfrtn_1_5/a_120_74#
+ sky130_fd_sc_hs__dfrtn_1_5/a_1547_508# sky130_fd_sc_hs__dfrtn_1_5/a_922_127# sky130_fd_sc_hs__dfrtn_1_5/a_33_74#
+ sky130_fd_sc_hs__dfrtn_1_5/a_714_127# sky130_fd_sc_hs__dfrtn_1_5/a_1934_94# sky130_fd_sc_hs__dfrtn_1_5/a_1550_119#
+ sky130_fd_sc_hs__dfrtn_1_5/a_1598_93# sky130_fd_sc_hs__dfrtn_1_5/a_300_74# sky130_fd_sc_hs__dfrtn_1_5/a_507_368#
+ sky130_fd_sc_hs__dfrtn_1_5/a_856_304# sky130_fd_sc_hs__dfrtn_1_5/a_850_127# sky130_fd_sc_hs__dfrtn_1
Xsky130_fd_sc_hs__o211ai_1_4 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__maj3_1_3/C sky130_fd_sc_hs__o211ai_1_5/Y
+ sky130_fd_sc_hs__nand2_1_71/Y sky130_fd_sc_hs__maj3_1_1/C sky130_fd_sc_hs__maj3_1_1/A
+ sky130_fd_sc_hs__o211ai_1_5/a_31_74# sky130_fd_sc_hs__o211ai_1_5/a_311_74# sky130_fd_sc_hs__o211ai_1_5/a_116_368#
+ sky130_fd_sc_hs__o211ai_1
Xsky130_fd_sc_hs__inv_4_29 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_29/Y sky130_fd_sc_hs__inv_4_29/A
+ sky130_fd_sc_hs__inv_4
Xsky130_fd_sc_hs__inv_4_18 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_19/Y sky130_fd_sc_hs__inv_4_19/A
+ sky130_fd_sc_hs__inv_4
Xsky130_fd_sc_hs__dfrtp_4_70 DVSS DVDD sky130_fd_sc_hs__inv_4_49/Y DVDD DVSS sky130_fd_sc_hs__nor2b_1_19/Y
+ sky130_fd_sc_hs__dfstp_2_1/CLK sky130_fd_sc_hs__fa_2_21/B sky130_fd_sc_hs__dfrtp_4_71/a_37_78#
+ sky130_fd_sc_hs__dfrtp_4_71/a_494_366# sky130_fd_sc_hs__dfrtp_4_71/a_699_463# sky130_fd_sc_hs__dfrtp_4_71/a_313_74#
+ sky130_fd_sc_hs__dfrtp_4_71/a_1627_493# sky130_fd_sc_hs__dfrtp_4_71/a_1678_395#
+ sky130_fd_sc_hs__dfrtp_4_71/a_1827_81# sky130_fd_sc_hs__dfrtp_4_71/a_789_463# sky130_fd_sc_hs__dfrtp_4_71/a_1350_392#
+ sky130_fd_sc_hs__dfrtp_4_71/a_834_355# sky130_fd_sc_hs__dfrtp_4_71/a_812_138# sky130_fd_sc_hs__dfrtp_4_71/a_124_78#
+ sky130_fd_sc_hs__dfrtp_4_71/a_1647_81# sky130_fd_sc_hs__dfrtp_4_71/a_2010_409# sky130_fd_sc_hs__dfrtp_4_71/a_890_138#
+ sky130_fd_sc_hs__dfrtp_4
Xsky130_fd_sc_hs__a22o_1_3 DVSS DVDD DVDD DVSS osc_fine_con_final[2] manual_control_osc[2]
+ sky130_fd_sc_hs__inv_4_43/Y sky130_fd_sc_hs__fa_2_3/B fftl_en sky130_fd_sc_hs__a22o_1_3/a_222_392#
+ sky130_fd_sc_hs__a22o_1_3/a_230_79# sky130_fd_sc_hs__a22o_1_3/a_52_123# sky130_fd_sc_hs__a22o_1_3/a_132_392#
+ sky130_fd_sc_hs__a22o_1
Xsky130_fd_sc_hs__dfrtp_4_81 DVSS DVDD sky130_fd_sc_hs__clkbuf_8_1/X DVDD DVSS sky130_fd_sc_hs__o21a_1_43/X
+ sky130_fd_sc_hs__clkbuf_2_1/X sky130_fd_sc_hs__inv_4_73/A sky130_fd_sc_hs__dfrtp_4_81/a_37_78#
+ sky130_fd_sc_hs__dfrtp_4_81/a_494_366# sky130_fd_sc_hs__dfrtp_4_81/a_699_463# sky130_fd_sc_hs__dfrtp_4_81/a_313_74#
+ sky130_fd_sc_hs__dfrtp_4_81/a_1627_493# sky130_fd_sc_hs__dfrtp_4_81/a_1678_395#
+ sky130_fd_sc_hs__dfrtp_4_81/a_1827_81# sky130_fd_sc_hs__dfrtp_4_81/a_789_463# sky130_fd_sc_hs__dfrtp_4_81/a_1350_392#
+ sky130_fd_sc_hs__dfrtp_4_81/a_834_355# sky130_fd_sc_hs__dfrtp_4_81/a_812_138# sky130_fd_sc_hs__dfrtp_4_81/a_124_78#
+ sky130_fd_sc_hs__dfrtp_4_81/a_1647_81# sky130_fd_sc_hs__dfrtp_4_81/a_2010_409# sky130_fd_sc_hs__dfrtp_4_81/a_890_138#
+ sky130_fd_sc_hs__dfrtp_4
Xsky130_fd_sc_hs__fa_2_6 DVSS DVDD sky130_fd_sc_hs__fa_2_9/B DVDD DVSS sky130_fd_sc_hs__fa_2_7/CIN
+ sky130_fd_sc_hs__fa_2_7/B sky130_fd_sc_hs__fa_2_7/COUT sky130_fd_sc_hs__fa_2_7/SUM
+ sky130_fd_sc_hs__fa_2_7/a_27_378# sky130_fd_sc_hs__fa_2_7/a_701_79# sky130_fd_sc_hs__fa_2_7/a_484_347#
+ sky130_fd_sc_hs__fa_2_7/a_1094_347# sky130_fd_sc_hs__fa_2_7/a_1205_79# sky130_fd_sc_hs__fa_2_7/a_27_79#
+ sky130_fd_sc_hs__fa_2_7/a_1202_368# sky130_fd_sc_hs__fa_2_7/a_336_347# sky130_fd_sc_hs__fa_2_7/a_992_347#
+ sky130_fd_sc_hs__fa_2_7/a_1119_79# sky130_fd_sc_hs__fa_2_7/a_487_79# sky130_fd_sc_hs__fa_2_7/a_683_347#
+ sky130_fd_sc_hs__fa_2
Xsky130_fd_sc_hs__nor2b_1_1 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__fa_2_1/SUM sky130_fd_sc_hs__nor2b_1_1/Y
+ sky130_fd_sc_hs__or2_1_1/A sky130_fd_sc_hs__nor2b_1_1/a_278_368# sky130_fd_sc_hs__nor2b_1_1/a_27_112#
+ sky130_fd_sc_hs__nor2b_1
Xsky130_fd_sc_hs__nand2_1_3 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nor2_1_5/Y sky130_fd_sc_hs__nor2_1_7/B
+ sky130_fd_sc_hs__o21a_1_1/A1 sky130_fd_sc_hs__nand2_1_3/a_117_74# sky130_fd_sc_hs__nand2_1
Xsky130_fd_sc_hs__a21oi_1_40 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nor2_1_29/Y sky130_fd_sc_hs__dfrtn_1_7/D
+ sky130_fd_sc_hs__nor2_1_29/B sky130_fd_sc_hs__inv_4_53/Y sky130_fd_sc_hs__a21oi_1_41/a_117_74#
+ sky130_fd_sc_hs__a21oi_1_41/a_29_368# sky130_fd_sc_hs__a21oi_1
Xsky130_fd_sc_hs__a21oi_1_73 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nor2_1_75/Y sky130_fd_sc_hs__dfrtn_1_19/D
+ sky130_fd_sc_hs__nor2_1_75/B sky130_fd_sc_hs__inv_4_75/Y sky130_fd_sc_hs__a21oi_1_73/a_117_74#
+ sky130_fd_sc_hs__a21oi_1_73/a_29_368# sky130_fd_sc_hs__a21oi_1
Xsky130_fd_sc_hs__a21oi_1_62 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nor2_1_43/Y sky130_fd_sc_hs__dfrbp_1_15/D
+ sky130_fd_sc_hs__nor2_1_43/B sky130_fd_sc_hs__inv_4_67/Y sky130_fd_sc_hs__a21oi_1_63/a_117_74#
+ sky130_fd_sc_hs__a21oi_1_63/a_29_368# sky130_fd_sc_hs__a21oi_1
Xsky130_fd_sc_hs__a21oi_1_51 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nor2_1_41/Y sky130_fd_sc_hs__dfrbp_1_5/D
+ sky130_fd_sc_hs__nor2_1_41/B sky130_fd_sc_hs__inv_4_51/Y sky130_fd_sc_hs__a21oi_1_51/a_117_74#
+ sky130_fd_sc_hs__a21oi_1_51/a_29_368# sky130_fd_sc_hs__a21oi_1
Xsky130_fd_sc_hs__a21oi_1_95 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nor4_1_3/D sky130_fd_sc_hs__o31ai_1_7/A1
+ sky130_fd_sc_hs__or2_1_3/X sky130_fd_sc_hs__a22oi_1_23/Y sky130_fd_sc_hs__a21oi_1_95/a_117_74#
+ sky130_fd_sc_hs__a21oi_1_95/a_29_368# sky130_fd_sc_hs__a21oi_1
Xsky130_fd_sc_hs__a21oi_1_84 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nor2_1_83/Y sky130_fd_sc_hs__dfrbp_1_19/D
+ sky130_fd_sc_hs__nor2_1_83/B sky130_fd_sc_hs__inv_4_89/Y sky130_fd_sc_hs__a21oi_1_85/a_117_74#
+ sky130_fd_sc_hs__a21oi_1_85/a_29_368# sky130_fd_sc_hs__a21oi_1
Xsky130_fd_sc_hs__dfrbp_1_18 DVSS DVDD sky130_fd_sc_hs__clkbuf_8_1/X DVDD DVSS sky130_fd_sc_hs__inv_4_89/A
+ sky130_fd_sc_hs__clkbuf_2_1/X sky130_fd_sc_hs__dfrbp_1_19/D sky130_fd_sc_hs__dfrbp_1_19/Q_N
+ sky130_fd_sc_hs__dfrbp_1_19/a_498_360# sky130_fd_sc_hs__dfrbp_1_19/a_1224_74# sky130_fd_sc_hs__dfrbp_1_19/a_2026_424#
+ sky130_fd_sc_hs__dfrbp_1_19/a_1482_48# sky130_fd_sc_hs__dfrbp_1_19/a_125_78# sky130_fd_sc_hs__dfrbp_1_19/a_796_463#
+ sky130_fd_sc_hs__dfrbp_1_19/a_910_118# sky130_fd_sc_hs__dfrbp_1_19/a_1465_471# sky130_fd_sc_hs__dfrbp_1_19/a_832_118#
+ sky130_fd_sc_hs__dfrbp_1_19/a_841_401# sky130_fd_sc_hs__dfrbp_1_19/a_38_78# sky130_fd_sc_hs__dfrbp_1_19/a_1434_74#
+ sky130_fd_sc_hs__dfrbp_1_19/a_706_463# sky130_fd_sc_hs__dfrbp_1_19/a_319_360# sky130_fd_sc_hs__dfrbp_1_19/a_1624_74#
+ sky130_fd_sc_hs__dfrbp_1
Xsky130_fd_sc_hs__dfrbp_1_29 DVSS DVDD sky130_fd_sc_hs__clkbuf_8_1/X DVDD DVSS sky130_fd_sc_hs__nor2_1_97/A
+ ref_clk sky130_fd_sc_hs__dfrbp_1_29/D sky130_fd_sc_hs__dfrbp_1_29/Q_N sky130_fd_sc_hs__dfrbp_1_29/a_498_360#
+ sky130_fd_sc_hs__dfrbp_1_29/a_1224_74# sky130_fd_sc_hs__dfrbp_1_29/a_2026_424# sky130_fd_sc_hs__dfrbp_1_29/a_1482_48#
+ sky130_fd_sc_hs__dfrbp_1_29/a_125_78# sky130_fd_sc_hs__dfrbp_1_29/a_796_463# sky130_fd_sc_hs__dfrbp_1_29/a_910_118#
+ sky130_fd_sc_hs__dfrbp_1_29/a_1465_471# sky130_fd_sc_hs__dfrbp_1_29/a_832_118# sky130_fd_sc_hs__dfrbp_1_29/a_841_401#
+ sky130_fd_sc_hs__dfrbp_1_29/a_38_78# sky130_fd_sc_hs__dfrbp_1_29/a_1434_74# sky130_fd_sc_hs__dfrbp_1_29/a_706_463#
+ sky130_fd_sc_hs__dfrbp_1_29/a_319_360# sky130_fd_sc_hs__dfrbp_1_29/a_1624_74# sky130_fd_sc_hs__dfrbp_1
Xsky130_fd_sc_hs__xor2_1_7 DVSS DVDD DVDD DVSS fine_con_step_size[3] sky130_fd_sc_hs__fa_2_9/B
+ sky130_fd_sc_hs__fa_2_1/A sky130_fd_sc_hs__xor2_1_7/a_194_125# sky130_fd_sc_hs__xor2_1_7/a_355_368#
+ sky130_fd_sc_hs__xor2_1_7/a_455_87# sky130_fd_sc_hs__xor2_1_7/a_158_392# sky130_fd_sc_hs__xor2_1
Xsky130_fd_sc_hs__a21oi_1_9 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nor2_1_7/Y sky130_fd_sc_hs__a21oi_1_9/Y
+ sky130_fd_sc_hs__nor2_1_7/B sky130_fd_sc_hs__nor2_1_7/A sky130_fd_sc_hs__a21oi_1_9/a_117_74#
+ sky130_fd_sc_hs__a21oi_1_9/a_29_368# sky130_fd_sc_hs__a21oi_1
Xsky130_fd_sc_hs__dfrtn_1_19 DVSS DVDD sky130_fd_sc_hs__clkbuf_8_1/X DVDD DVSS sky130_fd_sc_hs__clkbuf_2_1/X
+ sky130_fd_sc_hs__inv_4_75/A sky130_fd_sc_hs__dfrtn_1_19/D sky130_fd_sc_hs__dfrtn_1_19/a_1266_119#
+ sky130_fd_sc_hs__dfrtn_1_19/a_1736_119# sky130_fd_sc_hs__dfrtn_1_19/a_817_508# sky130_fd_sc_hs__dfrtn_1_19/a_120_74#
+ sky130_fd_sc_hs__dfrtn_1_19/a_1547_508# sky130_fd_sc_hs__dfrtn_1_19/a_922_127# sky130_fd_sc_hs__dfrtn_1_19/a_33_74#
+ sky130_fd_sc_hs__dfrtn_1_19/a_714_127# sky130_fd_sc_hs__dfrtn_1_19/a_1934_94# sky130_fd_sc_hs__dfrtn_1_19/a_1550_119#
+ sky130_fd_sc_hs__dfrtn_1_19/a_1598_93# sky130_fd_sc_hs__dfrtn_1_19/a_300_74# sky130_fd_sc_hs__dfrtn_1_19/a_507_368#
+ sky130_fd_sc_hs__dfrtn_1_19/a_856_304# sky130_fd_sc_hs__dfrtn_1_19/a_850_127# sky130_fd_sc_hs__dfrtn_1
Xsky130_fd_sc_hs__nand2b_1_5 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__xnor2_1_3/Y sky130_fd_sc_hs__inv_4_91/A
+ sky130_fd_sc_hs__nor2_2_1/A sky130_fd_sc_hs__nand2b_1_5/a_269_74# sky130_fd_sc_hs__nand2b_1_5/a_27_112#
+ sky130_fd_sc_hs__nand2b_1
Xsky130_fd_sc_hs__dfrbp_1_7 DVSS DVDD sky130_fd_sc_hs__clkbuf_8_1/X DVDD DVSS sky130_fd_sc_hs__dfrbp_1_7/Q
+ sky130_fd_sc_hs__clkbuf_2_1/X sky130_fd_sc_hs__o21a_1_41/X sky130_fd_sc_hs__dfrbp_1_7/Q_N
+ sky130_fd_sc_hs__dfrbp_1_7/a_498_360# sky130_fd_sc_hs__dfrbp_1_7/a_1224_74# sky130_fd_sc_hs__dfrbp_1_7/a_2026_424#
+ sky130_fd_sc_hs__dfrbp_1_7/a_1482_48# sky130_fd_sc_hs__dfrbp_1_7/a_125_78# sky130_fd_sc_hs__dfrbp_1_7/a_796_463#
+ sky130_fd_sc_hs__dfrbp_1_7/a_910_118# sky130_fd_sc_hs__dfrbp_1_7/a_1465_471# sky130_fd_sc_hs__dfrbp_1_7/a_832_118#
+ sky130_fd_sc_hs__dfrbp_1_7/a_841_401# sky130_fd_sc_hs__dfrbp_1_7/a_38_78# sky130_fd_sc_hs__dfrbp_1_7/a_1434_74#
+ sky130_fd_sc_hs__dfrbp_1_7/a_706_463# sky130_fd_sc_hs__dfrbp_1_7/a_319_360# sky130_fd_sc_hs__dfrbp_1_7/a_1624_74#
+ sky130_fd_sc_hs__dfrbp_1
Xsky130_fd_sc_hs__a32oi_1_4 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_25/A sky130_fd_sc_hs__o31ai_1_1/B1
+ sky130_fd_sc_hs__o22ai_1_1/A2 sky130_fd_sc_hs__o31ai_1_1/B1 sky130_fd_sc_hs__a32oi_1_5/Y
+ sky130_fd_sc_hs__a32oi_1_5/A1 sky130_fd_sc_hs__a32oi_1_5/a_391_74# sky130_fd_sc_hs__a32oi_1_5/a_27_368#
+ sky130_fd_sc_hs__a32oi_1_5/a_119_74# sky130_fd_sc_hs__a32oi_1_5/a_469_74# sky130_fd_sc_hs__a32oi_1
Xsky130_fd_sc_hs__o21a_1_0 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__o21a_1_1/X sky130_fd_sc_hs__nor2_1_5/Y
+ sky130_fd_sc_hs__nor2_1_7/B sky130_fd_sc_hs__o21a_1_1/A1 sky130_fd_sc_hs__o21a_1_1/a_320_74#
+ sky130_fd_sc_hs__o21a_1_1/a_376_387# sky130_fd_sc_hs__o21a_1_1/a_83_244# sky130_fd_sc_hs__o21a_1
Xsky130_fd_sc_hs__dfrtn_1_5 DVSS DVDD sky130_fd_sc_hs__clkbuf_8_1/X DVDD DVSS sky130_fd_sc_hs__clkbuf_2_1/X
+ sky130_fd_sc_hs__inv_4_55/A sky130_fd_sc_hs__o21a_1_33/X sky130_fd_sc_hs__dfrtn_1_5/a_1266_119#
+ sky130_fd_sc_hs__dfrtn_1_5/a_1736_119# sky130_fd_sc_hs__dfrtn_1_5/a_817_508# sky130_fd_sc_hs__dfrtn_1_5/a_120_74#
+ sky130_fd_sc_hs__dfrtn_1_5/a_1547_508# sky130_fd_sc_hs__dfrtn_1_5/a_922_127# sky130_fd_sc_hs__dfrtn_1_5/a_33_74#
+ sky130_fd_sc_hs__dfrtn_1_5/a_714_127# sky130_fd_sc_hs__dfrtn_1_5/a_1934_94# sky130_fd_sc_hs__dfrtn_1_5/a_1550_119#
+ sky130_fd_sc_hs__dfrtn_1_5/a_1598_93# sky130_fd_sc_hs__dfrtn_1_5/a_300_74# sky130_fd_sc_hs__dfrtn_1_5/a_507_368#
+ sky130_fd_sc_hs__dfrtn_1_5/a_856_304# sky130_fd_sc_hs__dfrtn_1_5/a_850_127# sky130_fd_sc_hs__dfrtn_1
Xsky130_fd_sc_hs__o211ai_1_5 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__maj3_1_3/C sky130_fd_sc_hs__o211ai_1_5/Y
+ sky130_fd_sc_hs__nand2_1_71/Y sky130_fd_sc_hs__maj3_1_1/C sky130_fd_sc_hs__maj3_1_1/A
+ sky130_fd_sc_hs__o211ai_1_5/a_31_74# sky130_fd_sc_hs__o211ai_1_5/a_311_74# sky130_fd_sc_hs__o211ai_1_5/a_116_368#
+ sky130_fd_sc_hs__o211ai_1
Xsky130_fd_sc_hs__nand3b_2_0 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nor2_1_91/B rst
+ sky130_fd_sc_hs__inv_4_91/A sky130_fd_sc_hs__inv_4_87/Y sky130_fd_sc_hs__nand3b_2_1/a_27_94#
+ sky130_fd_sc_hs__nand3b_2_1/a_403_54# sky130_fd_sc_hs__nand3b_2_1/a_206_74# sky130_fd_sc_hs__nand3b_2
Xsky130_fd_sc_hs__inv_4_19 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_19/Y sky130_fd_sc_hs__inv_4_19/A
+ sky130_fd_sc_hs__inv_4
Xsky130_fd_sc_hs__o21a_1_70 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__o21a_1_71/X sky130_fd_sc_hs__o21a_1_71/A2
+ sky130_fd_sc_hs__o21a_1_71/B1 sky130_fd_sc_hs__o21a_1_71/A1 sky130_fd_sc_hs__o21a_1_71/a_320_74#
+ sky130_fd_sc_hs__o21a_1_71/a_376_387# sky130_fd_sc_hs__o21a_1_71/a_83_244# sky130_fd_sc_hs__o21a_1
Xsky130_fd_sc_hs__dfrtp_4_71 DVSS DVDD sky130_fd_sc_hs__inv_4_49/Y DVDD DVSS sky130_fd_sc_hs__nor2b_1_19/Y
+ sky130_fd_sc_hs__dfstp_2_1/CLK sky130_fd_sc_hs__fa_2_21/B sky130_fd_sc_hs__dfrtp_4_71/a_37_78#
+ sky130_fd_sc_hs__dfrtp_4_71/a_494_366# sky130_fd_sc_hs__dfrtp_4_71/a_699_463# sky130_fd_sc_hs__dfrtp_4_71/a_313_74#
+ sky130_fd_sc_hs__dfrtp_4_71/a_1627_493# sky130_fd_sc_hs__dfrtp_4_71/a_1678_395#
+ sky130_fd_sc_hs__dfrtp_4_71/a_1827_81# sky130_fd_sc_hs__dfrtp_4_71/a_789_463# sky130_fd_sc_hs__dfrtp_4_71/a_1350_392#
+ sky130_fd_sc_hs__dfrtp_4_71/a_834_355# sky130_fd_sc_hs__dfrtp_4_71/a_812_138# sky130_fd_sc_hs__dfrtp_4_71/a_124_78#
+ sky130_fd_sc_hs__dfrtp_4_71/a_1647_81# sky130_fd_sc_hs__dfrtp_4_71/a_2010_409# sky130_fd_sc_hs__dfrtp_4_71/a_890_138#
+ sky130_fd_sc_hs__dfrtp_4
Xsky130_fd_sc_hs__dfrtp_4_60 DVSS DVDD sky130_fd_sc_hs__inv_4_49/Y DVDD DVSS sky130_fd_sc_hs__nor2b_1_13/Y
+ sky130_fd_sc_hs__dfstp_2_1/CLK sky130_fd_sc_hs__fa_2_13/B sky130_fd_sc_hs__dfrtp_4_61/a_37_78#
+ sky130_fd_sc_hs__dfrtp_4_61/a_494_366# sky130_fd_sc_hs__dfrtp_4_61/a_699_463# sky130_fd_sc_hs__dfrtp_4_61/a_313_74#
+ sky130_fd_sc_hs__dfrtp_4_61/a_1627_493# sky130_fd_sc_hs__dfrtp_4_61/a_1678_395#
+ sky130_fd_sc_hs__dfrtp_4_61/a_1827_81# sky130_fd_sc_hs__dfrtp_4_61/a_789_463# sky130_fd_sc_hs__dfrtp_4_61/a_1350_392#
+ sky130_fd_sc_hs__dfrtp_4_61/a_834_355# sky130_fd_sc_hs__dfrtp_4_61/a_812_138# sky130_fd_sc_hs__dfrtp_4_61/a_124_78#
+ sky130_fd_sc_hs__dfrtp_4_61/a_1647_81# sky130_fd_sc_hs__dfrtp_4_61/a_2010_409# sky130_fd_sc_hs__dfrtp_4_61/a_890_138#
+ sky130_fd_sc_hs__dfrtp_4
Xsky130_fd_sc_hs__dfrtp_4_82 DVSS DVDD sky130_fd_sc_hs__clkbuf_8_1/X DVDD DVSS sky130_fd_sc_hs__dfrtp_4_83/D
+ sky130_fd_sc_hs__nand2_1_47/B sky130_fd_sc_hs__inv_4_45/A sky130_fd_sc_hs__dfrtp_4_83/a_37_78#
+ sky130_fd_sc_hs__dfrtp_4_83/a_494_366# sky130_fd_sc_hs__dfrtp_4_83/a_699_463# sky130_fd_sc_hs__dfrtp_4_83/a_313_74#
+ sky130_fd_sc_hs__dfrtp_4_83/a_1627_493# sky130_fd_sc_hs__dfrtp_4_83/a_1678_395#
+ sky130_fd_sc_hs__dfrtp_4_83/a_1827_81# sky130_fd_sc_hs__dfrtp_4_83/a_789_463# sky130_fd_sc_hs__dfrtp_4_83/a_1350_392#
+ sky130_fd_sc_hs__dfrtp_4_83/a_834_355# sky130_fd_sc_hs__dfrtp_4_83/a_812_138# sky130_fd_sc_hs__dfrtp_4_83/a_124_78#
+ sky130_fd_sc_hs__dfrtp_4_83/a_1647_81# sky130_fd_sc_hs__dfrtp_4_83/a_2010_409# sky130_fd_sc_hs__dfrtp_4_83/a_890_138#
+ sky130_fd_sc_hs__dfrtp_4
Xsky130_fd_sc_hs__a22o_1_4 DVSS DVDD DVDD DVSS osc_fine_con_final[1] manual_control_osc[1]
+ sky130_fd_sc_hs__inv_4_43/Y sky130_fd_sc_hs__fa_2_5/B fftl_en sky130_fd_sc_hs__a22o_1_5/a_222_392#
+ sky130_fd_sc_hs__a22o_1_5/a_230_79# sky130_fd_sc_hs__a22o_1_5/a_52_123# sky130_fd_sc_hs__a22o_1_5/a_132_392#
+ sky130_fd_sc_hs__a22o_1
Xsky130_fd_sc_hs__fa_2_7 DVSS DVDD sky130_fd_sc_hs__fa_2_9/B DVDD DVSS sky130_fd_sc_hs__fa_2_7/CIN
+ sky130_fd_sc_hs__fa_2_7/B sky130_fd_sc_hs__fa_2_7/COUT sky130_fd_sc_hs__fa_2_7/SUM
+ sky130_fd_sc_hs__fa_2_7/a_27_378# sky130_fd_sc_hs__fa_2_7/a_701_79# sky130_fd_sc_hs__fa_2_7/a_484_347#
+ sky130_fd_sc_hs__fa_2_7/a_1094_347# sky130_fd_sc_hs__fa_2_7/a_1205_79# sky130_fd_sc_hs__fa_2_7/a_27_79#
+ sky130_fd_sc_hs__fa_2_7/a_1202_368# sky130_fd_sc_hs__fa_2_7/a_336_347# sky130_fd_sc_hs__fa_2_7/a_992_347#
+ sky130_fd_sc_hs__fa_2_7/a_1119_79# sky130_fd_sc_hs__fa_2_7/a_487_79# sky130_fd_sc_hs__fa_2_7/a_683_347#
+ sky130_fd_sc_hs__fa_2
Xsky130_fd_sc_hs__nor2b_1_2 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__fa_2_3/SUM sky130_fd_sc_hs__nor2b_1_3/Y
+ sky130_fd_sc_hs__or2_1_1/A sky130_fd_sc_hs__nor2b_1_3/a_278_368# sky130_fd_sc_hs__nor2b_1_3/a_27_112#
+ sky130_fd_sc_hs__nor2b_1
Xsky130_fd_sc_hs__nand2_1_4 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nor2_1_3/Y sky130_fd_sc_hs__o21a_1_5/B1
+ sky130_fd_sc_hs__o21a_1_5/A1 sky130_fd_sc_hs__nand2_1_5/a_117_74# sky130_fd_sc_hs__nand2_1
Xsky130_fd_sc_hs__nor2_1_0 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_1/Y sky130_fd_sc_hs__nor2_1_1/Y
+ sky130_fd_sc_hs__inv_4_5/Y sky130_fd_sc_hs__nor2_1_1/a_116_368# sky130_fd_sc_hs__nor2_1
Xsky130_fd_sc_hs__a21oi_1_30 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__o21a_1_7/A2 sky130_fd_sc_hs__dfrtp_4_57/D
+ sky130_fd_sc_hs__nor2_1_19/B sky130_fd_sc_hs__inv_4_29/Y sky130_fd_sc_hs__a21oi_1_31/a_117_74#
+ sky130_fd_sc_hs__a21oi_1_31/a_29_368# sky130_fd_sc_hs__a21oi_1
Xsky130_fd_sc_hs__a21oi_1_74 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__o22ai_1_9/Y sky130_fd_sc_hs__a31oi_1_1/A2
+ sky130_fd_sc_hs__inv_4_77/Y sky130_fd_sc_hs__a31oi_2_1/Y sky130_fd_sc_hs__a21oi_1_75/a_117_74#
+ sky130_fd_sc_hs__a21oi_1_75/a_29_368# sky130_fd_sc_hs__a21oi_1
Xsky130_fd_sc_hs__a21oi_1_63 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nor2_1_43/Y sky130_fd_sc_hs__dfrbp_1_15/D
+ sky130_fd_sc_hs__nor2_1_43/B sky130_fd_sc_hs__inv_4_67/Y sky130_fd_sc_hs__a21oi_1_63/a_117_74#
+ sky130_fd_sc_hs__a21oi_1_63/a_29_368# sky130_fd_sc_hs__a21oi_1
Xsky130_fd_sc_hs__a21oi_1_52 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nor2_1_35/Y sky130_fd_sc_hs__dfrtp_4_85/D
+ sky130_fd_sc_hs__nor2_1_35/B sky130_fd_sc_hs__inv_4_47/Y sky130_fd_sc_hs__a21oi_1_53/a_117_74#
+ sky130_fd_sc_hs__a21oi_1_53/a_29_368# sky130_fd_sc_hs__a21oi_1
Xsky130_fd_sc_hs__a21oi_1_41 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nor2_1_29/Y sky130_fd_sc_hs__dfrtn_1_7/D
+ sky130_fd_sc_hs__nor2_1_29/B sky130_fd_sc_hs__inv_4_53/Y sky130_fd_sc_hs__a21oi_1_41/a_117_74#
+ sky130_fd_sc_hs__a21oi_1_41/a_29_368# sky130_fd_sc_hs__a21oi_1
Xsky130_fd_sc_hs__a21oi_1_96 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__a22o_1_29/X sky130_fd_sc_hs__a21oi_1_97/Y
+ sky130_fd_sc_hs__or2_1_3/B sky130_fd_sc_hs__or2_1_3/A sky130_fd_sc_hs__a21oi_1_97/a_117_74#
+ sky130_fd_sc_hs__a21oi_1_97/a_29_368# sky130_fd_sc_hs__a21oi_1
Xsky130_fd_sc_hs__a21oi_1_85 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nor2_1_83/Y sky130_fd_sc_hs__dfrbp_1_19/D
+ sky130_fd_sc_hs__nor2_1_83/B sky130_fd_sc_hs__inv_4_89/Y sky130_fd_sc_hs__a21oi_1_85/a_117_74#
+ sky130_fd_sc_hs__a21oi_1_85/a_29_368# sky130_fd_sc_hs__a21oi_1
Xsky130_fd_sc_hs__dfrbp_1_19 DVSS DVDD sky130_fd_sc_hs__clkbuf_8_1/X DVDD DVSS sky130_fd_sc_hs__inv_4_89/A
+ sky130_fd_sc_hs__clkbuf_2_1/X sky130_fd_sc_hs__dfrbp_1_19/D sky130_fd_sc_hs__dfrbp_1_19/Q_N
+ sky130_fd_sc_hs__dfrbp_1_19/a_498_360# sky130_fd_sc_hs__dfrbp_1_19/a_1224_74# sky130_fd_sc_hs__dfrbp_1_19/a_2026_424#
+ sky130_fd_sc_hs__dfrbp_1_19/a_1482_48# sky130_fd_sc_hs__dfrbp_1_19/a_125_78# sky130_fd_sc_hs__dfrbp_1_19/a_796_463#
+ sky130_fd_sc_hs__dfrbp_1_19/a_910_118# sky130_fd_sc_hs__dfrbp_1_19/a_1465_471# sky130_fd_sc_hs__dfrbp_1_19/a_832_118#
+ sky130_fd_sc_hs__dfrbp_1_19/a_841_401# sky130_fd_sc_hs__dfrbp_1_19/a_38_78# sky130_fd_sc_hs__dfrbp_1_19/a_1434_74#
+ sky130_fd_sc_hs__dfrbp_1_19/a_706_463# sky130_fd_sc_hs__dfrbp_1_19/a_319_360# sky130_fd_sc_hs__dfrbp_1_19/a_1624_74#
+ sky130_fd_sc_hs__dfrbp_1
Xsky130_fd_sc_hs__xor2_1_8 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__xor2_1_9/A sky130_fd_sc_hs__fa_2_9/B
+ sky130_fd_sc_hs__xor2_1_9/X sky130_fd_sc_hs__xor2_1_9/a_194_125# sky130_fd_sc_hs__xor2_1_9/a_355_368#
+ sky130_fd_sc_hs__xor2_1_9/a_455_87# sky130_fd_sc_hs__xor2_1_9/a_158_392# sky130_fd_sc_hs__xor2_1
Xsky130_fd_sc_hs__nand2b_1_6 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__xnor2_1_7/B sky130_fd_sc_hs__nor3_1_7/Y
+ sky130_fd_sc_hs__nor2_1_89/A sky130_fd_sc_hs__nand2b_1_7/a_269_74# sky130_fd_sc_hs__nand2b_1_7/a_27_112#
+ sky130_fd_sc_hs__nand2b_1
Xsky130_fd_sc_hs__dfrbp_1_8 DVSS DVDD sky130_fd_sc_hs__clkbuf_8_1/X DVDD DVSS sky130_fd_sc_hs__inv_4_69/A
+ sky130_fd_sc_hs__clkbuf_2_1/X sky130_fd_sc_hs__o21a_1_45/X sky130_fd_sc_hs__dfrbp_1_9/Q_N
+ sky130_fd_sc_hs__dfrbp_1_9/a_498_360# sky130_fd_sc_hs__dfrbp_1_9/a_1224_74# sky130_fd_sc_hs__dfrbp_1_9/a_2026_424#
+ sky130_fd_sc_hs__dfrbp_1_9/a_1482_48# sky130_fd_sc_hs__dfrbp_1_9/a_125_78# sky130_fd_sc_hs__dfrbp_1_9/a_796_463#
+ sky130_fd_sc_hs__dfrbp_1_9/a_910_118# sky130_fd_sc_hs__dfrbp_1_9/a_1465_471# sky130_fd_sc_hs__dfrbp_1_9/a_832_118#
+ sky130_fd_sc_hs__dfrbp_1_9/a_841_401# sky130_fd_sc_hs__dfrbp_1_9/a_38_78# sky130_fd_sc_hs__dfrbp_1_9/a_1434_74#
+ sky130_fd_sc_hs__dfrbp_1_9/a_706_463# sky130_fd_sc_hs__dfrbp_1_9/a_319_360# sky130_fd_sc_hs__dfrbp_1_9/a_1624_74#
+ sky130_fd_sc_hs__dfrbp_1
Xsky130_fd_sc_hs__a32oi_1_5 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_25/A sky130_fd_sc_hs__o31ai_1_1/B1
+ sky130_fd_sc_hs__o22ai_1_1/A2 sky130_fd_sc_hs__o31ai_1_1/B1 sky130_fd_sc_hs__a32oi_1_5/Y
+ sky130_fd_sc_hs__a32oi_1_5/A1 sky130_fd_sc_hs__a32oi_1_5/a_391_74# sky130_fd_sc_hs__a32oi_1_5/a_27_368#
+ sky130_fd_sc_hs__a32oi_1_5/a_119_74# sky130_fd_sc_hs__a32oi_1_5/a_469_74# sky130_fd_sc_hs__a32oi_1
Xsky130_fd_sc_hs__o21a_1_1 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__o21a_1_1/X sky130_fd_sc_hs__nor2_1_5/Y
+ sky130_fd_sc_hs__nor2_1_7/B sky130_fd_sc_hs__o21a_1_1/A1 sky130_fd_sc_hs__o21a_1_1/a_320_74#
+ sky130_fd_sc_hs__o21a_1_1/a_376_387# sky130_fd_sc_hs__o21a_1_1/a_83_244# sky130_fd_sc_hs__o21a_1
Xsky130_fd_sc_hs__fa_2_20 DVSS DVDD sky130_fd_sc_hs__fa_2_9/B DVDD DVSS sky130_fd_sc_hs__fa_2_21/CIN
+ sky130_fd_sc_hs__fa_2_21/B sky130_fd_sc_hs__fa_2_23/CIN sky130_fd_sc_hs__fa_2_21/SUM
+ sky130_fd_sc_hs__fa_2_21/a_27_378# sky130_fd_sc_hs__fa_2_21/a_701_79# sky130_fd_sc_hs__fa_2_21/a_484_347#
+ sky130_fd_sc_hs__fa_2_21/a_1094_347# sky130_fd_sc_hs__fa_2_21/a_1205_79# sky130_fd_sc_hs__fa_2_21/a_27_79#
+ sky130_fd_sc_hs__fa_2_21/a_1202_368# sky130_fd_sc_hs__fa_2_21/a_336_347# sky130_fd_sc_hs__fa_2_21/a_992_347#
+ sky130_fd_sc_hs__fa_2_21/a_1119_79# sky130_fd_sc_hs__fa_2_21/a_487_79# sky130_fd_sc_hs__fa_2_21/a_683_347#
+ sky130_fd_sc_hs__fa_2
Xsky130_fd_sc_hs__dfrtn_1_6 DVSS DVDD sky130_fd_sc_hs__clkbuf_8_1/X DVDD DVSS sky130_fd_sc_hs__clkbuf_2_1/X
+ sky130_fd_sc_hs__inv_4_53/A sky130_fd_sc_hs__dfrtn_1_7/D sky130_fd_sc_hs__dfrtn_1_7/a_1266_119#
+ sky130_fd_sc_hs__dfrtn_1_7/a_1736_119# sky130_fd_sc_hs__dfrtn_1_7/a_817_508# sky130_fd_sc_hs__dfrtn_1_7/a_120_74#
+ sky130_fd_sc_hs__dfrtn_1_7/a_1547_508# sky130_fd_sc_hs__dfrtn_1_7/a_922_127# sky130_fd_sc_hs__dfrtn_1_7/a_33_74#
+ sky130_fd_sc_hs__dfrtn_1_7/a_714_127# sky130_fd_sc_hs__dfrtn_1_7/a_1934_94# sky130_fd_sc_hs__dfrtn_1_7/a_1550_119#
+ sky130_fd_sc_hs__dfrtn_1_7/a_1598_93# sky130_fd_sc_hs__dfrtn_1_7/a_300_74# sky130_fd_sc_hs__dfrtn_1_7/a_507_368#
+ sky130_fd_sc_hs__dfrtn_1_7/a_856_304# sky130_fd_sc_hs__dfrtn_1_7/a_850_127# sky130_fd_sc_hs__dfrtn_1
Xsky130_fd_sc_hs__o211ai_1_6 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__a21oi_1_97/Y sky130_fd_sc_hs__nor3_1_3/A
+ sky130_fd_sc_hs__nor2_1_61/Y sky130_fd_sc_hs__maj3_1_3/B sky130_fd_sc_hs__maj3_1_3/A
+ sky130_fd_sc_hs__o211ai_1_7/a_31_74# sky130_fd_sc_hs__o211ai_1_7/a_311_74# sky130_fd_sc_hs__o211ai_1_7/a_116_368#
+ sky130_fd_sc_hs__o211ai_1
Xsky130_fd_sc_hs__nand3b_2_1 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nor2_1_91/B rst
+ sky130_fd_sc_hs__inv_4_91/A sky130_fd_sc_hs__inv_4_87/Y sky130_fd_sc_hs__nand3b_2_1/a_27_94#
+ sky130_fd_sc_hs__nand3b_2_1/a_403_54# sky130_fd_sc_hs__nand3b_2_1/a_206_74# sky130_fd_sc_hs__nand3b_2
Xsky130_fd_sc_hs__o21a_1_60 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__o21a_1_61/X sky130_fd_sc_hs__o21a_1_61/A2
+ sky130_fd_sc_hs__xnor2_1_5/B sky130_fd_sc_hs__maj3_1_3/A sky130_fd_sc_hs__o21a_1_61/a_320_74#
+ sky130_fd_sc_hs__o21a_1_61/a_376_387# sky130_fd_sc_hs__o21a_1_61/a_83_244# sky130_fd_sc_hs__o21a_1
Xsky130_fd_sc_hs__o21a_1_71 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__o21a_1_71/X sky130_fd_sc_hs__o21a_1_71/A2
+ sky130_fd_sc_hs__o21a_1_71/B1 sky130_fd_sc_hs__o21a_1_71/A1 sky130_fd_sc_hs__o21a_1_71/a_320_74#
+ sky130_fd_sc_hs__o21a_1_71/a_376_387# sky130_fd_sc_hs__o21a_1_71/a_83_244# sky130_fd_sc_hs__o21a_1
Xsky130_fd_sc_hs__dfrtp_4_61 DVSS DVDD sky130_fd_sc_hs__inv_4_49/Y DVDD DVSS sky130_fd_sc_hs__nor2b_1_13/Y
+ sky130_fd_sc_hs__dfstp_2_1/CLK sky130_fd_sc_hs__fa_2_13/B sky130_fd_sc_hs__dfrtp_4_61/a_37_78#
+ sky130_fd_sc_hs__dfrtp_4_61/a_494_366# sky130_fd_sc_hs__dfrtp_4_61/a_699_463# sky130_fd_sc_hs__dfrtp_4_61/a_313_74#
+ sky130_fd_sc_hs__dfrtp_4_61/a_1627_493# sky130_fd_sc_hs__dfrtp_4_61/a_1678_395#
+ sky130_fd_sc_hs__dfrtp_4_61/a_1827_81# sky130_fd_sc_hs__dfrtp_4_61/a_789_463# sky130_fd_sc_hs__dfrtp_4_61/a_1350_392#
+ sky130_fd_sc_hs__dfrtp_4_61/a_834_355# sky130_fd_sc_hs__dfrtp_4_61/a_812_138# sky130_fd_sc_hs__dfrtp_4_61/a_124_78#
+ sky130_fd_sc_hs__dfrtp_4_61/a_1647_81# sky130_fd_sc_hs__dfrtp_4_61/a_2010_409# sky130_fd_sc_hs__dfrtp_4_61/a_890_138#
+ sky130_fd_sc_hs__dfrtp_4
Xsky130_fd_sc_hs__dfrtp_4_50 DVSS DVDD sky130_fd_sc_hs__clkbuf_8_1/X DVDD DVSS sky130_fd_sc_hs__o21a_1_13/X
+ sky130_fd_sc_hs__nand2_1_47/B sky130_fd_sc_hs__o21a_1_13/A1 sky130_fd_sc_hs__dfrtp_4_51/a_37_78#
+ sky130_fd_sc_hs__dfrtp_4_51/a_494_366# sky130_fd_sc_hs__dfrtp_4_51/a_699_463# sky130_fd_sc_hs__dfrtp_4_51/a_313_74#
+ sky130_fd_sc_hs__dfrtp_4_51/a_1627_493# sky130_fd_sc_hs__dfrtp_4_51/a_1678_395#
+ sky130_fd_sc_hs__dfrtp_4_51/a_1827_81# sky130_fd_sc_hs__dfrtp_4_51/a_789_463# sky130_fd_sc_hs__dfrtp_4_51/a_1350_392#
+ sky130_fd_sc_hs__dfrtp_4_51/a_834_355# sky130_fd_sc_hs__dfrtp_4_51/a_812_138# sky130_fd_sc_hs__dfrtp_4_51/a_124_78#
+ sky130_fd_sc_hs__dfrtp_4_51/a_1647_81# sky130_fd_sc_hs__dfrtp_4_51/a_2010_409# sky130_fd_sc_hs__dfrtp_4_51/a_890_138#
+ sky130_fd_sc_hs__dfrtp_4
Xsky130_fd_sc_hs__dfrtp_4_83 DVSS DVDD sky130_fd_sc_hs__clkbuf_8_1/X DVDD DVSS sky130_fd_sc_hs__dfrtp_4_83/D
+ sky130_fd_sc_hs__nand2_1_47/B sky130_fd_sc_hs__inv_4_45/A sky130_fd_sc_hs__dfrtp_4_83/a_37_78#
+ sky130_fd_sc_hs__dfrtp_4_83/a_494_366# sky130_fd_sc_hs__dfrtp_4_83/a_699_463# sky130_fd_sc_hs__dfrtp_4_83/a_313_74#
+ sky130_fd_sc_hs__dfrtp_4_83/a_1627_493# sky130_fd_sc_hs__dfrtp_4_83/a_1678_395#
+ sky130_fd_sc_hs__dfrtp_4_83/a_1827_81# sky130_fd_sc_hs__dfrtp_4_83/a_789_463# sky130_fd_sc_hs__dfrtp_4_83/a_1350_392#
+ sky130_fd_sc_hs__dfrtp_4_83/a_834_355# sky130_fd_sc_hs__dfrtp_4_83/a_812_138# sky130_fd_sc_hs__dfrtp_4_83/a_124_78#
+ sky130_fd_sc_hs__dfrtp_4_83/a_1647_81# sky130_fd_sc_hs__dfrtp_4_83/a_2010_409# sky130_fd_sc_hs__dfrtp_4_83/a_890_138#
+ sky130_fd_sc_hs__dfrtp_4
Xsky130_fd_sc_hs__dfrtp_4_72 DVSS DVDD sky130_fd_sc_hs__inv_4_49/Y DVDD DVSS sky130_fd_sc_hs__nor2b_1_21/Y
+ sky130_fd_sc_hs__dfstp_2_1/CLK sky130_fd_sc_hs__fa_2_23/B sky130_fd_sc_hs__dfrtp_4_73/a_37_78#
+ sky130_fd_sc_hs__dfrtp_4_73/a_494_366# sky130_fd_sc_hs__dfrtp_4_73/a_699_463# sky130_fd_sc_hs__dfrtp_4_73/a_313_74#
+ sky130_fd_sc_hs__dfrtp_4_73/a_1627_493# sky130_fd_sc_hs__dfrtp_4_73/a_1678_395#
+ sky130_fd_sc_hs__dfrtp_4_73/a_1827_81# sky130_fd_sc_hs__dfrtp_4_73/a_789_463# sky130_fd_sc_hs__dfrtp_4_73/a_1350_392#
+ sky130_fd_sc_hs__dfrtp_4_73/a_834_355# sky130_fd_sc_hs__dfrtp_4_73/a_812_138# sky130_fd_sc_hs__dfrtp_4_73/a_124_78#
+ sky130_fd_sc_hs__dfrtp_4_73/a_1647_81# sky130_fd_sc_hs__dfrtp_4_73/a_2010_409# sky130_fd_sc_hs__dfrtp_4_73/a_890_138#
+ sky130_fd_sc_hs__dfrtp_4
Xsky130_fd_sc_hs__a22o_1_5 DVSS DVDD DVDD DVSS osc_fine_con_final[1] manual_control_osc[1]
+ sky130_fd_sc_hs__inv_4_43/Y sky130_fd_sc_hs__fa_2_5/B fftl_en sky130_fd_sc_hs__a22o_1_5/a_222_392#
+ sky130_fd_sc_hs__a22o_1_5/a_230_79# sky130_fd_sc_hs__a22o_1_5/a_52_123# sky130_fd_sc_hs__a22o_1_5/a_132_392#
+ sky130_fd_sc_hs__a22o_1
Xsky130_fd_sc_hs__fa_2_8 DVSS DVDD sky130_fd_sc_hs__fa_2_9/A DVDD DVSS sky130_fd_sc_hs__xor2_1_1/X
+ sky130_fd_sc_hs__fa_2_9/B sky130_fd_sc_hs__fa_2_5/CIN sky130_fd_sc_hs__fa_2_9/SUM
+ sky130_fd_sc_hs__fa_2_9/a_27_378# sky130_fd_sc_hs__fa_2_9/a_701_79# sky130_fd_sc_hs__fa_2_9/a_484_347#
+ sky130_fd_sc_hs__fa_2_9/a_1094_347# sky130_fd_sc_hs__fa_2_9/a_1205_79# sky130_fd_sc_hs__fa_2_9/a_27_79#
+ sky130_fd_sc_hs__fa_2_9/a_1202_368# sky130_fd_sc_hs__fa_2_9/a_336_347# sky130_fd_sc_hs__fa_2_9/a_992_347#
+ sky130_fd_sc_hs__fa_2_9/a_1119_79# sky130_fd_sc_hs__fa_2_9/a_487_79# sky130_fd_sc_hs__fa_2_9/a_683_347#
+ sky130_fd_sc_hs__fa_2
Xsky130_fd_sc_hs__o2bb2ai_1_0 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nor4_1_3/B sky130_fd_sc_hs__inv_4_73/Y
+ sky130_fd_sc_hs__inv_4_83/Y sky130_fd_sc_hs__nor2_1_65/A sky130_fd_sc_hs__dfrbp_1_7/Q
+ sky130_fd_sc_hs__o2bb2ai_1_1/a_114_74# sky130_fd_sc_hs__o2bb2ai_1_1/a_490_368# sky130_fd_sc_hs__o2bb2ai_1_1/a_397_74#
+ sky130_fd_sc_hs__o2bb2ai_1_1/a_131_383# sky130_fd_sc_hs__o2bb2ai_1
Xsky130_fd_sc_hs__nor2b_1_3 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__fa_2_3/SUM sky130_fd_sc_hs__nor2b_1_3/Y
+ sky130_fd_sc_hs__or2_1_1/A sky130_fd_sc_hs__nor2b_1_3/a_278_368# sky130_fd_sc_hs__nor2b_1_3/a_27_112#
+ sky130_fd_sc_hs__nor2b_1
Xsky130_fd_sc_hs__nand2_1_5 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nor2_1_3/Y sky130_fd_sc_hs__o21a_1_5/B1
+ sky130_fd_sc_hs__o21a_1_5/A1 sky130_fd_sc_hs__nand2_1_5/a_117_74# sky130_fd_sc_hs__nand2_1
Xsky130_fd_sc_hs__nor2_1_1 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_1/Y sky130_fd_sc_hs__nor2_1_1/Y
+ sky130_fd_sc_hs__inv_4_5/Y sky130_fd_sc_hs__nor2_1_1/a_116_368# sky130_fd_sc_hs__nor2_1
Xsky130_fd_sc_hs__a21oi_1_31 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__o21a_1_7/A2 sky130_fd_sc_hs__dfrtp_4_57/D
+ sky130_fd_sc_hs__nor2_1_19/B sky130_fd_sc_hs__inv_4_29/Y sky130_fd_sc_hs__a21oi_1_31/a_117_74#
+ sky130_fd_sc_hs__a21oi_1_31/a_29_368# sky130_fd_sc_hs__a21oi_1
Xsky130_fd_sc_hs__a21oi_1_20 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nor2_1_17/Y sky130_fd_sc_hs__dfrtp_4_35/D
+ sky130_fd_sc_hs__o21a_1_9/B1 sky130_fd_sc_hs__inv_4_15/Y sky130_fd_sc_hs__a21oi_1_21/a_117_74#
+ sky130_fd_sc_hs__a21oi_1_21/a_29_368# sky130_fd_sc_hs__a21oi_1
Xsky130_fd_sc_hs__a21oi_1_64 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nor2_1_63/Y sky130_fd_sc_hs__dfrbp_1_17/D
+ sky130_fd_sc_hs__nor2_1_63/B sky130_fd_sc_hs__inv_4_71/Y sky130_fd_sc_hs__a21oi_1_65/a_117_74#
+ sky130_fd_sc_hs__a21oi_1_65/a_29_368# sky130_fd_sc_hs__a21oi_1
Xsky130_fd_sc_hs__a21oi_1_53 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nor2_1_35/Y sky130_fd_sc_hs__dfrtp_4_85/D
+ sky130_fd_sc_hs__nor2_1_35/B sky130_fd_sc_hs__inv_4_47/Y sky130_fd_sc_hs__a21oi_1_53/a_117_74#
+ sky130_fd_sc_hs__a21oi_1_53/a_29_368# sky130_fd_sc_hs__a21oi_1
Xsky130_fd_sc_hs__a21oi_1_42 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nor2_1_25/Y sky130_fd_sc_hs__dfrtp_4_79/D
+ sky130_fd_sc_hs__nor2_1_25/B sky130_fd_sc_hs__inv_4_41/Y sky130_fd_sc_hs__a21oi_1_43/a_117_74#
+ sky130_fd_sc_hs__a21oi_1_43/a_29_368# sky130_fd_sc_hs__a21oi_1
Xsky130_fd_sc_hs__a21oi_1_97 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__a22o_1_29/X sky130_fd_sc_hs__a21oi_1_97/Y
+ sky130_fd_sc_hs__or2_1_3/B sky130_fd_sc_hs__or2_1_3/A sky130_fd_sc_hs__a21oi_1_97/a_117_74#
+ sky130_fd_sc_hs__a21oi_1_97/a_29_368# sky130_fd_sc_hs__a21oi_1
Xsky130_fd_sc_hs__a21oi_1_86 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nor3_1_1/C sky130_fd_sc_hs__maj3_1_1/B
+ sky130_fd_sc_hs__o31ai_1_5/Y sky130_fd_sc_hs__nand2_1_67/Y sky130_fd_sc_hs__a21oi_1_87/a_117_74#
+ sky130_fd_sc_hs__a21oi_1_87/a_29_368# sky130_fd_sc_hs__a21oi_1
Xsky130_fd_sc_hs__a21oi_1_75 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__o22ai_1_9/Y sky130_fd_sc_hs__a31oi_1_1/A2
+ sky130_fd_sc_hs__inv_4_77/Y sky130_fd_sc_hs__a31oi_2_1/Y sky130_fd_sc_hs__a21oi_1_75/a_117_74#
+ sky130_fd_sc_hs__a21oi_1_75/a_29_368# sky130_fd_sc_hs__a21oi_1
Xsky130_fd_sc_hs__xor2_1_9 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__xor2_1_9/A sky130_fd_sc_hs__fa_2_9/B
+ sky130_fd_sc_hs__xor2_1_9/X sky130_fd_sc_hs__xor2_1_9/a_194_125# sky130_fd_sc_hs__xor2_1_9/a_355_368#
+ sky130_fd_sc_hs__xor2_1_9/a_455_87# sky130_fd_sc_hs__xor2_1_9/a_158_392# sky130_fd_sc_hs__xor2_1
Xsky130_fd_sc_hs__nand2b_1_7 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__xnor2_1_7/B sky130_fd_sc_hs__nor3_1_7/Y
+ sky130_fd_sc_hs__nor2_1_89/A sky130_fd_sc_hs__nand2b_1_7/a_269_74# sky130_fd_sc_hs__nand2b_1_7/a_27_112#
+ sky130_fd_sc_hs__nand2b_1
Xsky130_fd_sc_hs__dfrbp_1_9 DVSS DVDD sky130_fd_sc_hs__clkbuf_8_1/X DVDD DVSS sky130_fd_sc_hs__inv_4_69/A
+ sky130_fd_sc_hs__clkbuf_2_1/X sky130_fd_sc_hs__o21a_1_45/X sky130_fd_sc_hs__dfrbp_1_9/Q_N
+ sky130_fd_sc_hs__dfrbp_1_9/a_498_360# sky130_fd_sc_hs__dfrbp_1_9/a_1224_74# sky130_fd_sc_hs__dfrbp_1_9/a_2026_424#
+ sky130_fd_sc_hs__dfrbp_1_9/a_1482_48# sky130_fd_sc_hs__dfrbp_1_9/a_125_78# sky130_fd_sc_hs__dfrbp_1_9/a_796_463#
+ sky130_fd_sc_hs__dfrbp_1_9/a_910_118# sky130_fd_sc_hs__dfrbp_1_9/a_1465_471# sky130_fd_sc_hs__dfrbp_1_9/a_832_118#
+ sky130_fd_sc_hs__dfrbp_1_9/a_841_401# sky130_fd_sc_hs__dfrbp_1_9/a_38_78# sky130_fd_sc_hs__dfrbp_1_9/a_1434_74#
+ sky130_fd_sc_hs__dfrbp_1_9/a_706_463# sky130_fd_sc_hs__dfrbp_1_9/a_319_360# sky130_fd_sc_hs__dfrbp_1_9/a_1624_74#
+ sky130_fd_sc_hs__dfrbp_1
Xsky130_fd_sc_hs__a32oi_1_6 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__o21ai_1_3/Y fine_control_avg_window_select[0]
+ sky130_fd_sc_hs__a32oi_1_7/B1 sky130_fd_sc_hs__inv_4_33/Y sky130_fd_sc_hs__a32oi_1_7/Y
+ sky130_fd_sc_hs__a32oi_1_7/A1 sky130_fd_sc_hs__a32oi_1_7/a_391_74# sky130_fd_sc_hs__a32oi_1_7/a_27_368#
+ sky130_fd_sc_hs__a32oi_1_7/a_119_74# sky130_fd_sc_hs__a32oi_1_7/a_469_74# sky130_fd_sc_hs__a32oi_1
Xsky130_fd_sc_hs__o21a_1_2 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__o21a_1_3/X sky130_fd_sc_hs__nor2_1_1/Y
+ sky130_fd_sc_hs__nor2_1_3/B sky130_fd_sc_hs__o21a_1_3/A1 sky130_fd_sc_hs__o21a_1_3/a_320_74#
+ sky130_fd_sc_hs__o21a_1_3/a_376_387# sky130_fd_sc_hs__o21a_1_3/a_83_244# sky130_fd_sc_hs__o21a_1
Xsky130_fd_sc_hs__fa_2_21 DVSS DVDD sky130_fd_sc_hs__fa_2_9/B DVDD DVSS sky130_fd_sc_hs__fa_2_21/CIN
+ sky130_fd_sc_hs__fa_2_21/B sky130_fd_sc_hs__fa_2_23/CIN sky130_fd_sc_hs__fa_2_21/SUM
+ sky130_fd_sc_hs__fa_2_21/a_27_378# sky130_fd_sc_hs__fa_2_21/a_701_79# sky130_fd_sc_hs__fa_2_21/a_484_347#
+ sky130_fd_sc_hs__fa_2_21/a_1094_347# sky130_fd_sc_hs__fa_2_21/a_1205_79# sky130_fd_sc_hs__fa_2_21/a_27_79#
+ sky130_fd_sc_hs__fa_2_21/a_1202_368# sky130_fd_sc_hs__fa_2_21/a_336_347# sky130_fd_sc_hs__fa_2_21/a_992_347#
+ sky130_fd_sc_hs__fa_2_21/a_1119_79# sky130_fd_sc_hs__fa_2_21/a_487_79# sky130_fd_sc_hs__fa_2_21/a_683_347#
+ sky130_fd_sc_hs__fa_2
Xsky130_fd_sc_hs__fa_2_10 DVSS DVDD sky130_fd_sc_hs__fa_2_9/B DVDD DVSS sky130_fd_sc_hs__fa_2_7/COUT
+ sky130_fd_sc_hs__fa_2_11/B sky130_fd_sc_hs__fa_2_13/CIN sky130_fd_sc_hs__fa_2_11/SUM
+ sky130_fd_sc_hs__fa_2_11/a_27_378# sky130_fd_sc_hs__fa_2_11/a_701_79# sky130_fd_sc_hs__fa_2_11/a_484_347#
+ sky130_fd_sc_hs__fa_2_11/a_1094_347# sky130_fd_sc_hs__fa_2_11/a_1205_79# sky130_fd_sc_hs__fa_2_11/a_27_79#
+ sky130_fd_sc_hs__fa_2_11/a_1202_368# sky130_fd_sc_hs__fa_2_11/a_336_347# sky130_fd_sc_hs__fa_2_11/a_992_347#
+ sky130_fd_sc_hs__fa_2_11/a_1119_79# sky130_fd_sc_hs__fa_2_11/a_487_79# sky130_fd_sc_hs__fa_2_11/a_683_347#
+ sky130_fd_sc_hs__fa_2
Xsky130_fd_sc_hs__dfrtn_1_7 DVSS DVDD sky130_fd_sc_hs__clkbuf_8_1/X DVDD DVSS sky130_fd_sc_hs__clkbuf_2_1/X
+ sky130_fd_sc_hs__inv_4_53/A sky130_fd_sc_hs__dfrtn_1_7/D sky130_fd_sc_hs__dfrtn_1_7/a_1266_119#
+ sky130_fd_sc_hs__dfrtn_1_7/a_1736_119# sky130_fd_sc_hs__dfrtn_1_7/a_817_508# sky130_fd_sc_hs__dfrtn_1_7/a_120_74#
+ sky130_fd_sc_hs__dfrtn_1_7/a_1547_508# sky130_fd_sc_hs__dfrtn_1_7/a_922_127# sky130_fd_sc_hs__dfrtn_1_7/a_33_74#
+ sky130_fd_sc_hs__dfrtn_1_7/a_714_127# sky130_fd_sc_hs__dfrtn_1_7/a_1934_94# sky130_fd_sc_hs__dfrtn_1_7/a_1550_119#
+ sky130_fd_sc_hs__dfrtn_1_7/a_1598_93# sky130_fd_sc_hs__dfrtn_1_7/a_300_74# sky130_fd_sc_hs__dfrtn_1_7/a_507_368#
+ sky130_fd_sc_hs__dfrtn_1_7/a_856_304# sky130_fd_sc_hs__dfrtn_1_7/a_850_127# sky130_fd_sc_hs__dfrtn_1
Xsky130_fd_sc_hs__o211ai_1_7 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__a21oi_1_97/Y sky130_fd_sc_hs__nor3_1_3/A
+ sky130_fd_sc_hs__nor2_1_61/Y sky130_fd_sc_hs__maj3_1_3/B sky130_fd_sc_hs__maj3_1_3/A
+ sky130_fd_sc_hs__o211ai_1_7/a_31_74# sky130_fd_sc_hs__o211ai_1_7/a_311_74# sky130_fd_sc_hs__o211ai_1_7/a_116_368#
+ sky130_fd_sc_hs__o211ai_1
Xsky130_fd_sc_hs__o21a_1_50 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__o21a_1_51/X sky130_fd_sc_hs__nor2_1_83/Y
+ sky130_fd_sc_hs__o21a_1_51/B1 sky130_fd_sc_hs__maj3_1_1/A sky130_fd_sc_hs__o21a_1_51/a_320_74#
+ sky130_fd_sc_hs__o21a_1_51/a_376_387# sky130_fd_sc_hs__o21a_1_51/a_83_244# sky130_fd_sc_hs__o21a_1
Xsky130_fd_sc_hs__o21a_1_61 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__o21a_1_61/X sky130_fd_sc_hs__o21a_1_61/A2
+ sky130_fd_sc_hs__xnor2_1_5/B sky130_fd_sc_hs__maj3_1_3/A sky130_fd_sc_hs__o21a_1_61/a_320_74#
+ sky130_fd_sc_hs__o21a_1_61/a_376_387# sky130_fd_sc_hs__o21a_1_61/a_83_244# sky130_fd_sc_hs__o21a_1
Xsky130_fd_sc_hs__o21a_1_72 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__o21a_1_73/X sky130_fd_sc_hs__o21a_1_73/A2
+ sky130_fd_sc_hs__o21a_1_73/B1 sky130_fd_sc_hs__or2_1_3/A sky130_fd_sc_hs__o21a_1_73/a_320_74#
+ sky130_fd_sc_hs__o21a_1_73/a_376_387# sky130_fd_sc_hs__o21a_1_73/a_83_244# sky130_fd_sc_hs__o21a_1
Xsky130_fd_sc_hs__dfrtp_4_62 DVSS DVDD sky130_fd_sc_hs__clkbuf_8_1/X DVDD DVSS sky130_fd_sc_hs__o21a_1_25/X
+ sky130_fd_sc_hs__nand2_1_47/B sky130_fd_sc_hs__o21a_1_25/A1 sky130_fd_sc_hs__dfrtp_4_63/a_37_78#
+ sky130_fd_sc_hs__dfrtp_4_63/a_494_366# sky130_fd_sc_hs__dfrtp_4_63/a_699_463# sky130_fd_sc_hs__dfrtp_4_63/a_313_74#
+ sky130_fd_sc_hs__dfrtp_4_63/a_1627_493# sky130_fd_sc_hs__dfrtp_4_63/a_1678_395#
+ sky130_fd_sc_hs__dfrtp_4_63/a_1827_81# sky130_fd_sc_hs__dfrtp_4_63/a_789_463# sky130_fd_sc_hs__dfrtp_4_63/a_1350_392#
+ sky130_fd_sc_hs__dfrtp_4_63/a_834_355# sky130_fd_sc_hs__dfrtp_4_63/a_812_138# sky130_fd_sc_hs__dfrtp_4_63/a_124_78#
+ sky130_fd_sc_hs__dfrtp_4_63/a_1647_81# sky130_fd_sc_hs__dfrtp_4_63/a_2010_409# sky130_fd_sc_hs__dfrtp_4_63/a_890_138#
+ sky130_fd_sc_hs__dfrtp_4
Xsky130_fd_sc_hs__dfrtp_4_51 DVSS DVDD sky130_fd_sc_hs__clkbuf_8_1/X DVDD DVSS sky130_fd_sc_hs__o21a_1_13/X
+ sky130_fd_sc_hs__nand2_1_47/B sky130_fd_sc_hs__o21a_1_13/A1 sky130_fd_sc_hs__dfrtp_4_51/a_37_78#
+ sky130_fd_sc_hs__dfrtp_4_51/a_494_366# sky130_fd_sc_hs__dfrtp_4_51/a_699_463# sky130_fd_sc_hs__dfrtp_4_51/a_313_74#
+ sky130_fd_sc_hs__dfrtp_4_51/a_1627_493# sky130_fd_sc_hs__dfrtp_4_51/a_1678_395#
+ sky130_fd_sc_hs__dfrtp_4_51/a_1827_81# sky130_fd_sc_hs__dfrtp_4_51/a_789_463# sky130_fd_sc_hs__dfrtp_4_51/a_1350_392#
+ sky130_fd_sc_hs__dfrtp_4_51/a_834_355# sky130_fd_sc_hs__dfrtp_4_51/a_812_138# sky130_fd_sc_hs__dfrtp_4_51/a_124_78#
+ sky130_fd_sc_hs__dfrtp_4_51/a_1647_81# sky130_fd_sc_hs__dfrtp_4_51/a_2010_409# sky130_fd_sc_hs__dfrtp_4_51/a_890_138#
+ sky130_fd_sc_hs__dfrtp_4
Xsky130_fd_sc_hs__dfrtp_4_40 DVSS DVDD sky130_fd_sc_hs__clkbuf_8_1/X DVDD DVSS sky130_fd_sc_hs__o21a_1_17/X
+ sky130_fd_sc_hs__nand2_1_47/B sky130_fd_sc_hs__o21a_1_17/A1 sky130_fd_sc_hs__dfrtp_4_41/a_37_78#
+ sky130_fd_sc_hs__dfrtp_4_41/a_494_366# sky130_fd_sc_hs__dfrtp_4_41/a_699_463# sky130_fd_sc_hs__dfrtp_4_41/a_313_74#
+ sky130_fd_sc_hs__dfrtp_4_41/a_1627_493# sky130_fd_sc_hs__dfrtp_4_41/a_1678_395#
+ sky130_fd_sc_hs__dfrtp_4_41/a_1827_81# sky130_fd_sc_hs__dfrtp_4_41/a_789_463# sky130_fd_sc_hs__dfrtp_4_41/a_1350_392#
+ sky130_fd_sc_hs__dfrtp_4_41/a_834_355# sky130_fd_sc_hs__dfrtp_4_41/a_812_138# sky130_fd_sc_hs__dfrtp_4_41/a_124_78#
+ sky130_fd_sc_hs__dfrtp_4_41/a_1647_81# sky130_fd_sc_hs__dfrtp_4_41/a_2010_409# sky130_fd_sc_hs__dfrtp_4_41/a_890_138#
+ sky130_fd_sc_hs__dfrtp_4
Xsky130_fd_sc_hs__dfrtp_4_84 DVSS DVDD sky130_fd_sc_hs__clkbuf_8_1/X DVDD DVSS sky130_fd_sc_hs__dfrtp_4_85/D
+ sky130_fd_sc_hs__nand2_1_47/B sky130_fd_sc_hs__inv_4_47/A sky130_fd_sc_hs__dfrtp_4_85/a_37_78#
+ sky130_fd_sc_hs__dfrtp_4_85/a_494_366# sky130_fd_sc_hs__dfrtp_4_85/a_699_463# sky130_fd_sc_hs__dfrtp_4_85/a_313_74#
+ sky130_fd_sc_hs__dfrtp_4_85/a_1627_493# sky130_fd_sc_hs__dfrtp_4_85/a_1678_395#
+ sky130_fd_sc_hs__dfrtp_4_85/a_1827_81# sky130_fd_sc_hs__dfrtp_4_85/a_789_463# sky130_fd_sc_hs__dfrtp_4_85/a_1350_392#
+ sky130_fd_sc_hs__dfrtp_4_85/a_834_355# sky130_fd_sc_hs__dfrtp_4_85/a_812_138# sky130_fd_sc_hs__dfrtp_4_85/a_124_78#
+ sky130_fd_sc_hs__dfrtp_4_85/a_1647_81# sky130_fd_sc_hs__dfrtp_4_85/a_2010_409# sky130_fd_sc_hs__dfrtp_4_85/a_890_138#
+ sky130_fd_sc_hs__dfrtp_4
Xsky130_fd_sc_hs__dfrtp_4_73 DVSS DVDD sky130_fd_sc_hs__inv_4_49/Y DVDD DVSS sky130_fd_sc_hs__nor2b_1_21/Y
+ sky130_fd_sc_hs__dfstp_2_1/CLK sky130_fd_sc_hs__fa_2_23/B sky130_fd_sc_hs__dfrtp_4_73/a_37_78#
+ sky130_fd_sc_hs__dfrtp_4_73/a_494_366# sky130_fd_sc_hs__dfrtp_4_73/a_699_463# sky130_fd_sc_hs__dfrtp_4_73/a_313_74#
+ sky130_fd_sc_hs__dfrtp_4_73/a_1627_493# sky130_fd_sc_hs__dfrtp_4_73/a_1678_395#
+ sky130_fd_sc_hs__dfrtp_4_73/a_1827_81# sky130_fd_sc_hs__dfrtp_4_73/a_789_463# sky130_fd_sc_hs__dfrtp_4_73/a_1350_392#
+ sky130_fd_sc_hs__dfrtp_4_73/a_834_355# sky130_fd_sc_hs__dfrtp_4_73/a_812_138# sky130_fd_sc_hs__dfrtp_4_73/a_124_78#
+ sky130_fd_sc_hs__dfrtp_4_73/a_1647_81# sky130_fd_sc_hs__dfrtp_4_73/a_2010_409# sky130_fd_sc_hs__dfrtp_4_73/a_890_138#
+ sky130_fd_sc_hs__dfrtp_4
Xsky130_fd_sc_hs__a22o_1_6 DVSS DVDD DVDD DVSS osc_fine_con_final[12] manual_control_osc[12]
+ sky130_fd_sc_hs__inv_4_43/Y sky130_fd_sc_hs__xor2_1_9/A fftl_en sky130_fd_sc_hs__a22o_1_7/a_222_392#
+ sky130_fd_sc_hs__a22o_1_7/a_230_79# sky130_fd_sc_hs__a22o_1_7/a_52_123# sky130_fd_sc_hs__a22o_1_7/a_132_392#
+ sky130_fd_sc_hs__a22o_1
Xsky130_fd_sc_hs__fa_2_9 DVSS DVDD sky130_fd_sc_hs__fa_2_9/A DVDD DVSS sky130_fd_sc_hs__xor2_1_1/X
+ sky130_fd_sc_hs__fa_2_9/B sky130_fd_sc_hs__fa_2_5/CIN sky130_fd_sc_hs__fa_2_9/SUM
+ sky130_fd_sc_hs__fa_2_9/a_27_378# sky130_fd_sc_hs__fa_2_9/a_701_79# sky130_fd_sc_hs__fa_2_9/a_484_347#
+ sky130_fd_sc_hs__fa_2_9/a_1094_347# sky130_fd_sc_hs__fa_2_9/a_1205_79# sky130_fd_sc_hs__fa_2_9/a_27_79#
+ sky130_fd_sc_hs__fa_2_9/a_1202_368# sky130_fd_sc_hs__fa_2_9/a_336_347# sky130_fd_sc_hs__fa_2_9/a_992_347#
+ sky130_fd_sc_hs__fa_2_9/a_1119_79# sky130_fd_sc_hs__fa_2_9/a_487_79# sky130_fd_sc_hs__fa_2_9/a_683_347#
+ sky130_fd_sc_hs__fa_2
Xsky130_fd_sc_hs__o2bb2ai_1_1 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nor4_1_3/B sky130_fd_sc_hs__inv_4_73/Y
+ sky130_fd_sc_hs__inv_4_83/Y sky130_fd_sc_hs__nor2_1_65/A sky130_fd_sc_hs__dfrbp_1_7/Q
+ sky130_fd_sc_hs__o2bb2ai_1_1/a_114_74# sky130_fd_sc_hs__o2bb2ai_1_1/a_490_368# sky130_fd_sc_hs__o2bb2ai_1_1/a_397_74#
+ sky130_fd_sc_hs__o2bb2ai_1_1/a_131_383# sky130_fd_sc_hs__o2bb2ai_1
Xsky130_fd_sc_hs__nor2b_1_4 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__fa_2_5/SUM sky130_fd_sc_hs__nor2b_1_5/Y
+ sky130_fd_sc_hs__or2_1_1/A sky130_fd_sc_hs__nor2b_1_5/a_278_368# sky130_fd_sc_hs__nor2b_1_5/a_27_112#
+ sky130_fd_sc_hs__nor2b_1
Xsky130_fd_sc_hs__nand2_1_6 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nor2_1_9/Y sky130_fd_sc_hs__o21a_1_9/B1
+ sky130_fd_sc_hs__o21a_1_9/A1 sky130_fd_sc_hs__nand2_1_7/a_117_74# sky130_fd_sc_hs__nand2_1
Xsky130_fd_sc_hs__nor2_1_2 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nor2_1_3/B sky130_fd_sc_hs__nor2_1_3/Y
+ sky130_fd_sc_hs__inv_4_3/Y sky130_fd_sc_hs__nor2_1_3/a_116_368# sky130_fd_sc_hs__nor2_1
Xsky130_fd_sc_hs__a21oi_1_21 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nor2_1_17/Y sky130_fd_sc_hs__dfrtp_4_35/D
+ sky130_fd_sc_hs__o21a_1_9/B1 sky130_fd_sc_hs__inv_4_15/Y sky130_fd_sc_hs__a21oi_1_21/a_117_74#
+ sky130_fd_sc_hs__a21oi_1_21/a_29_368# sky130_fd_sc_hs__a21oi_1
Xsky130_fd_sc_hs__a21oi_1_10 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nor2_1_11/Y sky130_fd_sc_hs__dfrtp_4_25/D
+ sky130_fd_sc_hs__o21a_1_5/B1 sky130_fd_sc_hs__inv_4_13/Y sky130_fd_sc_hs__a21oi_1_11/a_117_74#
+ sky130_fd_sc_hs__a21oi_1_11/a_29_368# sky130_fd_sc_hs__a21oi_1
Xsky130_fd_sc_hs__a21oi_1_65 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nor2_1_63/Y sky130_fd_sc_hs__dfrbp_1_17/D
+ sky130_fd_sc_hs__nor2_1_63/B sky130_fd_sc_hs__inv_4_71/Y sky130_fd_sc_hs__a21oi_1_65/a_117_74#
+ sky130_fd_sc_hs__a21oi_1_65/a_29_368# sky130_fd_sc_hs__a21oi_1
Xsky130_fd_sc_hs__a21oi_1_54 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nor2_1_49/Y sky130_fd_sc_hs__dfrtn_1_13/D
+ sky130_fd_sc_hs__nor2_1_49/B sky130_fd_sc_hs__inv_4_59/Y sky130_fd_sc_hs__a21oi_1_55/a_117_74#
+ sky130_fd_sc_hs__a21oi_1_55/a_29_368# sky130_fd_sc_hs__a21oi_1
Xsky130_fd_sc_hs__a21oi_1_43 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nor2_1_25/Y sky130_fd_sc_hs__dfrtp_4_79/D
+ sky130_fd_sc_hs__nor2_1_25/B sky130_fd_sc_hs__inv_4_41/Y sky130_fd_sc_hs__a21oi_1_43/a_117_74#
+ sky130_fd_sc_hs__a21oi_1_43/a_29_368# sky130_fd_sc_hs__a21oi_1
Xsky130_fd_sc_hs__a21oi_1_32 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nor2_1_21/Y sky130_fd_sc_hs__dfrtp_4_59/D
+ sky130_fd_sc_hs__nor2_1_21/B sky130_fd_sc_hs__inv_4_31/Y sky130_fd_sc_hs__a21oi_1_33/a_117_74#
+ sky130_fd_sc_hs__a21oi_1_33/a_29_368# sky130_fd_sc_hs__a21oi_1
Xsky130_fd_sc_hs__a21oi_1_98 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nor3_1_9/C sky130_fd_sc_hs__o22ai_1_9/A1
+ sky130_fd_sc_hs__o211ai_1_9/C1 sky130_fd_sc_hs__nor3_1_9/B sky130_fd_sc_hs__a21oi_1_99/a_117_74#
+ sky130_fd_sc_hs__a21oi_1_99/a_29_368# sky130_fd_sc_hs__a21oi_1
Xsky130_fd_sc_hs__a21oi_1_87 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nor3_1_1/C sky130_fd_sc_hs__maj3_1_1/B
+ sky130_fd_sc_hs__o31ai_1_5/Y sky130_fd_sc_hs__nand2_1_67/Y sky130_fd_sc_hs__a21oi_1_87/a_117_74#
+ sky130_fd_sc_hs__a21oi_1_87/a_29_368# sky130_fd_sc_hs__a21oi_1
Xsky130_fd_sc_hs__a21oi_1_76 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nor4_1_1/D sky130_fd_sc_hs__a31oi_2_1/A1
+ sky130_fd_sc_hs__nand2_1_59/Y sky130_fd_sc_hs__nor4_1_1/C sky130_fd_sc_hs__a21oi_1_77/a_117_74#
+ sky130_fd_sc_hs__a21oi_1_77/a_29_368# sky130_fd_sc_hs__a21oi_1
Xsky130_fd_sc_hs__nand2b_1_8 DVSS DVDD DVDD DVSS rst sky130_fd_sc_hs__nor2_1_81/Y
+ sky130_fd_sc_hs__nor2b_1_41/A sky130_fd_sc_hs__nand2b_1_9/a_269_74# sky130_fd_sc_hs__nand2b_1_9/a_27_112#
+ sky130_fd_sc_hs__nand2b_1
Xsky130_fd_sc_hs__a32oi_1_7 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__o21ai_1_3/Y fine_control_avg_window_select[0]
+ sky130_fd_sc_hs__a32oi_1_7/B1 sky130_fd_sc_hs__inv_4_33/Y sky130_fd_sc_hs__a32oi_1_7/Y
+ sky130_fd_sc_hs__a32oi_1_7/A1 sky130_fd_sc_hs__a32oi_1_7/a_391_74# sky130_fd_sc_hs__a32oi_1_7/a_27_368#
+ sky130_fd_sc_hs__a32oi_1_7/a_119_74# sky130_fd_sc_hs__a32oi_1_7/a_469_74# sky130_fd_sc_hs__a32oi_1
Xsky130_fd_sc_hs__o21a_1_3 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__o21a_1_3/X sky130_fd_sc_hs__nor2_1_1/Y
+ sky130_fd_sc_hs__nor2_1_3/B sky130_fd_sc_hs__o21a_1_3/A1 sky130_fd_sc_hs__o21a_1_3/a_320_74#
+ sky130_fd_sc_hs__o21a_1_3/a_376_387# sky130_fd_sc_hs__o21a_1_3/a_83_244# sky130_fd_sc_hs__o21a_1
Xsky130_fd_sc_hs__fa_2_22 DVSS DVDD sky130_fd_sc_hs__fa_2_9/B DVDD DVSS sky130_fd_sc_hs__fa_2_23/CIN
+ sky130_fd_sc_hs__fa_2_23/B sky130_fd_sc_hs__fa_2_15/CIN sky130_fd_sc_hs__fa_2_23/SUM
+ sky130_fd_sc_hs__fa_2_23/a_27_378# sky130_fd_sc_hs__fa_2_23/a_701_79# sky130_fd_sc_hs__fa_2_23/a_484_347#
+ sky130_fd_sc_hs__fa_2_23/a_1094_347# sky130_fd_sc_hs__fa_2_23/a_1205_79# sky130_fd_sc_hs__fa_2_23/a_27_79#
+ sky130_fd_sc_hs__fa_2_23/a_1202_368# sky130_fd_sc_hs__fa_2_23/a_336_347# sky130_fd_sc_hs__fa_2_23/a_992_347#
+ sky130_fd_sc_hs__fa_2_23/a_1119_79# sky130_fd_sc_hs__fa_2_23/a_487_79# sky130_fd_sc_hs__fa_2_23/a_683_347#
+ sky130_fd_sc_hs__fa_2
Xsky130_fd_sc_hs__fa_2_11 DVSS DVDD sky130_fd_sc_hs__fa_2_9/B DVDD DVSS sky130_fd_sc_hs__fa_2_7/COUT
+ sky130_fd_sc_hs__fa_2_11/B sky130_fd_sc_hs__fa_2_13/CIN sky130_fd_sc_hs__fa_2_11/SUM
+ sky130_fd_sc_hs__fa_2_11/a_27_378# sky130_fd_sc_hs__fa_2_11/a_701_79# sky130_fd_sc_hs__fa_2_11/a_484_347#
+ sky130_fd_sc_hs__fa_2_11/a_1094_347# sky130_fd_sc_hs__fa_2_11/a_1205_79# sky130_fd_sc_hs__fa_2_11/a_27_79#
+ sky130_fd_sc_hs__fa_2_11/a_1202_368# sky130_fd_sc_hs__fa_2_11/a_336_347# sky130_fd_sc_hs__fa_2_11/a_992_347#
+ sky130_fd_sc_hs__fa_2_11/a_1119_79# sky130_fd_sc_hs__fa_2_11/a_487_79# sky130_fd_sc_hs__fa_2_11/a_683_347#
+ sky130_fd_sc_hs__fa_2
Xsky130_fd_sc_hs__dfrtn_1_8 DVSS DVDD sky130_fd_sc_hs__clkbuf_8_1/X DVDD DVSS sky130_fd_sc_hs__clkbuf_2_1/X
+ sky130_fd_sc_hs__nor2_1_65/A sky130_fd_sc_hs__o21a_1_37/X sky130_fd_sc_hs__dfrtn_1_9/a_1266_119#
+ sky130_fd_sc_hs__dfrtn_1_9/a_1736_119# sky130_fd_sc_hs__dfrtn_1_9/a_817_508# sky130_fd_sc_hs__dfrtn_1_9/a_120_74#
+ sky130_fd_sc_hs__dfrtn_1_9/a_1547_508# sky130_fd_sc_hs__dfrtn_1_9/a_922_127# sky130_fd_sc_hs__dfrtn_1_9/a_33_74#
+ sky130_fd_sc_hs__dfrtn_1_9/a_714_127# sky130_fd_sc_hs__dfrtn_1_9/a_1934_94# sky130_fd_sc_hs__dfrtn_1_9/a_1550_119#
+ sky130_fd_sc_hs__dfrtn_1_9/a_1598_93# sky130_fd_sc_hs__dfrtn_1_9/a_300_74# sky130_fd_sc_hs__dfrtn_1_9/a_507_368#
+ sky130_fd_sc_hs__dfrtn_1_9/a_856_304# sky130_fd_sc_hs__dfrtn_1_9/a_850_127# sky130_fd_sc_hs__dfrtn_1
Xsky130_fd_sc_hs__o211ai_1_8 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_109/A sky130_fd_sc_hs__o22ai_1_9/B1
+ sky130_fd_sc_hs__o211ai_1_9/C1 sky130_fd_sc_hs__inv_4_107/Y sky130_fd_sc_hs__inv_4_105/A
+ sky130_fd_sc_hs__o211ai_1_9/a_31_74# sky130_fd_sc_hs__o211ai_1_9/a_311_74# sky130_fd_sc_hs__o211ai_1_9/a_116_368#
+ sky130_fd_sc_hs__o211ai_1
Xsky130_fd_sc_hs__o21a_1_51 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__o21a_1_51/X sky130_fd_sc_hs__nor2_1_83/Y
+ sky130_fd_sc_hs__o21a_1_51/B1 sky130_fd_sc_hs__maj3_1_1/A sky130_fd_sc_hs__o21a_1_51/a_320_74#
+ sky130_fd_sc_hs__o21a_1_51/a_376_387# sky130_fd_sc_hs__o21a_1_51/a_83_244# sky130_fd_sc_hs__o21a_1
Xsky130_fd_sc_hs__o21a_1_40 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__o21a_1_41/X sky130_fd_sc_hs__nor2_1_63/Y
+ sky130_fd_sc_hs__nor2_1_43/B sky130_fd_sc_hs__dfrbp_1_7/Q sky130_fd_sc_hs__o21a_1_41/a_320_74#
+ sky130_fd_sc_hs__o21a_1_41/a_376_387# sky130_fd_sc_hs__o21a_1_41/a_83_244# sky130_fd_sc_hs__o21a_1
Xsky130_fd_sc_hs__o21a_1_62 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__o21a_1_63/X sky130_fd_sc_hs__o21a_1_63/A2
+ sky130_fd_sc_hs__nor2_1_63/B sky130_fd_sc_hs__o21a_1_63/A1 sky130_fd_sc_hs__o21a_1_63/a_320_74#
+ sky130_fd_sc_hs__o21a_1_63/a_376_387# sky130_fd_sc_hs__o21a_1_63/a_83_244# sky130_fd_sc_hs__o21a_1
Xsky130_fd_sc_hs__o21a_1_73 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__o21a_1_73/X sky130_fd_sc_hs__o21a_1_73/A2
+ sky130_fd_sc_hs__o21a_1_73/B1 sky130_fd_sc_hs__or2_1_3/A sky130_fd_sc_hs__o21a_1_73/a_320_74#
+ sky130_fd_sc_hs__o21a_1_73/a_376_387# sky130_fd_sc_hs__o21a_1_73/a_83_244# sky130_fd_sc_hs__o21a_1
Xsky130_fd_sc_hs__dfrtp_4_52 DVSS DVDD sky130_fd_sc_hs__inv_4_49/Y DVDD DVSS sky130_fd_sc_hs__nor2b_1_9/Y
+ sky130_fd_sc_hs__dfstp_2_1/CLK sky130_fd_sc_hs__fa_2_11/B sky130_fd_sc_hs__dfrtp_4_53/a_37_78#
+ sky130_fd_sc_hs__dfrtp_4_53/a_494_366# sky130_fd_sc_hs__dfrtp_4_53/a_699_463# sky130_fd_sc_hs__dfrtp_4_53/a_313_74#
+ sky130_fd_sc_hs__dfrtp_4_53/a_1627_493# sky130_fd_sc_hs__dfrtp_4_53/a_1678_395#
+ sky130_fd_sc_hs__dfrtp_4_53/a_1827_81# sky130_fd_sc_hs__dfrtp_4_53/a_789_463# sky130_fd_sc_hs__dfrtp_4_53/a_1350_392#
+ sky130_fd_sc_hs__dfrtp_4_53/a_834_355# sky130_fd_sc_hs__dfrtp_4_53/a_812_138# sky130_fd_sc_hs__dfrtp_4_53/a_124_78#
+ sky130_fd_sc_hs__dfrtp_4_53/a_1647_81# sky130_fd_sc_hs__dfrtp_4_53/a_2010_409# sky130_fd_sc_hs__dfrtp_4_53/a_890_138#
+ sky130_fd_sc_hs__dfrtp_4
Xsky130_fd_sc_hs__dfrtp_4_41 DVSS DVDD sky130_fd_sc_hs__clkbuf_8_1/X DVDD DVSS sky130_fd_sc_hs__o21a_1_17/X
+ sky130_fd_sc_hs__nand2_1_47/B sky130_fd_sc_hs__o21a_1_17/A1 sky130_fd_sc_hs__dfrtp_4_41/a_37_78#
+ sky130_fd_sc_hs__dfrtp_4_41/a_494_366# sky130_fd_sc_hs__dfrtp_4_41/a_699_463# sky130_fd_sc_hs__dfrtp_4_41/a_313_74#
+ sky130_fd_sc_hs__dfrtp_4_41/a_1627_493# sky130_fd_sc_hs__dfrtp_4_41/a_1678_395#
+ sky130_fd_sc_hs__dfrtp_4_41/a_1827_81# sky130_fd_sc_hs__dfrtp_4_41/a_789_463# sky130_fd_sc_hs__dfrtp_4_41/a_1350_392#
+ sky130_fd_sc_hs__dfrtp_4_41/a_834_355# sky130_fd_sc_hs__dfrtp_4_41/a_812_138# sky130_fd_sc_hs__dfrtp_4_41/a_124_78#
+ sky130_fd_sc_hs__dfrtp_4_41/a_1647_81# sky130_fd_sc_hs__dfrtp_4_41/a_2010_409# sky130_fd_sc_hs__dfrtp_4_41/a_890_138#
+ sky130_fd_sc_hs__dfrtp_4
Xsky130_fd_sc_hs__dfrtp_4_30 DVSS DVDD sky130_fd_sc_hs__clkbuf_8_1/X DVDD DVSS sky130_fd_sc_hs__dfrtp_4_31/D
+ sky130_fd_sc_hs__nand2_1_47/B sky130_fd_sc_hs__inv_4_19/A sky130_fd_sc_hs__dfrtp_4_31/a_37_78#
+ sky130_fd_sc_hs__dfrtp_4_31/a_494_366# sky130_fd_sc_hs__dfrtp_4_31/a_699_463# sky130_fd_sc_hs__dfrtp_4_31/a_313_74#
+ sky130_fd_sc_hs__dfrtp_4_31/a_1627_493# sky130_fd_sc_hs__dfrtp_4_31/a_1678_395#
+ sky130_fd_sc_hs__dfrtp_4_31/a_1827_81# sky130_fd_sc_hs__dfrtp_4_31/a_789_463# sky130_fd_sc_hs__dfrtp_4_31/a_1350_392#
+ sky130_fd_sc_hs__dfrtp_4_31/a_834_355# sky130_fd_sc_hs__dfrtp_4_31/a_812_138# sky130_fd_sc_hs__dfrtp_4_31/a_124_78#
+ sky130_fd_sc_hs__dfrtp_4_31/a_1647_81# sky130_fd_sc_hs__dfrtp_4_31/a_2010_409# sky130_fd_sc_hs__dfrtp_4_31/a_890_138#
+ sky130_fd_sc_hs__dfrtp_4
Xsky130_fd_sc_hs__dfrtp_4_85 DVSS DVDD sky130_fd_sc_hs__clkbuf_8_1/X DVDD DVSS sky130_fd_sc_hs__dfrtp_4_85/D
+ sky130_fd_sc_hs__nand2_1_47/B sky130_fd_sc_hs__inv_4_47/A sky130_fd_sc_hs__dfrtp_4_85/a_37_78#
+ sky130_fd_sc_hs__dfrtp_4_85/a_494_366# sky130_fd_sc_hs__dfrtp_4_85/a_699_463# sky130_fd_sc_hs__dfrtp_4_85/a_313_74#
+ sky130_fd_sc_hs__dfrtp_4_85/a_1627_493# sky130_fd_sc_hs__dfrtp_4_85/a_1678_395#
+ sky130_fd_sc_hs__dfrtp_4_85/a_1827_81# sky130_fd_sc_hs__dfrtp_4_85/a_789_463# sky130_fd_sc_hs__dfrtp_4_85/a_1350_392#
+ sky130_fd_sc_hs__dfrtp_4_85/a_834_355# sky130_fd_sc_hs__dfrtp_4_85/a_812_138# sky130_fd_sc_hs__dfrtp_4_85/a_124_78#
+ sky130_fd_sc_hs__dfrtp_4_85/a_1647_81# sky130_fd_sc_hs__dfrtp_4_85/a_2010_409# sky130_fd_sc_hs__dfrtp_4_85/a_890_138#
+ sky130_fd_sc_hs__dfrtp_4
Xsky130_fd_sc_hs__dfrtp_4_74 DVSS DVDD sky130_fd_sc_hs__inv_4_49/Y DVDD DVSS sky130_fd_sc_hs__nor2b_1_17/Y
+ sky130_fd_sc_hs__dfstp_2_1/CLK sky130_fd_sc_hs__fa_2_17/B sky130_fd_sc_hs__dfrtp_4_75/a_37_78#
+ sky130_fd_sc_hs__dfrtp_4_75/a_494_366# sky130_fd_sc_hs__dfrtp_4_75/a_699_463# sky130_fd_sc_hs__dfrtp_4_75/a_313_74#
+ sky130_fd_sc_hs__dfrtp_4_75/a_1627_493# sky130_fd_sc_hs__dfrtp_4_75/a_1678_395#
+ sky130_fd_sc_hs__dfrtp_4_75/a_1827_81# sky130_fd_sc_hs__dfrtp_4_75/a_789_463# sky130_fd_sc_hs__dfrtp_4_75/a_1350_392#
+ sky130_fd_sc_hs__dfrtp_4_75/a_834_355# sky130_fd_sc_hs__dfrtp_4_75/a_812_138# sky130_fd_sc_hs__dfrtp_4_75/a_124_78#
+ sky130_fd_sc_hs__dfrtp_4_75/a_1647_81# sky130_fd_sc_hs__dfrtp_4_75/a_2010_409# sky130_fd_sc_hs__dfrtp_4_75/a_890_138#
+ sky130_fd_sc_hs__dfrtp_4
Xsky130_fd_sc_hs__dfrtp_4_63 DVSS DVDD sky130_fd_sc_hs__clkbuf_8_1/X DVDD DVSS sky130_fd_sc_hs__o21a_1_25/X
+ sky130_fd_sc_hs__nand2_1_47/B sky130_fd_sc_hs__o21a_1_25/A1 sky130_fd_sc_hs__dfrtp_4_63/a_37_78#
+ sky130_fd_sc_hs__dfrtp_4_63/a_494_366# sky130_fd_sc_hs__dfrtp_4_63/a_699_463# sky130_fd_sc_hs__dfrtp_4_63/a_313_74#
+ sky130_fd_sc_hs__dfrtp_4_63/a_1627_493# sky130_fd_sc_hs__dfrtp_4_63/a_1678_395#
+ sky130_fd_sc_hs__dfrtp_4_63/a_1827_81# sky130_fd_sc_hs__dfrtp_4_63/a_789_463# sky130_fd_sc_hs__dfrtp_4_63/a_1350_392#
+ sky130_fd_sc_hs__dfrtp_4_63/a_834_355# sky130_fd_sc_hs__dfrtp_4_63/a_812_138# sky130_fd_sc_hs__dfrtp_4_63/a_124_78#
+ sky130_fd_sc_hs__dfrtp_4_63/a_1647_81# sky130_fd_sc_hs__dfrtp_4_63/a_2010_409# sky130_fd_sc_hs__dfrtp_4_63/a_890_138#
+ sky130_fd_sc_hs__dfrtp_4
Xsky130_fd_sc_hs__a22o_1_7 DVSS DVDD DVDD DVSS osc_fine_con_final[12] manual_control_osc[12]
+ sky130_fd_sc_hs__inv_4_43/Y sky130_fd_sc_hs__xor2_1_9/A fftl_en sky130_fd_sc_hs__a22o_1_7/a_222_392#
+ sky130_fd_sc_hs__a22o_1_7/a_230_79# sky130_fd_sc_hs__a22o_1_7/a_52_123# sky130_fd_sc_hs__a22o_1_7/a_132_392#
+ sky130_fd_sc_hs__a22o_1
Xsky130_fd_sc_hs__nor2b_1_5 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__fa_2_5/SUM sky130_fd_sc_hs__nor2b_1_5/Y
+ sky130_fd_sc_hs__or2_1_1/A sky130_fd_sc_hs__nor2b_1_5/a_278_368# sky130_fd_sc_hs__nor2b_1_5/a_27_112#
+ sky130_fd_sc_hs__nor2b_1
Xsky130_fd_sc_hs__nand2_1_7 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nor2_1_9/Y sky130_fd_sc_hs__o21a_1_9/B1
+ sky130_fd_sc_hs__o21a_1_9/A1 sky130_fd_sc_hs__nand2_1_7/a_117_74# sky130_fd_sc_hs__nand2_1
Xsky130_fd_sc_hs__nor2_1_3 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nor2_1_3/B sky130_fd_sc_hs__nor2_1_3/Y
+ sky130_fd_sc_hs__inv_4_3/Y sky130_fd_sc_hs__nor2_1_3/a_116_368# sky130_fd_sc_hs__nor2_1
Xsky130_fd_sc_hs__a21oi_1_22 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nor2_1_13/Y sky130_fd_sc_hs__dfrtp_4_43/D
+ sky130_fd_sc_hs__nor2_1_13/B sky130_fd_sc_hs__inv_4_17/Y sky130_fd_sc_hs__a21oi_1_23/a_117_74#
+ sky130_fd_sc_hs__a21oi_1_23/a_29_368# sky130_fd_sc_hs__a21oi_1
Xsky130_fd_sc_hs__a21oi_1_11 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nor2_1_11/Y sky130_fd_sc_hs__dfrtp_4_25/D
+ sky130_fd_sc_hs__o21a_1_5/B1 sky130_fd_sc_hs__inv_4_13/Y sky130_fd_sc_hs__a21oi_1_11/a_117_74#
+ sky130_fd_sc_hs__a21oi_1_11/a_29_368# sky130_fd_sc_hs__a21oi_1
Xsky130_fd_sc_hs__a21oi_1_55 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nor2_1_49/Y sky130_fd_sc_hs__dfrtn_1_13/D
+ sky130_fd_sc_hs__nor2_1_49/B sky130_fd_sc_hs__inv_4_59/Y sky130_fd_sc_hs__a21oi_1_55/a_117_74#
+ sky130_fd_sc_hs__a21oi_1_55/a_29_368# sky130_fd_sc_hs__a21oi_1
Xsky130_fd_sc_hs__a21oi_1_44 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nor2_1_31/Y sky130_fd_sc_hs__dfrtp_4_83/D
+ sky130_fd_sc_hs__nor2_1_31/B sky130_fd_sc_hs__inv_4_45/Y sky130_fd_sc_hs__a21oi_1_45/a_117_74#
+ sky130_fd_sc_hs__a21oi_1_45/a_29_368# sky130_fd_sc_hs__a21oi_1
Xsky130_fd_sc_hs__a21oi_1_33 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nor2_1_21/Y sky130_fd_sc_hs__dfrtp_4_59/D
+ sky130_fd_sc_hs__nor2_1_21/B sky130_fd_sc_hs__inv_4_31/Y sky130_fd_sc_hs__a21oi_1_33/a_117_74#
+ sky130_fd_sc_hs__a21oi_1_33/a_29_368# sky130_fd_sc_hs__a21oi_1
Xsky130_fd_sc_hs__a21oi_1_88 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nor2_1_87/Y sky130_fd_sc_hs__dfrtn_1_23/D
+ sky130_fd_sc_hs__nor2_1_87/B sky130_fd_sc_hs__inv_4_81/Y sky130_fd_sc_hs__a21oi_1_89/a_117_74#
+ sky130_fd_sc_hs__a21oi_1_89/a_29_368# sky130_fd_sc_hs__a21oi_1
Xsky130_fd_sc_hs__a21oi_1_77 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nor4_1_1/D sky130_fd_sc_hs__a31oi_2_1/A1
+ sky130_fd_sc_hs__nand2_1_59/Y sky130_fd_sc_hs__nor4_1_1/C sky130_fd_sc_hs__a21oi_1_77/a_117_74#
+ sky130_fd_sc_hs__a21oi_1_77/a_29_368# sky130_fd_sc_hs__a21oi_1
Xsky130_fd_sc_hs__a21oi_1_66 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nor2_1_47/Y sky130_fd_sc_hs__dfrtn_1_15/D
+ sky130_fd_sc_hs__nor2_1_47/B sky130_fd_sc_hs__inv_4_65/Y sky130_fd_sc_hs__a21oi_1_67/a_117_74#
+ sky130_fd_sc_hs__a21oi_1_67/a_29_368# sky130_fd_sc_hs__a21oi_1
Xsky130_fd_sc_hs__a21oi_1_99 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nor3_1_9/C sky130_fd_sc_hs__o22ai_1_9/A1
+ sky130_fd_sc_hs__o211ai_1_9/C1 sky130_fd_sc_hs__nor3_1_9/B sky130_fd_sc_hs__a21oi_1_99/a_117_74#
+ sky130_fd_sc_hs__a21oi_1_99/a_29_368# sky130_fd_sc_hs__a21oi_1
Xsky130_fd_sc_hs__a211oi_4_0 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__clkbuf_8_1/A sky130_fd_sc_hs__o22ai_1_1/Y
+ rst sky130_fd_sc_hs__o31ai_1_1/Y sky130_fd_sc_hs__inv_4_33/Y sky130_fd_sc_hs__a211oi_4_1/a_901_368#
+ sky130_fd_sc_hs__a211oi_4_1/a_77_368# sky130_fd_sc_hs__a211oi_4_1/a_92_74# sky130_fd_sc_hs__a211oi_4
Xsky130_fd_sc_hs__nand2b_1_9 DVSS DVDD DVDD DVSS rst sky130_fd_sc_hs__nor2_1_81/Y
+ sky130_fd_sc_hs__nor2b_1_41/A sky130_fd_sc_hs__nand2b_1_9/a_269_74# sky130_fd_sc_hs__nand2b_1_9/a_27_112#
+ sky130_fd_sc_hs__nand2b_1
Xsky130_fd_sc_hs__a32oi_1_8 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_1_51/Y sky130_fd_sc_hs__o21ai_1_5/B1
+ sky130_fd_sc_hs__o22ai_1_3/Y sky130_fd_sc_hs__o21ai_1_5/B1 sky130_fd_sc_hs__a32oi_1_9/Y
+ sky130_fd_sc_hs__o31ai_1_3/Y sky130_fd_sc_hs__a32oi_1_9/a_391_74# sky130_fd_sc_hs__a32oi_1_9/a_27_368#
+ sky130_fd_sc_hs__a32oi_1_9/a_119_74# sky130_fd_sc_hs__a32oi_1_9/a_469_74# sky130_fd_sc_hs__a32oi_1
Xsky130_fd_sc_hs__o21a_1_4 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__o21a_1_5/X sky130_fd_sc_hs__nor2_1_3/Y
+ sky130_fd_sc_hs__o21a_1_5/B1 sky130_fd_sc_hs__o21a_1_5/A1 sky130_fd_sc_hs__o21a_1_5/a_320_74#
+ sky130_fd_sc_hs__o21a_1_5/a_376_387# sky130_fd_sc_hs__o21a_1_5/a_83_244# sky130_fd_sc_hs__o21a_1
Xsky130_fd_sc_hs__fa_2_23 DVSS DVDD sky130_fd_sc_hs__fa_2_9/B DVDD DVSS sky130_fd_sc_hs__fa_2_23/CIN
+ sky130_fd_sc_hs__fa_2_23/B sky130_fd_sc_hs__fa_2_15/CIN sky130_fd_sc_hs__fa_2_23/SUM
+ sky130_fd_sc_hs__fa_2_23/a_27_378# sky130_fd_sc_hs__fa_2_23/a_701_79# sky130_fd_sc_hs__fa_2_23/a_484_347#
+ sky130_fd_sc_hs__fa_2_23/a_1094_347# sky130_fd_sc_hs__fa_2_23/a_1205_79# sky130_fd_sc_hs__fa_2_23/a_27_79#
+ sky130_fd_sc_hs__fa_2_23/a_1202_368# sky130_fd_sc_hs__fa_2_23/a_336_347# sky130_fd_sc_hs__fa_2_23/a_992_347#
+ sky130_fd_sc_hs__fa_2_23/a_1119_79# sky130_fd_sc_hs__fa_2_23/a_487_79# sky130_fd_sc_hs__fa_2_23/a_683_347#
+ sky130_fd_sc_hs__fa_2
Xsky130_fd_sc_hs__fa_2_12 DVSS DVDD sky130_fd_sc_hs__fa_2_9/B DVDD DVSS sky130_fd_sc_hs__fa_2_13/CIN
+ sky130_fd_sc_hs__fa_2_13/B sky130_fd_sc_hs__fa_2_17/CIN sky130_fd_sc_hs__fa_2_13/SUM
+ sky130_fd_sc_hs__fa_2_13/a_27_378# sky130_fd_sc_hs__fa_2_13/a_701_79# sky130_fd_sc_hs__fa_2_13/a_484_347#
+ sky130_fd_sc_hs__fa_2_13/a_1094_347# sky130_fd_sc_hs__fa_2_13/a_1205_79# sky130_fd_sc_hs__fa_2_13/a_27_79#
+ sky130_fd_sc_hs__fa_2_13/a_1202_368# sky130_fd_sc_hs__fa_2_13/a_336_347# sky130_fd_sc_hs__fa_2_13/a_992_347#
+ sky130_fd_sc_hs__fa_2_13/a_1119_79# sky130_fd_sc_hs__fa_2_13/a_487_79# sky130_fd_sc_hs__fa_2_13/a_683_347#
+ sky130_fd_sc_hs__fa_2
Xsky130_fd_sc_hs__dfrtn_1_9 DVSS DVDD sky130_fd_sc_hs__clkbuf_8_1/X DVDD DVSS sky130_fd_sc_hs__clkbuf_2_1/X
+ sky130_fd_sc_hs__nor2_1_65/A sky130_fd_sc_hs__o21a_1_37/X sky130_fd_sc_hs__dfrtn_1_9/a_1266_119#
+ sky130_fd_sc_hs__dfrtn_1_9/a_1736_119# sky130_fd_sc_hs__dfrtn_1_9/a_817_508# sky130_fd_sc_hs__dfrtn_1_9/a_120_74#
+ sky130_fd_sc_hs__dfrtn_1_9/a_1547_508# sky130_fd_sc_hs__dfrtn_1_9/a_922_127# sky130_fd_sc_hs__dfrtn_1_9/a_33_74#
+ sky130_fd_sc_hs__dfrtn_1_9/a_714_127# sky130_fd_sc_hs__dfrtn_1_9/a_1934_94# sky130_fd_sc_hs__dfrtn_1_9/a_1550_119#
+ sky130_fd_sc_hs__dfrtn_1_9/a_1598_93# sky130_fd_sc_hs__dfrtn_1_9/a_300_74# sky130_fd_sc_hs__dfrtn_1_9/a_507_368#
+ sky130_fd_sc_hs__dfrtn_1_9/a_856_304# sky130_fd_sc_hs__dfrtn_1_9/a_850_127# sky130_fd_sc_hs__dfrtn_1
Xsky130_fd_sc_hs__o211ai_1_9 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_109/A sky130_fd_sc_hs__o22ai_1_9/B1
+ sky130_fd_sc_hs__o211ai_1_9/C1 sky130_fd_sc_hs__inv_4_107/Y sky130_fd_sc_hs__inv_4_105/A
+ sky130_fd_sc_hs__o211ai_1_9/a_31_74# sky130_fd_sc_hs__o211ai_1_9/a_311_74# sky130_fd_sc_hs__o211ai_1_9/a_116_368#
+ sky130_fd_sc_hs__o211ai_1
Xsky130_fd_sc_hs__o21a_1_41 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__o21a_1_41/X sky130_fd_sc_hs__nor2_1_63/Y
+ sky130_fd_sc_hs__nor2_1_43/B sky130_fd_sc_hs__dfrbp_1_7/Q sky130_fd_sc_hs__o21a_1_41/a_320_74#
+ sky130_fd_sc_hs__o21a_1_41/a_376_387# sky130_fd_sc_hs__o21a_1_41/a_83_244# sky130_fd_sc_hs__o21a_1
Xsky130_fd_sc_hs__o21a_1_30 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__o21a_1_31/X sky130_fd_sc_hs__nor2_1_35/Y
+ sky130_fd_sc_hs__nor2_1_37/B sky130_fd_sc_hs__o21ai_1_3/B1 sky130_fd_sc_hs__o21a_1_31/a_320_74#
+ sky130_fd_sc_hs__o21a_1_31/a_376_387# sky130_fd_sc_hs__o21a_1_31/a_83_244# sky130_fd_sc_hs__o21a_1
Xsky130_fd_sc_hs__o21a_1_63 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__o21a_1_63/X sky130_fd_sc_hs__o21a_1_63/A2
+ sky130_fd_sc_hs__nor2_1_63/B sky130_fd_sc_hs__o21a_1_63/A1 sky130_fd_sc_hs__o21a_1_63/a_320_74#
+ sky130_fd_sc_hs__o21a_1_63/a_376_387# sky130_fd_sc_hs__o21a_1_63/a_83_244# sky130_fd_sc_hs__o21a_1
Xsky130_fd_sc_hs__o21a_1_74 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__o21a_1_75/X sky130_fd_sc_hs__o21a_1_75/A2
+ sky130_fd_sc_hs__o21a_1_75/B1 sky130_fd_sc_hs__o21a_1_75/A1 sky130_fd_sc_hs__o21a_1_75/a_320_74#
+ sky130_fd_sc_hs__o21a_1_75/a_376_387# sky130_fd_sc_hs__o21a_1_75/a_83_244# sky130_fd_sc_hs__o21a_1
Xsky130_fd_sc_hs__o21a_1_52 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__o21a_1_53/X sky130_fd_sc_hs__nor2_1_73/Y
+ sky130_fd_sc_hs__o21a_1_53/B1 sky130_fd_sc_hs__o22ai_1_7/A1 sky130_fd_sc_hs__o21a_1_53/a_320_74#
+ sky130_fd_sc_hs__o21a_1_53/a_376_387# sky130_fd_sc_hs__o21a_1_53/a_83_244# sky130_fd_sc_hs__o21a_1
Xsky130_fd_sc_hs__dfrtp_4_53 DVSS DVDD sky130_fd_sc_hs__inv_4_49/Y DVDD DVSS sky130_fd_sc_hs__nor2b_1_9/Y
+ sky130_fd_sc_hs__dfstp_2_1/CLK sky130_fd_sc_hs__fa_2_11/B sky130_fd_sc_hs__dfrtp_4_53/a_37_78#
+ sky130_fd_sc_hs__dfrtp_4_53/a_494_366# sky130_fd_sc_hs__dfrtp_4_53/a_699_463# sky130_fd_sc_hs__dfrtp_4_53/a_313_74#
+ sky130_fd_sc_hs__dfrtp_4_53/a_1627_493# sky130_fd_sc_hs__dfrtp_4_53/a_1678_395#
+ sky130_fd_sc_hs__dfrtp_4_53/a_1827_81# sky130_fd_sc_hs__dfrtp_4_53/a_789_463# sky130_fd_sc_hs__dfrtp_4_53/a_1350_392#
+ sky130_fd_sc_hs__dfrtp_4_53/a_834_355# sky130_fd_sc_hs__dfrtp_4_53/a_812_138# sky130_fd_sc_hs__dfrtp_4_53/a_124_78#
+ sky130_fd_sc_hs__dfrtp_4_53/a_1647_81# sky130_fd_sc_hs__dfrtp_4_53/a_2010_409# sky130_fd_sc_hs__dfrtp_4_53/a_890_138#
+ sky130_fd_sc_hs__dfrtp_4
Xsky130_fd_sc_hs__dfrtp_4_42 DVSS DVDD sky130_fd_sc_hs__clkbuf_8_1/X DVDD DVSS sky130_fd_sc_hs__dfrtp_4_43/D
+ sky130_fd_sc_hs__nand2_1_47/B sky130_fd_sc_hs__inv_4_17/A sky130_fd_sc_hs__dfrtp_4_43/a_37_78#
+ sky130_fd_sc_hs__dfrtp_4_43/a_494_366# sky130_fd_sc_hs__dfrtp_4_43/a_699_463# sky130_fd_sc_hs__dfrtp_4_43/a_313_74#
+ sky130_fd_sc_hs__dfrtp_4_43/a_1627_493# sky130_fd_sc_hs__dfrtp_4_43/a_1678_395#
+ sky130_fd_sc_hs__dfrtp_4_43/a_1827_81# sky130_fd_sc_hs__dfrtp_4_43/a_789_463# sky130_fd_sc_hs__dfrtp_4_43/a_1350_392#
+ sky130_fd_sc_hs__dfrtp_4_43/a_834_355# sky130_fd_sc_hs__dfrtp_4_43/a_812_138# sky130_fd_sc_hs__dfrtp_4_43/a_124_78#
+ sky130_fd_sc_hs__dfrtp_4_43/a_1647_81# sky130_fd_sc_hs__dfrtp_4_43/a_2010_409# sky130_fd_sc_hs__dfrtp_4_43/a_890_138#
+ sky130_fd_sc_hs__dfrtp_4
Xsky130_fd_sc_hs__dfrtp_4_31 DVSS DVDD sky130_fd_sc_hs__clkbuf_8_1/X DVDD DVSS sky130_fd_sc_hs__dfrtp_4_31/D
+ sky130_fd_sc_hs__nand2_1_47/B sky130_fd_sc_hs__inv_4_19/A sky130_fd_sc_hs__dfrtp_4_31/a_37_78#
+ sky130_fd_sc_hs__dfrtp_4_31/a_494_366# sky130_fd_sc_hs__dfrtp_4_31/a_699_463# sky130_fd_sc_hs__dfrtp_4_31/a_313_74#
+ sky130_fd_sc_hs__dfrtp_4_31/a_1627_493# sky130_fd_sc_hs__dfrtp_4_31/a_1678_395#
+ sky130_fd_sc_hs__dfrtp_4_31/a_1827_81# sky130_fd_sc_hs__dfrtp_4_31/a_789_463# sky130_fd_sc_hs__dfrtp_4_31/a_1350_392#
+ sky130_fd_sc_hs__dfrtp_4_31/a_834_355# sky130_fd_sc_hs__dfrtp_4_31/a_812_138# sky130_fd_sc_hs__dfrtp_4_31/a_124_78#
+ sky130_fd_sc_hs__dfrtp_4_31/a_1647_81# sky130_fd_sc_hs__dfrtp_4_31/a_2010_409# sky130_fd_sc_hs__dfrtp_4_31/a_890_138#
+ sky130_fd_sc_hs__dfrtp_4
Xsky130_fd_sc_hs__dfrtp_4_20 DVSS DVDD sky130_fd_sc_hs__clkbuf_8_1/X DVDD DVSS sky130_fd_sc_hs__o21a_1_11/X
+ sky130_fd_sc_hs__nand2_1_47/B sky130_fd_sc_hs__nand2_1_9/A sky130_fd_sc_hs__dfrtp_4_21/a_37_78#
+ sky130_fd_sc_hs__dfrtp_4_21/a_494_366# sky130_fd_sc_hs__dfrtp_4_21/a_699_463# sky130_fd_sc_hs__dfrtp_4_21/a_313_74#
+ sky130_fd_sc_hs__dfrtp_4_21/a_1627_493# sky130_fd_sc_hs__dfrtp_4_21/a_1678_395#
+ sky130_fd_sc_hs__dfrtp_4_21/a_1827_81# sky130_fd_sc_hs__dfrtp_4_21/a_789_463# sky130_fd_sc_hs__dfrtp_4_21/a_1350_392#
+ sky130_fd_sc_hs__dfrtp_4_21/a_834_355# sky130_fd_sc_hs__dfrtp_4_21/a_812_138# sky130_fd_sc_hs__dfrtp_4_21/a_124_78#
+ sky130_fd_sc_hs__dfrtp_4_21/a_1647_81# sky130_fd_sc_hs__dfrtp_4_21/a_2010_409# sky130_fd_sc_hs__dfrtp_4_21/a_890_138#
+ sky130_fd_sc_hs__dfrtp_4
Xsky130_fd_sc_hs__dfrtp_4_86 DVSS DVDD sky130_fd_sc_hs__clkbuf_8_1/X DVDD DVSS sky130_fd_sc_hs__o21a_1_31/X
+ sky130_fd_sc_hs__nand2_1_47/B sky130_fd_sc_hs__o21ai_1_3/B1 sky130_fd_sc_hs__dfrtp_4_87/a_37_78#
+ sky130_fd_sc_hs__dfrtp_4_87/a_494_366# sky130_fd_sc_hs__dfrtp_4_87/a_699_463# sky130_fd_sc_hs__dfrtp_4_87/a_313_74#
+ sky130_fd_sc_hs__dfrtp_4_87/a_1627_493# sky130_fd_sc_hs__dfrtp_4_87/a_1678_395#
+ sky130_fd_sc_hs__dfrtp_4_87/a_1827_81# sky130_fd_sc_hs__dfrtp_4_87/a_789_463# sky130_fd_sc_hs__dfrtp_4_87/a_1350_392#
+ sky130_fd_sc_hs__dfrtp_4_87/a_834_355# sky130_fd_sc_hs__dfrtp_4_87/a_812_138# sky130_fd_sc_hs__dfrtp_4_87/a_124_78#
+ sky130_fd_sc_hs__dfrtp_4_87/a_1647_81# sky130_fd_sc_hs__dfrtp_4_87/a_2010_409# sky130_fd_sc_hs__dfrtp_4_87/a_890_138#
+ sky130_fd_sc_hs__dfrtp_4
Xsky130_fd_sc_hs__dfrtp_4_75 DVSS DVDD sky130_fd_sc_hs__inv_4_49/Y DVDD DVSS sky130_fd_sc_hs__nor2b_1_17/Y
+ sky130_fd_sc_hs__dfstp_2_1/CLK sky130_fd_sc_hs__fa_2_17/B sky130_fd_sc_hs__dfrtp_4_75/a_37_78#
+ sky130_fd_sc_hs__dfrtp_4_75/a_494_366# sky130_fd_sc_hs__dfrtp_4_75/a_699_463# sky130_fd_sc_hs__dfrtp_4_75/a_313_74#
+ sky130_fd_sc_hs__dfrtp_4_75/a_1627_493# sky130_fd_sc_hs__dfrtp_4_75/a_1678_395#
+ sky130_fd_sc_hs__dfrtp_4_75/a_1827_81# sky130_fd_sc_hs__dfrtp_4_75/a_789_463# sky130_fd_sc_hs__dfrtp_4_75/a_1350_392#
+ sky130_fd_sc_hs__dfrtp_4_75/a_834_355# sky130_fd_sc_hs__dfrtp_4_75/a_812_138# sky130_fd_sc_hs__dfrtp_4_75/a_124_78#
+ sky130_fd_sc_hs__dfrtp_4_75/a_1647_81# sky130_fd_sc_hs__dfrtp_4_75/a_2010_409# sky130_fd_sc_hs__dfrtp_4_75/a_890_138#
+ sky130_fd_sc_hs__dfrtp_4
Xsky130_fd_sc_hs__dfrtp_4_64 DVSS DVDD sky130_fd_sc_hs__clkbuf_8_1/X DVDD DVSS sky130_fd_sc_hs__o21a_1_27/X
+ sky130_fd_sc_hs__nand2_1_47/B sky130_fd_sc_hs__o21a_1_27/A1 sky130_fd_sc_hs__dfrtp_4_65/a_37_78#
+ sky130_fd_sc_hs__dfrtp_4_65/a_494_366# sky130_fd_sc_hs__dfrtp_4_65/a_699_463# sky130_fd_sc_hs__dfrtp_4_65/a_313_74#
+ sky130_fd_sc_hs__dfrtp_4_65/a_1627_493# sky130_fd_sc_hs__dfrtp_4_65/a_1678_395#
+ sky130_fd_sc_hs__dfrtp_4_65/a_1827_81# sky130_fd_sc_hs__dfrtp_4_65/a_789_463# sky130_fd_sc_hs__dfrtp_4_65/a_1350_392#
+ sky130_fd_sc_hs__dfrtp_4_65/a_834_355# sky130_fd_sc_hs__dfrtp_4_65/a_812_138# sky130_fd_sc_hs__dfrtp_4_65/a_124_78#
+ sky130_fd_sc_hs__dfrtp_4_65/a_1647_81# sky130_fd_sc_hs__dfrtp_4_65/a_2010_409# sky130_fd_sc_hs__dfrtp_4_65/a_890_138#
+ sky130_fd_sc_hs__dfrtp_4
Xsky130_fd_sc_hs__a22o_1_8 DVSS DVDD DVDD DVSS osc_fine_con_final[4] manual_control_osc[4]
+ sky130_fd_sc_hs__inv_4_43/Y sky130_fd_sc_hs__fa_2_7/B fftl_en sky130_fd_sc_hs__a22o_1_9/a_222_392#
+ sky130_fd_sc_hs__a22o_1_9/a_230_79# sky130_fd_sc_hs__a22o_1_9/a_52_123# sky130_fd_sc_hs__a22o_1_9/a_132_392#
+ sky130_fd_sc_hs__a22o_1
Xsky130_fd_sc_hs__a2bb2oi_1_0 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__a2bb2oi_1_1/Y sky130_fd_sc_hs__inv_2_5/A
+ sky130_fd_sc_hs__inv_2_9/Y div_ratio_half[0] sky130_fd_sc_hs__inv_2_3/A sky130_fd_sc_hs__a2bb2oi_1_1/a_399_368#
+ sky130_fd_sc_hs__a2bb2oi_1_1/a_126_112# sky130_fd_sc_hs__a2bb2oi_1_1/a_117_392#
+ sky130_fd_sc_hs__a2bb2oi_1_1/a_488_74# sky130_fd_sc_hs__a2bb2oi_1
Xsky130_fd_sc_hs__nor2b_1_6 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__fa_2_7/SUM sky130_fd_sc_hs__nor2b_1_7/Y
+ sky130_fd_sc_hs__or2_1_1/A sky130_fd_sc_hs__nor2b_1_7/a_278_368# sky130_fd_sc_hs__nor2b_1_7/a_27_112#
+ sky130_fd_sc_hs__nor2b_1
Xsky130_fd_sc_hs__nand2_1_8 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nor2_1_15/Y sky130_fd_sc_hs__nor2_1_13/B
+ sky130_fd_sc_hs__nand2_1_9/A sky130_fd_sc_hs__nand2_1_9/a_117_74# sky130_fd_sc_hs__nand2_1
Xsky130_fd_sc_hs__nor2_1_4 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nor2_1_5/B sky130_fd_sc_hs__nor2_1_5/Y
+ sky130_fd_sc_hs__inv_4_7/Y sky130_fd_sc_hs__nor2_1_5/a_116_368# sky130_fd_sc_hs__nor2_1
Xsky130_fd_sc_hs__a21oi_1_12 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nor2_1_15/Y sky130_fd_sc_hs__dfrtp_4_31/D
+ sky130_fd_sc_hs__nor2_1_15/B sky130_fd_sc_hs__inv_4_19/Y sky130_fd_sc_hs__a21oi_1_13/a_117_74#
+ sky130_fd_sc_hs__a21oi_1_13/a_29_368# sky130_fd_sc_hs__a21oi_1
Xsky130_fd_sc_hs__a21oi_1_56 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nor2_1_51/Y sky130_fd_sc_hs__dfrbp_1_3/D
+ sky130_fd_sc_hs__nor2_1_51/B sky130_fd_sc_hs__inv_4_61/Y sky130_fd_sc_hs__a21oi_1_57/a_117_74#
+ sky130_fd_sc_hs__a21oi_1_57/a_29_368# sky130_fd_sc_hs__a21oi_1
Xsky130_fd_sc_hs__a21oi_1_45 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nor2_1_31/Y sky130_fd_sc_hs__dfrtp_4_83/D
+ sky130_fd_sc_hs__nor2_1_31/B sky130_fd_sc_hs__inv_4_45/Y sky130_fd_sc_hs__a21oi_1_45/a_117_74#
+ sky130_fd_sc_hs__a21oi_1_45/a_29_368# sky130_fd_sc_hs__a21oi_1
Xsky130_fd_sc_hs__a21oi_1_34 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__a222o_1_1/X sky130_fd_sc_hs__a32oi_1_7/B1
+ sky130_fd_sc_hs__nor2_1_33/Y sky130_fd_sc_hs__inv_4_5/A sky130_fd_sc_hs__a21oi_1_35/a_117_74#
+ sky130_fd_sc_hs__a21oi_1_35/a_29_368# sky130_fd_sc_hs__a21oi_1
Xsky130_fd_sc_hs__a21oi_1_23 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nor2_1_13/Y sky130_fd_sc_hs__dfrtp_4_43/D
+ sky130_fd_sc_hs__nor2_1_13/B sky130_fd_sc_hs__inv_4_17/Y sky130_fd_sc_hs__a21oi_1_23/a_117_74#
+ sky130_fd_sc_hs__a21oi_1_23/a_29_368# sky130_fd_sc_hs__a21oi_1
Xsky130_fd_sc_hs__a21oi_1_89 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nor2_1_87/Y sky130_fd_sc_hs__dfrtn_1_23/D
+ sky130_fd_sc_hs__nor2_1_87/B sky130_fd_sc_hs__inv_4_81/Y sky130_fd_sc_hs__a21oi_1_89/a_117_74#
+ sky130_fd_sc_hs__a21oi_1_89/a_29_368# sky130_fd_sc_hs__a21oi_1
Xsky130_fd_sc_hs__a21oi_1_78 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__o21ai_1_5/Y sky130_fd_sc_hs__nand4_1_5/A
+ sky130_fd_sc_hs__inv_4_81/Y sky130_fd_sc_hs__inv_4_71/A sky130_fd_sc_hs__a21oi_1_79/a_117_74#
+ sky130_fd_sc_hs__a21oi_1_79/a_29_368# sky130_fd_sc_hs__a21oi_1
Xsky130_fd_sc_hs__a21oi_1_67 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nor2_1_47/Y sky130_fd_sc_hs__dfrtn_1_15/D
+ sky130_fd_sc_hs__nor2_1_47/B sky130_fd_sc_hs__inv_4_65/Y sky130_fd_sc_hs__a21oi_1_67/a_117_74#
+ sky130_fd_sc_hs__a21oi_1_67/a_29_368# sky130_fd_sc_hs__a21oi_1
Xsky130_fd_sc_hs__a211oi_4_1 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__clkbuf_8_1/A sky130_fd_sc_hs__o22ai_1_1/Y
+ rst sky130_fd_sc_hs__o31ai_1_1/Y sky130_fd_sc_hs__inv_4_33/Y sky130_fd_sc_hs__a211oi_4_1/a_901_368#
+ sky130_fd_sc_hs__a211oi_4_1/a_77_368# sky130_fd_sc_hs__a211oi_4_1/a_92_74# sky130_fd_sc_hs__a211oi_4
Xsky130_fd_sc_hs__a32oi_1_9 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_1_51/Y sky130_fd_sc_hs__o21ai_1_5/B1
+ sky130_fd_sc_hs__o22ai_1_3/Y sky130_fd_sc_hs__o21ai_1_5/B1 sky130_fd_sc_hs__a32oi_1_9/Y
+ sky130_fd_sc_hs__o31ai_1_3/Y sky130_fd_sc_hs__a32oi_1_9/a_391_74# sky130_fd_sc_hs__a32oi_1_9/a_27_368#
+ sky130_fd_sc_hs__a32oi_1_9/a_119_74# sky130_fd_sc_hs__a32oi_1_9/a_469_74# sky130_fd_sc_hs__a32oi_1
Xsky130_fd_sc_hs__o21a_1_5 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__o21a_1_5/X sky130_fd_sc_hs__nor2_1_3/Y
+ sky130_fd_sc_hs__o21a_1_5/B1 sky130_fd_sc_hs__o21a_1_5/A1 sky130_fd_sc_hs__o21a_1_5/a_320_74#
+ sky130_fd_sc_hs__o21a_1_5/a_376_387# sky130_fd_sc_hs__o21a_1_5/a_83_244# sky130_fd_sc_hs__o21a_1
Xsky130_fd_sc_hs__fa_2_13 DVSS DVDD sky130_fd_sc_hs__fa_2_9/B DVDD DVSS sky130_fd_sc_hs__fa_2_13/CIN
+ sky130_fd_sc_hs__fa_2_13/B sky130_fd_sc_hs__fa_2_17/CIN sky130_fd_sc_hs__fa_2_13/SUM
+ sky130_fd_sc_hs__fa_2_13/a_27_378# sky130_fd_sc_hs__fa_2_13/a_701_79# sky130_fd_sc_hs__fa_2_13/a_484_347#
+ sky130_fd_sc_hs__fa_2_13/a_1094_347# sky130_fd_sc_hs__fa_2_13/a_1205_79# sky130_fd_sc_hs__fa_2_13/a_27_79#
+ sky130_fd_sc_hs__fa_2_13/a_1202_368# sky130_fd_sc_hs__fa_2_13/a_336_347# sky130_fd_sc_hs__fa_2_13/a_992_347#
+ sky130_fd_sc_hs__fa_2_13/a_1119_79# sky130_fd_sc_hs__fa_2_13/a_487_79# sky130_fd_sc_hs__fa_2_13/a_683_347#
+ sky130_fd_sc_hs__fa_2
Xsky130_fd_sc_hs__o21a_1_42 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__o21a_1_43/X sky130_fd_sc_hs__nor2_1_43/Y
+ sky130_fd_sc_hs__nor2_1_41/B sky130_fd_sc_hs__inv_4_73/A sky130_fd_sc_hs__o21a_1_43/a_320_74#
+ sky130_fd_sc_hs__o21a_1_43/a_376_387# sky130_fd_sc_hs__o21a_1_43/a_83_244# sky130_fd_sc_hs__o21a_1
Xsky130_fd_sc_hs__o21a_1_31 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__o21a_1_31/X sky130_fd_sc_hs__nor2_1_35/Y
+ sky130_fd_sc_hs__nor2_1_37/B sky130_fd_sc_hs__o21ai_1_3/B1 sky130_fd_sc_hs__o21a_1_31/a_320_74#
+ sky130_fd_sc_hs__o21a_1_31/a_376_387# sky130_fd_sc_hs__o21a_1_31/a_83_244# sky130_fd_sc_hs__o21a_1
Xsky130_fd_sc_hs__o21a_1_20 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__o21a_1_21/X sky130_fd_sc_hs__nor2_1_13/Y
+ sky130_fd_sc_hs__nor2_1_25/B sky130_fd_sc_hs__o21a_1_21/A1 sky130_fd_sc_hs__o21a_1_21/a_320_74#
+ sky130_fd_sc_hs__o21a_1_21/a_376_387# sky130_fd_sc_hs__o21a_1_21/a_83_244# sky130_fd_sc_hs__o21a_1
Xsky130_fd_sc_hs__o21a_1_64 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__o21a_1_65/X sky130_fd_sc_hs__nor2_1_99/Y
+ sky130_fd_sc_hs__o21a_1_65/B1 sky130_fd_sc_hs__inv_4_101/A sky130_fd_sc_hs__o21a_1_65/a_320_74#
+ sky130_fd_sc_hs__o21a_1_65/a_376_387# sky130_fd_sc_hs__o21a_1_65/a_83_244# sky130_fd_sc_hs__o21a_1
Xsky130_fd_sc_hs__o21a_1_75 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__o21a_1_75/X sky130_fd_sc_hs__o21a_1_75/A2
+ sky130_fd_sc_hs__o21a_1_75/B1 sky130_fd_sc_hs__o21a_1_75/A1 sky130_fd_sc_hs__o21a_1_75/a_320_74#
+ sky130_fd_sc_hs__o21a_1_75/a_376_387# sky130_fd_sc_hs__o21a_1_75/a_83_244# sky130_fd_sc_hs__o21a_1
Xsky130_fd_sc_hs__o21a_1_53 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__o21a_1_53/X sky130_fd_sc_hs__nor2_1_73/Y
+ sky130_fd_sc_hs__o21a_1_53/B1 sky130_fd_sc_hs__o22ai_1_7/A1 sky130_fd_sc_hs__o21a_1_53/a_320_74#
+ sky130_fd_sc_hs__o21a_1_53/a_376_387# sky130_fd_sc_hs__o21a_1_53/a_83_244# sky130_fd_sc_hs__o21a_1
Xsky130_fd_sc_hs__dfrtp_4_10 DVSS DVDD sky130_fd_sc_hs__clkbuf_8_1/X DVDD DVSS sky130_fd_sc_hs__a21oi_1_1/Y
+ sky130_fd_sc_hs__nand2_1_47/B sky130_fd_sc_hs__inv_4_5/A sky130_fd_sc_hs__dfrtp_4_11/a_37_78#
+ sky130_fd_sc_hs__dfrtp_4_11/a_494_366# sky130_fd_sc_hs__dfrtp_4_11/a_699_463# sky130_fd_sc_hs__dfrtp_4_11/a_313_74#
+ sky130_fd_sc_hs__dfrtp_4_11/a_1627_493# sky130_fd_sc_hs__dfrtp_4_11/a_1678_395#
+ sky130_fd_sc_hs__dfrtp_4_11/a_1827_81# sky130_fd_sc_hs__dfrtp_4_11/a_789_463# sky130_fd_sc_hs__dfrtp_4_11/a_1350_392#
+ sky130_fd_sc_hs__dfrtp_4_11/a_834_355# sky130_fd_sc_hs__dfrtp_4_11/a_812_138# sky130_fd_sc_hs__dfrtp_4_11/a_124_78#
+ sky130_fd_sc_hs__dfrtp_4_11/a_1647_81# sky130_fd_sc_hs__dfrtp_4_11/a_2010_409# sky130_fd_sc_hs__dfrtp_4_11/a_890_138#
+ sky130_fd_sc_hs__dfrtp_4
Xsky130_fd_sc_hs__dfrtp_4_43 DVSS DVDD sky130_fd_sc_hs__clkbuf_8_1/X DVDD DVSS sky130_fd_sc_hs__dfrtp_4_43/D
+ sky130_fd_sc_hs__nand2_1_47/B sky130_fd_sc_hs__inv_4_17/A sky130_fd_sc_hs__dfrtp_4_43/a_37_78#
+ sky130_fd_sc_hs__dfrtp_4_43/a_494_366# sky130_fd_sc_hs__dfrtp_4_43/a_699_463# sky130_fd_sc_hs__dfrtp_4_43/a_313_74#
+ sky130_fd_sc_hs__dfrtp_4_43/a_1627_493# sky130_fd_sc_hs__dfrtp_4_43/a_1678_395#
+ sky130_fd_sc_hs__dfrtp_4_43/a_1827_81# sky130_fd_sc_hs__dfrtp_4_43/a_789_463# sky130_fd_sc_hs__dfrtp_4_43/a_1350_392#
+ sky130_fd_sc_hs__dfrtp_4_43/a_834_355# sky130_fd_sc_hs__dfrtp_4_43/a_812_138# sky130_fd_sc_hs__dfrtp_4_43/a_124_78#
+ sky130_fd_sc_hs__dfrtp_4_43/a_1647_81# sky130_fd_sc_hs__dfrtp_4_43/a_2010_409# sky130_fd_sc_hs__dfrtp_4_43/a_890_138#
+ sky130_fd_sc_hs__dfrtp_4
Xsky130_fd_sc_hs__dfrtp_4_32 DVSS DVDD sky130_fd_sc_hs__clkbuf_8_1/X DVDD DVSS sky130_fd_sc_hs__a21oi_1_9/Y
+ sky130_fd_sc_hs__nand2_1_47/B sky130_fd_sc_hs__inv_4_11/A sky130_fd_sc_hs__dfrtp_4_33/a_37_78#
+ sky130_fd_sc_hs__dfrtp_4_33/a_494_366# sky130_fd_sc_hs__dfrtp_4_33/a_699_463# sky130_fd_sc_hs__dfrtp_4_33/a_313_74#
+ sky130_fd_sc_hs__dfrtp_4_33/a_1627_493# sky130_fd_sc_hs__dfrtp_4_33/a_1678_395#
+ sky130_fd_sc_hs__dfrtp_4_33/a_1827_81# sky130_fd_sc_hs__dfrtp_4_33/a_789_463# sky130_fd_sc_hs__dfrtp_4_33/a_1350_392#
+ sky130_fd_sc_hs__dfrtp_4_33/a_834_355# sky130_fd_sc_hs__dfrtp_4_33/a_812_138# sky130_fd_sc_hs__dfrtp_4_33/a_124_78#
+ sky130_fd_sc_hs__dfrtp_4_33/a_1647_81# sky130_fd_sc_hs__dfrtp_4_33/a_2010_409# sky130_fd_sc_hs__dfrtp_4_33/a_890_138#
+ sky130_fd_sc_hs__dfrtp_4
Xsky130_fd_sc_hs__dfrtp_4_21 DVSS DVDD sky130_fd_sc_hs__clkbuf_8_1/X DVDD DVSS sky130_fd_sc_hs__o21a_1_11/X
+ sky130_fd_sc_hs__nand2_1_47/B sky130_fd_sc_hs__nand2_1_9/A sky130_fd_sc_hs__dfrtp_4_21/a_37_78#
+ sky130_fd_sc_hs__dfrtp_4_21/a_494_366# sky130_fd_sc_hs__dfrtp_4_21/a_699_463# sky130_fd_sc_hs__dfrtp_4_21/a_313_74#
+ sky130_fd_sc_hs__dfrtp_4_21/a_1627_493# sky130_fd_sc_hs__dfrtp_4_21/a_1678_395#
+ sky130_fd_sc_hs__dfrtp_4_21/a_1827_81# sky130_fd_sc_hs__dfrtp_4_21/a_789_463# sky130_fd_sc_hs__dfrtp_4_21/a_1350_392#
+ sky130_fd_sc_hs__dfrtp_4_21/a_834_355# sky130_fd_sc_hs__dfrtp_4_21/a_812_138# sky130_fd_sc_hs__dfrtp_4_21/a_124_78#
+ sky130_fd_sc_hs__dfrtp_4_21/a_1647_81# sky130_fd_sc_hs__dfrtp_4_21/a_2010_409# sky130_fd_sc_hs__dfrtp_4_21/a_890_138#
+ sky130_fd_sc_hs__dfrtp_4
Xsky130_fd_sc_hs__dfrtp_4_76 DVSS DVDD sky130_fd_sc_hs__clkbuf_8_1/A DVDD DVSS sky130_fd_sc_hs__dfrtp_4_77/D
+ sky130_fd_sc_hs__nand2_1_47/B sky130_fd_sc_hs__inv_4_35/A sky130_fd_sc_hs__dfrtp_4_77/a_37_78#
+ sky130_fd_sc_hs__dfrtp_4_77/a_494_366# sky130_fd_sc_hs__dfrtp_4_77/a_699_463# sky130_fd_sc_hs__dfrtp_4_77/a_313_74#
+ sky130_fd_sc_hs__dfrtp_4_77/a_1627_493# sky130_fd_sc_hs__dfrtp_4_77/a_1678_395#
+ sky130_fd_sc_hs__dfrtp_4_77/a_1827_81# sky130_fd_sc_hs__dfrtp_4_77/a_789_463# sky130_fd_sc_hs__dfrtp_4_77/a_1350_392#
+ sky130_fd_sc_hs__dfrtp_4_77/a_834_355# sky130_fd_sc_hs__dfrtp_4_77/a_812_138# sky130_fd_sc_hs__dfrtp_4_77/a_124_78#
+ sky130_fd_sc_hs__dfrtp_4_77/a_1647_81# sky130_fd_sc_hs__dfrtp_4_77/a_2010_409# sky130_fd_sc_hs__dfrtp_4_77/a_890_138#
+ sky130_fd_sc_hs__dfrtp_4
Xsky130_fd_sc_hs__dfrtp_4_65 DVSS DVDD sky130_fd_sc_hs__clkbuf_8_1/X DVDD DVSS sky130_fd_sc_hs__o21a_1_27/X
+ sky130_fd_sc_hs__nand2_1_47/B sky130_fd_sc_hs__o21a_1_27/A1 sky130_fd_sc_hs__dfrtp_4_65/a_37_78#
+ sky130_fd_sc_hs__dfrtp_4_65/a_494_366# sky130_fd_sc_hs__dfrtp_4_65/a_699_463# sky130_fd_sc_hs__dfrtp_4_65/a_313_74#
+ sky130_fd_sc_hs__dfrtp_4_65/a_1627_493# sky130_fd_sc_hs__dfrtp_4_65/a_1678_395#
+ sky130_fd_sc_hs__dfrtp_4_65/a_1827_81# sky130_fd_sc_hs__dfrtp_4_65/a_789_463# sky130_fd_sc_hs__dfrtp_4_65/a_1350_392#
+ sky130_fd_sc_hs__dfrtp_4_65/a_834_355# sky130_fd_sc_hs__dfrtp_4_65/a_812_138# sky130_fd_sc_hs__dfrtp_4_65/a_124_78#
+ sky130_fd_sc_hs__dfrtp_4_65/a_1647_81# sky130_fd_sc_hs__dfrtp_4_65/a_2010_409# sky130_fd_sc_hs__dfrtp_4_65/a_890_138#
+ sky130_fd_sc_hs__dfrtp_4
Xsky130_fd_sc_hs__dfrtp_4_54 DVSS DVDD sky130_fd_sc_hs__clkbuf_8_1/A DVDD DVSS sky130_fd_sc_hs__o21a_1_23/X
+ sky130_fd_sc_hs__nand2_1_47/B sky130_fd_sc_hs__o21a_1_23/A1 sky130_fd_sc_hs__dfrtp_4_55/a_37_78#
+ sky130_fd_sc_hs__dfrtp_4_55/a_494_366# sky130_fd_sc_hs__dfrtp_4_55/a_699_463# sky130_fd_sc_hs__dfrtp_4_55/a_313_74#
+ sky130_fd_sc_hs__dfrtp_4_55/a_1627_493# sky130_fd_sc_hs__dfrtp_4_55/a_1678_395#
+ sky130_fd_sc_hs__dfrtp_4_55/a_1827_81# sky130_fd_sc_hs__dfrtp_4_55/a_789_463# sky130_fd_sc_hs__dfrtp_4_55/a_1350_392#
+ sky130_fd_sc_hs__dfrtp_4_55/a_834_355# sky130_fd_sc_hs__dfrtp_4_55/a_812_138# sky130_fd_sc_hs__dfrtp_4_55/a_124_78#
+ sky130_fd_sc_hs__dfrtp_4_55/a_1647_81# sky130_fd_sc_hs__dfrtp_4_55/a_2010_409# sky130_fd_sc_hs__dfrtp_4_55/a_890_138#
+ sky130_fd_sc_hs__dfrtp_4
Xsky130_fd_sc_hs__a22o_1_9 DVSS DVDD DVDD DVSS osc_fine_con_final[4] manual_control_osc[4]
+ sky130_fd_sc_hs__inv_4_43/Y sky130_fd_sc_hs__fa_2_7/B fftl_en sky130_fd_sc_hs__a22o_1_9/a_222_392#
+ sky130_fd_sc_hs__a22o_1_9/a_230_79# sky130_fd_sc_hs__a22o_1_9/a_52_123# sky130_fd_sc_hs__a22o_1_9/a_132_392#
+ sky130_fd_sc_hs__a22o_1
Xsky130_fd_sc_hs__dfrtp_4_87 DVSS DVDD sky130_fd_sc_hs__clkbuf_8_1/X DVDD DVSS sky130_fd_sc_hs__o21a_1_31/X
+ sky130_fd_sc_hs__nand2_1_47/B sky130_fd_sc_hs__o21ai_1_3/B1 sky130_fd_sc_hs__dfrtp_4_87/a_37_78#
+ sky130_fd_sc_hs__dfrtp_4_87/a_494_366# sky130_fd_sc_hs__dfrtp_4_87/a_699_463# sky130_fd_sc_hs__dfrtp_4_87/a_313_74#
+ sky130_fd_sc_hs__dfrtp_4_87/a_1627_493# sky130_fd_sc_hs__dfrtp_4_87/a_1678_395#
+ sky130_fd_sc_hs__dfrtp_4_87/a_1827_81# sky130_fd_sc_hs__dfrtp_4_87/a_789_463# sky130_fd_sc_hs__dfrtp_4_87/a_1350_392#
+ sky130_fd_sc_hs__dfrtp_4_87/a_834_355# sky130_fd_sc_hs__dfrtp_4_87/a_812_138# sky130_fd_sc_hs__dfrtp_4_87/a_124_78#
+ sky130_fd_sc_hs__dfrtp_4_87/a_1647_81# sky130_fd_sc_hs__dfrtp_4_87/a_2010_409# sky130_fd_sc_hs__dfrtp_4_87/a_890_138#
+ sky130_fd_sc_hs__dfrtp_4
Xsky130_fd_sc_hs__a2bb2oi_1_1 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__a2bb2oi_1_1/Y sky130_fd_sc_hs__inv_2_5/A
+ sky130_fd_sc_hs__inv_2_9/Y div_ratio_half[0] sky130_fd_sc_hs__inv_2_3/A sky130_fd_sc_hs__a2bb2oi_1_1/a_399_368#
+ sky130_fd_sc_hs__a2bb2oi_1_1/a_126_112# sky130_fd_sc_hs__a2bb2oi_1_1/a_117_392#
+ sky130_fd_sc_hs__a2bb2oi_1_1/a_488_74# sky130_fd_sc_hs__a2bb2oi_1
Xsky130_fd_sc_hs__nor2b_1_7 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__fa_2_7/SUM sky130_fd_sc_hs__nor2b_1_7/Y
+ sky130_fd_sc_hs__or2_1_1/A sky130_fd_sc_hs__nor2b_1_7/a_278_368# sky130_fd_sc_hs__nor2b_1_7/a_27_112#
+ sky130_fd_sc_hs__nor2b_1
Xsky130_fd_sc_hs__nand2_1_9 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nor2_1_15/Y sky130_fd_sc_hs__nor2_1_13/B
+ sky130_fd_sc_hs__nand2_1_9/A sky130_fd_sc_hs__nand2_1_9/a_117_74# sky130_fd_sc_hs__nand2_1
Xsky130_fd_sc_hs__nor2_1_5 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nor2_1_5/B sky130_fd_sc_hs__nor2_1_5/Y
+ sky130_fd_sc_hs__inv_4_7/Y sky130_fd_sc_hs__nor2_1_5/a_116_368# sky130_fd_sc_hs__nor2_1
Xsky130_fd_sc_hs__a21oi_1_13 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nor2_1_15/Y sky130_fd_sc_hs__dfrtp_4_31/D
+ sky130_fd_sc_hs__nor2_1_15/B sky130_fd_sc_hs__inv_4_19/Y sky130_fd_sc_hs__a21oi_1_13/a_117_74#
+ sky130_fd_sc_hs__a21oi_1_13/a_29_368# sky130_fd_sc_hs__a21oi_1
Xsky130_fd_sc_hs__a21oi_1_46 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nor2_1_37/Y sky130_fd_sc_hs__dfrtp_4_77/D
+ sky130_fd_sc_hs__nor2_1_37/B sky130_fd_sc_hs__inv_4_35/Y sky130_fd_sc_hs__a21oi_1_47/a_117_74#
+ sky130_fd_sc_hs__a21oi_1_47/a_29_368# sky130_fd_sc_hs__a21oi_1
Xsky130_fd_sc_hs__a21oi_1_35 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__a222o_1_1/X sky130_fd_sc_hs__a32oi_1_7/B1
+ sky130_fd_sc_hs__nor2_1_33/Y sky130_fd_sc_hs__inv_4_5/A sky130_fd_sc_hs__a21oi_1_35/a_117_74#
+ sky130_fd_sc_hs__a21oi_1_35/a_29_368# sky130_fd_sc_hs__a21oi_1
Xsky130_fd_sc_hs__a21oi_1_24 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__a21oi_1_15/Y sky130_fd_sc_hs__a32oi_1_3/B1
+ sky130_fd_sc_hs__a211oi_1_1/Y sky130_fd_sc_hs__a22oi_1_15/Y sky130_fd_sc_hs__a21oi_1_25/a_117_74#
+ sky130_fd_sc_hs__a21oi_1_25/a_29_368# sky130_fd_sc_hs__a21oi_1
Xsky130_fd_sc_hs__a21oi_1_79 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__o21ai_1_5/Y sky130_fd_sc_hs__nand4_1_5/A
+ sky130_fd_sc_hs__inv_4_81/Y sky130_fd_sc_hs__inv_4_71/A sky130_fd_sc_hs__a21oi_1_79/a_117_74#
+ sky130_fd_sc_hs__a21oi_1_79/a_29_368# sky130_fd_sc_hs__a21oi_1
Xsky130_fd_sc_hs__a21oi_1_68 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nor2_1_57/Y sky130_fd_sc_hs__dfrbp_1_11/D
+ sky130_fd_sc_hs__nor2_1_57/B sky130_fd_sc_hs__inv_4_79/Y sky130_fd_sc_hs__a21oi_1_69/a_117_74#
+ sky130_fd_sc_hs__a21oi_1_69/a_29_368# sky130_fd_sc_hs__a21oi_1
Xsky130_fd_sc_hs__a21oi_1_57 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nor2_1_51/Y sky130_fd_sc_hs__dfrbp_1_3/D
+ sky130_fd_sc_hs__nor2_1_51/B sky130_fd_sc_hs__inv_4_61/Y sky130_fd_sc_hs__a21oi_1_57/a_117_74#
+ sky130_fd_sc_hs__a21oi_1_57/a_29_368# sky130_fd_sc_hs__a21oi_1
Xsky130_fd_sc_hs__clkbuf_8_0 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__clkbuf_8_1/X sky130_fd_sc_hs__clkbuf_8_1/A
+ sky130_fd_sc_hs__clkbuf_8_1/a_125_368# sky130_fd_sc_hs__clkbuf_8
Xsky130_fd_sc_hs__o21a_1_6 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__o21a_1_7/X sky130_fd_sc_hs__o21a_1_7/A2
+ sky130_fd_sc_hs__nor2_1_5/B sky130_fd_sc_hs__o21a_1_7/A1 sky130_fd_sc_hs__o21a_1_7/a_320_74#
+ sky130_fd_sc_hs__o21a_1_7/a_376_387# sky130_fd_sc_hs__o21a_1_7/a_83_244# sky130_fd_sc_hs__o21a_1
Xsky130_fd_sc_hs__nor2_1_120 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__o21a_1_75/B1 sky130_fd_sc_hs__o21a_1_61/A2
+ sky130_fd_sc_hs__inv_4_135/Y sky130_fd_sc_hs__nor2_1_121/a_116_368# sky130_fd_sc_hs__nor2_1
Xsky130_fd_sc_hs__fa_2_14 DVSS DVDD sky130_fd_sc_hs__fa_2_9/B DVDD DVSS sky130_fd_sc_hs__fa_2_15/CIN
+ sky130_fd_sc_hs__fa_2_15/B sky130_fd_sc_hs__xor2_1_11/B sky130_fd_sc_hs__fa_2_15/SUM
+ sky130_fd_sc_hs__fa_2_15/a_27_378# sky130_fd_sc_hs__fa_2_15/a_701_79# sky130_fd_sc_hs__fa_2_15/a_484_347#
+ sky130_fd_sc_hs__fa_2_15/a_1094_347# sky130_fd_sc_hs__fa_2_15/a_1205_79# sky130_fd_sc_hs__fa_2_15/a_27_79#
+ sky130_fd_sc_hs__fa_2_15/a_1202_368# sky130_fd_sc_hs__fa_2_15/a_336_347# sky130_fd_sc_hs__fa_2_15/a_992_347#
+ sky130_fd_sc_hs__fa_2_15/a_1119_79# sky130_fd_sc_hs__fa_2_15/a_487_79# sky130_fd_sc_hs__fa_2_15/a_683_347#
+ sky130_fd_sc_hs__fa_2
Xsky130_fd_sc_hs__o21a_1_32 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__o21a_1_33/X sky130_fd_sc_hs__nor2_1_27/Y
+ sky130_fd_sc_hs__nor2_1_49/B sky130_fd_sc_hs__inv_4_55/A sky130_fd_sc_hs__o21a_1_33/a_320_74#
+ sky130_fd_sc_hs__o21a_1_33/a_376_387# sky130_fd_sc_hs__o21a_1_33/a_83_244# sky130_fd_sc_hs__o21a_1
Xsky130_fd_sc_hs__o21a_1_21 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__o21a_1_21/X sky130_fd_sc_hs__nor2_1_13/Y
+ sky130_fd_sc_hs__nor2_1_25/B sky130_fd_sc_hs__o21a_1_21/A1 sky130_fd_sc_hs__o21a_1_21/a_320_74#
+ sky130_fd_sc_hs__o21a_1_21/a_376_387# sky130_fd_sc_hs__o21a_1_21/a_83_244# sky130_fd_sc_hs__o21a_1
Xsky130_fd_sc_hs__o21a_1_10 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__o21a_1_11/X sky130_fd_sc_hs__nor2_1_15/Y
+ sky130_fd_sc_hs__nor2_1_13/B sky130_fd_sc_hs__nand2_1_9/A sky130_fd_sc_hs__o21a_1_11/a_320_74#
+ sky130_fd_sc_hs__o21a_1_11/a_376_387# sky130_fd_sc_hs__o21a_1_11/a_83_244# sky130_fd_sc_hs__o21a_1
Xsky130_fd_sc_hs__o21a_1_65 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__o21a_1_65/X sky130_fd_sc_hs__nor2_1_99/Y
+ sky130_fd_sc_hs__o21a_1_65/B1 sky130_fd_sc_hs__inv_4_101/A sky130_fd_sc_hs__o21a_1_65/a_320_74#
+ sky130_fd_sc_hs__o21a_1_65/a_376_387# sky130_fd_sc_hs__o21a_1_65/a_83_244# sky130_fd_sc_hs__o21a_1
Xsky130_fd_sc_hs__o21a_1_76 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__o21a_1_77/X sky130_fd_sc_hs__o21a_1_77/A2
+ sky130_fd_sc_hs__o21a_1_77/B1 sky130_fd_sc_hs__inv_4_113/A sky130_fd_sc_hs__o21a_1_77/a_320_74#
+ sky130_fd_sc_hs__o21a_1_77/a_376_387# sky130_fd_sc_hs__o21a_1_77/a_83_244# sky130_fd_sc_hs__o21a_1
Xsky130_fd_sc_hs__o21a_1_54 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__o21a_1_55/X sky130_fd_sc_hs__nor2_1_75/Y
+ sky130_fd_sc_hs__nor2_1_99/B sky130_fd_sc_hs__inv_4_97/A sky130_fd_sc_hs__o21a_1_55/a_320_74#
+ sky130_fd_sc_hs__o21a_1_55/a_376_387# sky130_fd_sc_hs__o21a_1_55/a_83_244# sky130_fd_sc_hs__o21a_1
Xsky130_fd_sc_hs__o21a_1_43 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__o21a_1_43/X sky130_fd_sc_hs__nor2_1_43/Y
+ sky130_fd_sc_hs__nor2_1_41/B sky130_fd_sc_hs__inv_4_73/A sky130_fd_sc_hs__o21a_1_43/a_320_74#
+ sky130_fd_sc_hs__o21a_1_43/a_376_387# sky130_fd_sc_hs__o21a_1_43/a_83_244# sky130_fd_sc_hs__o21a_1
Xsky130_fd_sc_hs__dfrtp_4_44 DVSS DVDD sky130_fd_sc_hs__clkbuf_8_1/A DVDD DVSS sky130_fd_sc_hs__o21a_1_19/X
+ sky130_fd_sc_hs__nand2_1_47/B sky130_fd_sc_hs__o21a_1_19/A1 sky130_fd_sc_hs__dfrtp_4_45/a_37_78#
+ sky130_fd_sc_hs__dfrtp_4_45/a_494_366# sky130_fd_sc_hs__dfrtp_4_45/a_699_463# sky130_fd_sc_hs__dfrtp_4_45/a_313_74#
+ sky130_fd_sc_hs__dfrtp_4_45/a_1627_493# sky130_fd_sc_hs__dfrtp_4_45/a_1678_395#
+ sky130_fd_sc_hs__dfrtp_4_45/a_1827_81# sky130_fd_sc_hs__dfrtp_4_45/a_789_463# sky130_fd_sc_hs__dfrtp_4_45/a_1350_392#
+ sky130_fd_sc_hs__dfrtp_4_45/a_834_355# sky130_fd_sc_hs__dfrtp_4_45/a_812_138# sky130_fd_sc_hs__dfrtp_4_45/a_124_78#
+ sky130_fd_sc_hs__dfrtp_4_45/a_1647_81# sky130_fd_sc_hs__dfrtp_4_45/a_2010_409# sky130_fd_sc_hs__dfrtp_4_45/a_890_138#
+ sky130_fd_sc_hs__dfrtp_4
Xsky130_fd_sc_hs__dfrtp_4_33 DVSS DVDD sky130_fd_sc_hs__clkbuf_8_1/X DVDD DVSS sky130_fd_sc_hs__a21oi_1_9/Y
+ sky130_fd_sc_hs__nand2_1_47/B sky130_fd_sc_hs__inv_4_11/A sky130_fd_sc_hs__dfrtp_4_33/a_37_78#
+ sky130_fd_sc_hs__dfrtp_4_33/a_494_366# sky130_fd_sc_hs__dfrtp_4_33/a_699_463# sky130_fd_sc_hs__dfrtp_4_33/a_313_74#
+ sky130_fd_sc_hs__dfrtp_4_33/a_1627_493# sky130_fd_sc_hs__dfrtp_4_33/a_1678_395#
+ sky130_fd_sc_hs__dfrtp_4_33/a_1827_81# sky130_fd_sc_hs__dfrtp_4_33/a_789_463# sky130_fd_sc_hs__dfrtp_4_33/a_1350_392#
+ sky130_fd_sc_hs__dfrtp_4_33/a_834_355# sky130_fd_sc_hs__dfrtp_4_33/a_812_138# sky130_fd_sc_hs__dfrtp_4_33/a_124_78#
+ sky130_fd_sc_hs__dfrtp_4_33/a_1647_81# sky130_fd_sc_hs__dfrtp_4_33/a_2010_409# sky130_fd_sc_hs__dfrtp_4_33/a_890_138#
+ sky130_fd_sc_hs__dfrtp_4
Xsky130_fd_sc_hs__dfrtp_4_22 DVSS DVDD sky130_fd_sc_hs__clkbuf_8_1/A DVDD DVSS sky130_fd_sc_hs__o21a_1_3/X
+ sky130_fd_sc_hs__nand2_1_47/B sky130_fd_sc_hs__o21a_1_3/A1 sky130_fd_sc_hs__dfrtp_4_23/a_37_78#
+ sky130_fd_sc_hs__dfrtp_4_23/a_494_366# sky130_fd_sc_hs__dfrtp_4_23/a_699_463# sky130_fd_sc_hs__dfrtp_4_23/a_313_74#
+ sky130_fd_sc_hs__dfrtp_4_23/a_1627_493# sky130_fd_sc_hs__dfrtp_4_23/a_1678_395#
+ sky130_fd_sc_hs__dfrtp_4_23/a_1827_81# sky130_fd_sc_hs__dfrtp_4_23/a_789_463# sky130_fd_sc_hs__dfrtp_4_23/a_1350_392#
+ sky130_fd_sc_hs__dfrtp_4_23/a_834_355# sky130_fd_sc_hs__dfrtp_4_23/a_812_138# sky130_fd_sc_hs__dfrtp_4_23/a_124_78#
+ sky130_fd_sc_hs__dfrtp_4_23/a_1647_81# sky130_fd_sc_hs__dfrtp_4_23/a_2010_409# sky130_fd_sc_hs__dfrtp_4_23/a_890_138#
+ sky130_fd_sc_hs__dfrtp_4
Xsky130_fd_sc_hs__dfrtp_4_11 DVSS DVDD sky130_fd_sc_hs__clkbuf_8_1/X DVDD DVSS sky130_fd_sc_hs__a21oi_1_1/Y
+ sky130_fd_sc_hs__nand2_1_47/B sky130_fd_sc_hs__inv_4_5/A sky130_fd_sc_hs__dfrtp_4_11/a_37_78#
+ sky130_fd_sc_hs__dfrtp_4_11/a_494_366# sky130_fd_sc_hs__dfrtp_4_11/a_699_463# sky130_fd_sc_hs__dfrtp_4_11/a_313_74#
+ sky130_fd_sc_hs__dfrtp_4_11/a_1627_493# sky130_fd_sc_hs__dfrtp_4_11/a_1678_395#
+ sky130_fd_sc_hs__dfrtp_4_11/a_1827_81# sky130_fd_sc_hs__dfrtp_4_11/a_789_463# sky130_fd_sc_hs__dfrtp_4_11/a_1350_392#
+ sky130_fd_sc_hs__dfrtp_4_11/a_834_355# sky130_fd_sc_hs__dfrtp_4_11/a_812_138# sky130_fd_sc_hs__dfrtp_4_11/a_124_78#
+ sky130_fd_sc_hs__dfrtp_4_11/a_1647_81# sky130_fd_sc_hs__dfrtp_4_11/a_2010_409# sky130_fd_sc_hs__dfrtp_4_11/a_890_138#
+ sky130_fd_sc_hs__dfrtp_4
Xsky130_fd_sc_hs__dfrtp_4_77 DVSS DVDD sky130_fd_sc_hs__clkbuf_8_1/A DVDD DVSS sky130_fd_sc_hs__dfrtp_4_77/D
+ sky130_fd_sc_hs__nand2_1_47/B sky130_fd_sc_hs__inv_4_35/A sky130_fd_sc_hs__dfrtp_4_77/a_37_78#
+ sky130_fd_sc_hs__dfrtp_4_77/a_494_366# sky130_fd_sc_hs__dfrtp_4_77/a_699_463# sky130_fd_sc_hs__dfrtp_4_77/a_313_74#
+ sky130_fd_sc_hs__dfrtp_4_77/a_1627_493# sky130_fd_sc_hs__dfrtp_4_77/a_1678_395#
+ sky130_fd_sc_hs__dfrtp_4_77/a_1827_81# sky130_fd_sc_hs__dfrtp_4_77/a_789_463# sky130_fd_sc_hs__dfrtp_4_77/a_1350_392#
+ sky130_fd_sc_hs__dfrtp_4_77/a_834_355# sky130_fd_sc_hs__dfrtp_4_77/a_812_138# sky130_fd_sc_hs__dfrtp_4_77/a_124_78#
+ sky130_fd_sc_hs__dfrtp_4_77/a_1647_81# sky130_fd_sc_hs__dfrtp_4_77/a_2010_409# sky130_fd_sc_hs__dfrtp_4_77/a_890_138#
+ sky130_fd_sc_hs__dfrtp_4
Xsky130_fd_sc_hs__dfrtp_4_66 DVSS DVDD sky130_fd_sc_hs__inv_4_49/Y DVDD DVSS sky130_fd_sc_hs__nor2b_1_15/Y
+ sky130_fd_sc_hs__dfstp_2_1/CLK sky130_fd_sc_hs__fa_2_15/B sky130_fd_sc_hs__dfrtp_4_67/a_37_78#
+ sky130_fd_sc_hs__dfrtp_4_67/a_494_366# sky130_fd_sc_hs__dfrtp_4_67/a_699_463# sky130_fd_sc_hs__dfrtp_4_67/a_313_74#
+ sky130_fd_sc_hs__dfrtp_4_67/a_1627_493# sky130_fd_sc_hs__dfrtp_4_67/a_1678_395#
+ sky130_fd_sc_hs__dfrtp_4_67/a_1827_81# sky130_fd_sc_hs__dfrtp_4_67/a_789_463# sky130_fd_sc_hs__dfrtp_4_67/a_1350_392#
+ sky130_fd_sc_hs__dfrtp_4_67/a_834_355# sky130_fd_sc_hs__dfrtp_4_67/a_812_138# sky130_fd_sc_hs__dfrtp_4_67/a_124_78#
+ sky130_fd_sc_hs__dfrtp_4_67/a_1647_81# sky130_fd_sc_hs__dfrtp_4_67/a_2010_409# sky130_fd_sc_hs__dfrtp_4_67/a_890_138#
+ sky130_fd_sc_hs__dfrtp_4
Xsky130_fd_sc_hs__dfrtp_4_55 DVSS DVDD sky130_fd_sc_hs__clkbuf_8_1/A DVDD DVSS sky130_fd_sc_hs__o21a_1_23/X
+ sky130_fd_sc_hs__nand2_1_47/B sky130_fd_sc_hs__o21a_1_23/A1 sky130_fd_sc_hs__dfrtp_4_55/a_37_78#
+ sky130_fd_sc_hs__dfrtp_4_55/a_494_366# sky130_fd_sc_hs__dfrtp_4_55/a_699_463# sky130_fd_sc_hs__dfrtp_4_55/a_313_74#
+ sky130_fd_sc_hs__dfrtp_4_55/a_1627_493# sky130_fd_sc_hs__dfrtp_4_55/a_1678_395#
+ sky130_fd_sc_hs__dfrtp_4_55/a_1827_81# sky130_fd_sc_hs__dfrtp_4_55/a_789_463# sky130_fd_sc_hs__dfrtp_4_55/a_1350_392#
+ sky130_fd_sc_hs__dfrtp_4_55/a_834_355# sky130_fd_sc_hs__dfrtp_4_55/a_812_138# sky130_fd_sc_hs__dfrtp_4_55/a_124_78#
+ sky130_fd_sc_hs__dfrtp_4_55/a_1647_81# sky130_fd_sc_hs__dfrtp_4_55/a_2010_409# sky130_fd_sc_hs__dfrtp_4_55/a_890_138#
+ sky130_fd_sc_hs__dfrtp_4
Xsky130_fd_sc_hs__dfrtp_4_88 DVSS DVDD sky130_fd_sc_hs__inv_4_49/Y DVDD DVSS ref_clk
+ clk_out sky130_fd_sc_hs__nand2_1_47/B sky130_fd_sc_hs__dfrtp_4_89/a_37_78# sky130_fd_sc_hs__dfrtp_4_89/a_494_366#
+ sky130_fd_sc_hs__dfrtp_4_89/a_699_463# sky130_fd_sc_hs__dfrtp_4_89/a_313_74# sky130_fd_sc_hs__dfrtp_4_89/a_1627_493#
+ sky130_fd_sc_hs__dfrtp_4_89/a_1678_395# sky130_fd_sc_hs__dfrtp_4_89/a_1827_81# sky130_fd_sc_hs__dfrtp_4_89/a_789_463#
+ sky130_fd_sc_hs__dfrtp_4_89/a_1350_392# sky130_fd_sc_hs__dfrtp_4_89/a_834_355# sky130_fd_sc_hs__dfrtp_4_89/a_812_138#
+ sky130_fd_sc_hs__dfrtp_4_89/a_124_78# sky130_fd_sc_hs__dfrtp_4_89/a_1647_81# sky130_fd_sc_hs__dfrtp_4_89/a_2010_409#
+ sky130_fd_sc_hs__dfrtp_4_89/a_890_138# sky130_fd_sc_hs__dfrtp_4
Xsky130_fd_sc_hs__nor2b_1_8 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__fa_2_11/SUM sky130_fd_sc_hs__nor2b_1_9/Y
+ sky130_fd_sc_hs__or2_1_1/A sky130_fd_sc_hs__nor2b_1_9/a_278_368# sky130_fd_sc_hs__nor2b_1_9/a_27_112#
+ sky130_fd_sc_hs__nor2b_1
Xsky130_fd_sc_hs__nand2_1_90 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_1_91/B sky130_fd_sc_hs__nand2_1_99/A
+ sky130_fd_sc_hs__nand2_1_91/A sky130_fd_sc_hs__nand2_1_91/a_117_74# sky130_fd_sc_hs__nand2_1
Xsky130_fd_sc_hs__nor2_1_6 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nor2_1_7/B sky130_fd_sc_hs__nor2_1_7/Y
+ sky130_fd_sc_hs__nor2_1_7/A sky130_fd_sc_hs__nor2_1_7/a_116_368# sky130_fd_sc_hs__nor2_1
Xsky130_fd_sc_hs__a21oi_1_47 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nor2_1_37/Y sky130_fd_sc_hs__dfrtp_4_77/D
+ sky130_fd_sc_hs__nor2_1_37/B sky130_fd_sc_hs__inv_4_35/Y sky130_fd_sc_hs__a21oi_1_47/a_117_74#
+ sky130_fd_sc_hs__a21oi_1_47/a_29_368# sky130_fd_sc_hs__a21oi_1
Xsky130_fd_sc_hs__a21oi_1_36 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__a222o_1_1/X sky130_fd_sc_hs__o31ai_1_1/A3
+ sky130_fd_sc_hs__nor2_1_33/Y sky130_fd_sc_hs__inv_4_35/A sky130_fd_sc_hs__a21oi_1_37/a_117_74#
+ sky130_fd_sc_hs__a21oi_1_37/a_29_368# sky130_fd_sc_hs__a21oi_1
Xsky130_fd_sc_hs__a21oi_1_25 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__a21oi_1_15/Y sky130_fd_sc_hs__a32oi_1_3/B1
+ sky130_fd_sc_hs__a211oi_1_1/Y sky130_fd_sc_hs__a22oi_1_15/Y sky130_fd_sc_hs__a21oi_1_25/a_117_74#
+ sky130_fd_sc_hs__a21oi_1_25/a_29_368# sky130_fd_sc_hs__a21oi_1
Xsky130_fd_sc_hs__a21oi_1_14 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_2_3/Y sky130_fd_sc_hs__a21oi_1_15/Y
+ sky130_fd_sc_hs__nor2_1_33/Y sky130_fd_sc_hs__o21a_1_3/A1 sky130_fd_sc_hs__a21oi_1_15/a_117_74#
+ sky130_fd_sc_hs__a21oi_1_15/a_29_368# sky130_fd_sc_hs__a21oi_1
Xsky130_fd_sc_hs__a21oi_1_69 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nor2_1_57/Y sky130_fd_sc_hs__dfrbp_1_11/D
+ sky130_fd_sc_hs__nor2_1_57/B sky130_fd_sc_hs__inv_4_79/Y sky130_fd_sc_hs__a21oi_1_69/a_117_74#
+ sky130_fd_sc_hs__a21oi_1_69/a_29_368# sky130_fd_sc_hs__a21oi_1
Xsky130_fd_sc_hs__a21oi_1_58 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nor2_1_45/Y sky130_fd_sc_hs__dfrtn_1_17/D
+ sky130_fd_sc_hs__nor2_1_45/B sky130_fd_sc_hs__inv_4_63/Y sky130_fd_sc_hs__a21oi_1_59/a_117_74#
+ sky130_fd_sc_hs__a21oi_1_59/a_29_368# sky130_fd_sc_hs__a21oi_1
Xsky130_fd_sc_hs__clkbuf_8_1 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__clkbuf_8_1/X sky130_fd_sc_hs__clkbuf_8_1/A
+ sky130_fd_sc_hs__clkbuf_8_1/a_125_368# sky130_fd_sc_hs__clkbuf_8
Xsky130_fd_sc_hs__nor3_1_10 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__xnor2_1_7/B sky130_fd_sc_hs__xnor2_1_3/B
+ sky130_fd_sc_hs__nor3_1_11/B sky130_fd_sc_hs__xnor2_1_3/A sky130_fd_sc_hs__nor3_1_11/a_198_368#
+ sky130_fd_sc_hs__nor3_1_11/a_114_368# sky130_fd_sc_hs__nor3_1
Xsky130_fd_sc_hs__o21a_1_7 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__o21a_1_7/X sky130_fd_sc_hs__o21a_1_7/A2
+ sky130_fd_sc_hs__nor2_1_5/B sky130_fd_sc_hs__o21a_1_7/A1 sky130_fd_sc_hs__o21a_1_7/a_320_74#
+ sky130_fd_sc_hs__o21a_1_7/a_376_387# sky130_fd_sc_hs__o21a_1_7/a_83_244# sky130_fd_sc_hs__o21a_1
Xsky130_fd_sc_hs__nor2_1_110 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__o21a_1_65/B1 sky130_fd_sc_hs__o21a_1_71/A2
+ sky130_fd_sc_hs__inv_4_99/Y sky130_fd_sc_hs__nor2_1_111/a_116_368# sky130_fd_sc_hs__nor2_1
Xsky130_fd_sc_hs__nor2_1_121 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__o21a_1_75/B1 sky130_fd_sc_hs__o21a_1_61/A2
+ sky130_fd_sc_hs__inv_4_135/Y sky130_fd_sc_hs__nor2_1_121/a_116_368# sky130_fd_sc_hs__nor2_1
Xsky130_fd_sc_hs__fa_2_15 DVSS DVDD sky130_fd_sc_hs__fa_2_9/B DVDD DVSS sky130_fd_sc_hs__fa_2_15/CIN
+ sky130_fd_sc_hs__fa_2_15/B sky130_fd_sc_hs__xor2_1_11/B sky130_fd_sc_hs__fa_2_15/SUM
+ sky130_fd_sc_hs__fa_2_15/a_27_378# sky130_fd_sc_hs__fa_2_15/a_701_79# sky130_fd_sc_hs__fa_2_15/a_484_347#
+ sky130_fd_sc_hs__fa_2_15/a_1094_347# sky130_fd_sc_hs__fa_2_15/a_1205_79# sky130_fd_sc_hs__fa_2_15/a_27_79#
+ sky130_fd_sc_hs__fa_2_15/a_1202_368# sky130_fd_sc_hs__fa_2_15/a_336_347# sky130_fd_sc_hs__fa_2_15/a_992_347#
+ sky130_fd_sc_hs__fa_2_15/a_1119_79# sky130_fd_sc_hs__fa_2_15/a_487_79# sky130_fd_sc_hs__fa_2_15/a_683_347#
+ sky130_fd_sc_hs__fa_2
Xsky130_fd_sc_hs__o21a_1_33 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__o21a_1_33/X sky130_fd_sc_hs__nor2_1_27/Y
+ sky130_fd_sc_hs__nor2_1_49/B sky130_fd_sc_hs__inv_4_55/A sky130_fd_sc_hs__o21a_1_33/a_320_74#
+ sky130_fd_sc_hs__o21a_1_33/a_376_387# sky130_fd_sc_hs__o21a_1_33/a_83_244# sky130_fd_sc_hs__o21a_1
Xsky130_fd_sc_hs__o21a_1_22 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__o21a_1_23/X sky130_fd_sc_hs__nor2_1_17/Y
+ sky130_fd_sc_hs__xnor2_1_1/B sky130_fd_sc_hs__o21a_1_23/A1 sky130_fd_sc_hs__o21a_1_23/a_320_74#
+ sky130_fd_sc_hs__o21a_1_23/a_376_387# sky130_fd_sc_hs__o21a_1_23/a_83_244# sky130_fd_sc_hs__o21a_1
Xsky130_fd_sc_hs__o21a_1_11 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__o21a_1_11/X sky130_fd_sc_hs__nor2_1_15/Y
+ sky130_fd_sc_hs__nor2_1_13/B sky130_fd_sc_hs__nand2_1_9/A sky130_fd_sc_hs__o21a_1_11/a_320_74#
+ sky130_fd_sc_hs__o21a_1_11/a_376_387# sky130_fd_sc_hs__o21a_1_11/a_83_244# sky130_fd_sc_hs__o21a_1
Xsky130_fd_sc_hs__o21a_1_66 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__o21a_1_67/X sky130_fd_sc_hs__o21a_1_67/A2
+ sky130_fd_sc_hs__o21a_1_67/B1 sky130_fd_sc_hs__inv_4_133/A sky130_fd_sc_hs__o21a_1_67/a_320_74#
+ sky130_fd_sc_hs__o21a_1_67/a_376_387# sky130_fd_sc_hs__o21a_1_67/a_83_244# sky130_fd_sc_hs__o21a_1
Xsky130_fd_sc_hs__o21a_1_55 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__o21a_1_55/X sky130_fd_sc_hs__nor2_1_75/Y
+ sky130_fd_sc_hs__nor2_1_99/B sky130_fd_sc_hs__inv_4_97/A sky130_fd_sc_hs__o21a_1_55/a_320_74#
+ sky130_fd_sc_hs__o21a_1_55/a_376_387# sky130_fd_sc_hs__o21a_1_55/a_83_244# sky130_fd_sc_hs__o21a_1
Xsky130_fd_sc_hs__o21a_1_44 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__o21a_1_45/X sky130_fd_sc_hs__nor2_1_57/Y
+ sky130_fd_sc_hs__nor2_1_83/B sky130_fd_sc_hs__inv_4_69/A sky130_fd_sc_hs__o21a_1_45/a_320_74#
+ sky130_fd_sc_hs__o21a_1_45/a_376_387# sky130_fd_sc_hs__o21a_1_45/a_83_244# sky130_fd_sc_hs__o21a_1
Xsky130_fd_sc_hs__o21a_1_77 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__o21a_1_77/X sky130_fd_sc_hs__o21a_1_77/A2
+ sky130_fd_sc_hs__o21a_1_77/B1 sky130_fd_sc_hs__inv_4_113/A sky130_fd_sc_hs__o21a_1_77/a_320_74#
+ sky130_fd_sc_hs__o21a_1_77/a_376_387# sky130_fd_sc_hs__o21a_1_77/a_83_244# sky130_fd_sc_hs__o21a_1
Xsky130_fd_sc_hs__dfrtp_4_34 DVSS DVDD sky130_fd_sc_hs__clkbuf_8_1/A DVDD DVSS sky130_fd_sc_hs__dfrtp_4_35/D
+ sky130_fd_sc_hs__nand2_1_47/B sky130_fd_sc_hs__inv_4_15/A sky130_fd_sc_hs__dfrtp_4_35/a_37_78#
+ sky130_fd_sc_hs__dfrtp_4_35/a_494_366# sky130_fd_sc_hs__dfrtp_4_35/a_699_463# sky130_fd_sc_hs__dfrtp_4_35/a_313_74#
+ sky130_fd_sc_hs__dfrtp_4_35/a_1627_493# sky130_fd_sc_hs__dfrtp_4_35/a_1678_395#
+ sky130_fd_sc_hs__dfrtp_4_35/a_1827_81# sky130_fd_sc_hs__dfrtp_4_35/a_789_463# sky130_fd_sc_hs__dfrtp_4_35/a_1350_392#
+ sky130_fd_sc_hs__dfrtp_4_35/a_834_355# sky130_fd_sc_hs__dfrtp_4_35/a_812_138# sky130_fd_sc_hs__dfrtp_4_35/a_124_78#
+ sky130_fd_sc_hs__dfrtp_4_35/a_1647_81# sky130_fd_sc_hs__dfrtp_4_35/a_2010_409# sky130_fd_sc_hs__dfrtp_4_35/a_890_138#
+ sky130_fd_sc_hs__dfrtp_4
Xsky130_fd_sc_hs__dfrtp_4_23 DVSS DVDD sky130_fd_sc_hs__clkbuf_8_1/A DVDD DVSS sky130_fd_sc_hs__o21a_1_3/X
+ sky130_fd_sc_hs__nand2_1_47/B sky130_fd_sc_hs__o21a_1_3/A1 sky130_fd_sc_hs__dfrtp_4_23/a_37_78#
+ sky130_fd_sc_hs__dfrtp_4_23/a_494_366# sky130_fd_sc_hs__dfrtp_4_23/a_699_463# sky130_fd_sc_hs__dfrtp_4_23/a_313_74#
+ sky130_fd_sc_hs__dfrtp_4_23/a_1627_493# sky130_fd_sc_hs__dfrtp_4_23/a_1678_395#
+ sky130_fd_sc_hs__dfrtp_4_23/a_1827_81# sky130_fd_sc_hs__dfrtp_4_23/a_789_463# sky130_fd_sc_hs__dfrtp_4_23/a_1350_392#
+ sky130_fd_sc_hs__dfrtp_4_23/a_834_355# sky130_fd_sc_hs__dfrtp_4_23/a_812_138# sky130_fd_sc_hs__dfrtp_4_23/a_124_78#
+ sky130_fd_sc_hs__dfrtp_4_23/a_1647_81# sky130_fd_sc_hs__dfrtp_4_23/a_2010_409# sky130_fd_sc_hs__dfrtp_4_23/a_890_138#
+ sky130_fd_sc_hs__dfrtp_4
Xsky130_fd_sc_hs__dfrtp_4_12 DVSS DVDD sky130_fd_sc_hs__clkbuf_8_1/A DVDD DVSS sky130_fd_sc_hs__o21a_1_5/X
+ sky130_fd_sc_hs__nand2_1_47/B sky130_fd_sc_hs__o21a_1_5/A1 sky130_fd_sc_hs__dfrtp_4_13/a_37_78#
+ sky130_fd_sc_hs__dfrtp_4_13/a_494_366# sky130_fd_sc_hs__dfrtp_4_13/a_699_463# sky130_fd_sc_hs__dfrtp_4_13/a_313_74#
+ sky130_fd_sc_hs__dfrtp_4_13/a_1627_493# sky130_fd_sc_hs__dfrtp_4_13/a_1678_395#
+ sky130_fd_sc_hs__dfrtp_4_13/a_1827_81# sky130_fd_sc_hs__dfrtp_4_13/a_789_463# sky130_fd_sc_hs__dfrtp_4_13/a_1350_392#
+ sky130_fd_sc_hs__dfrtp_4_13/a_834_355# sky130_fd_sc_hs__dfrtp_4_13/a_812_138# sky130_fd_sc_hs__dfrtp_4_13/a_124_78#
+ sky130_fd_sc_hs__dfrtp_4_13/a_1647_81# sky130_fd_sc_hs__dfrtp_4_13/a_2010_409# sky130_fd_sc_hs__dfrtp_4_13/a_890_138#
+ sky130_fd_sc_hs__dfrtp_4
Xsky130_fd_sc_hs__dfrtp_4_67 DVSS DVDD sky130_fd_sc_hs__inv_4_49/Y DVDD DVSS sky130_fd_sc_hs__nor2b_1_15/Y
+ sky130_fd_sc_hs__dfstp_2_1/CLK sky130_fd_sc_hs__fa_2_15/B sky130_fd_sc_hs__dfrtp_4_67/a_37_78#
+ sky130_fd_sc_hs__dfrtp_4_67/a_494_366# sky130_fd_sc_hs__dfrtp_4_67/a_699_463# sky130_fd_sc_hs__dfrtp_4_67/a_313_74#
+ sky130_fd_sc_hs__dfrtp_4_67/a_1627_493# sky130_fd_sc_hs__dfrtp_4_67/a_1678_395#
+ sky130_fd_sc_hs__dfrtp_4_67/a_1827_81# sky130_fd_sc_hs__dfrtp_4_67/a_789_463# sky130_fd_sc_hs__dfrtp_4_67/a_1350_392#
+ sky130_fd_sc_hs__dfrtp_4_67/a_834_355# sky130_fd_sc_hs__dfrtp_4_67/a_812_138# sky130_fd_sc_hs__dfrtp_4_67/a_124_78#
+ sky130_fd_sc_hs__dfrtp_4_67/a_1647_81# sky130_fd_sc_hs__dfrtp_4_67/a_2010_409# sky130_fd_sc_hs__dfrtp_4_67/a_890_138#
+ sky130_fd_sc_hs__dfrtp_4
Xsky130_fd_sc_hs__dfrtp_4_56 DVSS DVDD sky130_fd_sc_hs__clkbuf_8_1/X DVDD DVSS sky130_fd_sc_hs__dfrtp_4_57/D
+ sky130_fd_sc_hs__nand2_1_47/B sky130_fd_sc_hs__inv_4_29/A sky130_fd_sc_hs__dfrtp_4_57/a_37_78#
+ sky130_fd_sc_hs__dfrtp_4_57/a_494_366# sky130_fd_sc_hs__dfrtp_4_57/a_699_463# sky130_fd_sc_hs__dfrtp_4_57/a_313_74#
+ sky130_fd_sc_hs__dfrtp_4_57/a_1627_493# sky130_fd_sc_hs__dfrtp_4_57/a_1678_395#
+ sky130_fd_sc_hs__dfrtp_4_57/a_1827_81# sky130_fd_sc_hs__dfrtp_4_57/a_789_463# sky130_fd_sc_hs__dfrtp_4_57/a_1350_392#
+ sky130_fd_sc_hs__dfrtp_4_57/a_834_355# sky130_fd_sc_hs__dfrtp_4_57/a_812_138# sky130_fd_sc_hs__dfrtp_4_57/a_124_78#
+ sky130_fd_sc_hs__dfrtp_4_57/a_1647_81# sky130_fd_sc_hs__dfrtp_4_57/a_2010_409# sky130_fd_sc_hs__dfrtp_4_57/a_890_138#
+ sky130_fd_sc_hs__dfrtp_4
Xsky130_fd_sc_hs__dfrtp_4_45 DVSS DVDD sky130_fd_sc_hs__clkbuf_8_1/A DVDD DVSS sky130_fd_sc_hs__o21a_1_19/X
+ sky130_fd_sc_hs__nand2_1_47/B sky130_fd_sc_hs__o21a_1_19/A1 sky130_fd_sc_hs__dfrtp_4_45/a_37_78#
+ sky130_fd_sc_hs__dfrtp_4_45/a_494_366# sky130_fd_sc_hs__dfrtp_4_45/a_699_463# sky130_fd_sc_hs__dfrtp_4_45/a_313_74#
+ sky130_fd_sc_hs__dfrtp_4_45/a_1627_493# sky130_fd_sc_hs__dfrtp_4_45/a_1678_395#
+ sky130_fd_sc_hs__dfrtp_4_45/a_1827_81# sky130_fd_sc_hs__dfrtp_4_45/a_789_463# sky130_fd_sc_hs__dfrtp_4_45/a_1350_392#
+ sky130_fd_sc_hs__dfrtp_4_45/a_834_355# sky130_fd_sc_hs__dfrtp_4_45/a_812_138# sky130_fd_sc_hs__dfrtp_4_45/a_124_78#
+ sky130_fd_sc_hs__dfrtp_4_45/a_1647_81# sky130_fd_sc_hs__dfrtp_4_45/a_2010_409# sky130_fd_sc_hs__dfrtp_4_45/a_890_138#
+ sky130_fd_sc_hs__dfrtp_4
Xsky130_fd_sc_hs__dfrtp_4_89 DVSS DVDD sky130_fd_sc_hs__inv_4_49/Y DVDD DVSS ref_clk
+ clk_out sky130_fd_sc_hs__nand2_1_47/B sky130_fd_sc_hs__dfrtp_4_89/a_37_78# sky130_fd_sc_hs__dfrtp_4_89/a_494_366#
+ sky130_fd_sc_hs__dfrtp_4_89/a_699_463# sky130_fd_sc_hs__dfrtp_4_89/a_313_74# sky130_fd_sc_hs__dfrtp_4_89/a_1627_493#
+ sky130_fd_sc_hs__dfrtp_4_89/a_1678_395# sky130_fd_sc_hs__dfrtp_4_89/a_1827_81# sky130_fd_sc_hs__dfrtp_4_89/a_789_463#
+ sky130_fd_sc_hs__dfrtp_4_89/a_1350_392# sky130_fd_sc_hs__dfrtp_4_89/a_834_355# sky130_fd_sc_hs__dfrtp_4_89/a_812_138#
+ sky130_fd_sc_hs__dfrtp_4_89/a_124_78# sky130_fd_sc_hs__dfrtp_4_89/a_1647_81# sky130_fd_sc_hs__dfrtp_4_89/a_2010_409#
+ sky130_fd_sc_hs__dfrtp_4_89/a_890_138# sky130_fd_sc_hs__dfrtp_4
Xsky130_fd_sc_hs__dfrtp_4_78 DVSS DVDD sky130_fd_sc_hs__clkbuf_8_1/X DVDD DVSS sky130_fd_sc_hs__dfrtp_4_79/D
+ sky130_fd_sc_hs__nand2_1_47/B sky130_fd_sc_hs__inv_4_41/A sky130_fd_sc_hs__dfrtp_4_79/a_37_78#
+ sky130_fd_sc_hs__dfrtp_4_79/a_494_366# sky130_fd_sc_hs__dfrtp_4_79/a_699_463# sky130_fd_sc_hs__dfrtp_4_79/a_313_74#
+ sky130_fd_sc_hs__dfrtp_4_79/a_1627_493# sky130_fd_sc_hs__dfrtp_4_79/a_1678_395#
+ sky130_fd_sc_hs__dfrtp_4_79/a_1827_81# sky130_fd_sc_hs__dfrtp_4_79/a_789_463# sky130_fd_sc_hs__dfrtp_4_79/a_1350_392#
+ sky130_fd_sc_hs__dfrtp_4_79/a_834_355# sky130_fd_sc_hs__dfrtp_4_79/a_812_138# sky130_fd_sc_hs__dfrtp_4_79/a_124_78#
+ sky130_fd_sc_hs__dfrtp_4_79/a_1647_81# sky130_fd_sc_hs__dfrtp_4_79/a_2010_409# sky130_fd_sc_hs__dfrtp_4_79/a_890_138#
+ sky130_fd_sc_hs__dfrtp_4
Xsky130_fd_sc_hs__nor2b_1_9 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__fa_2_11/SUM sky130_fd_sc_hs__nor2b_1_9/Y
+ sky130_fd_sc_hs__or2_1_1/A sky130_fd_sc_hs__nor2b_1_9/a_278_368# sky130_fd_sc_hs__nor2b_1_9/a_27_112#
+ sky130_fd_sc_hs__nor2b_1
Xsky130_fd_sc_hs__nand2_1_91 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_1_91/B sky130_fd_sc_hs__nand2_1_99/A
+ sky130_fd_sc_hs__nand2_1_91/A sky130_fd_sc_hs__nand2_1_91/a_117_74# sky130_fd_sc_hs__nand2_1
Xsky130_fd_sc_hs__nand2_1_80 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_2_3/A sky130_fd_sc_hs__nand2_1_91/A
+ sky130_fd_sc_hs__inv_2_5/Y sky130_fd_sc_hs__nand2_1_81/a_117_74# sky130_fd_sc_hs__nand2_1
Xsky130_fd_sc_hs__nor2_1_7 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nor2_1_7/B sky130_fd_sc_hs__nor2_1_7/Y
+ sky130_fd_sc_hs__nor2_1_7/A sky130_fd_sc_hs__nor2_1_7/a_116_368# sky130_fd_sc_hs__nor2_1
Xsky130_fd_sc_hs__a21oi_1_37 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__a222o_1_1/X sky130_fd_sc_hs__o31ai_1_1/A3
+ sky130_fd_sc_hs__nor2_1_33/Y sky130_fd_sc_hs__inv_4_35/A sky130_fd_sc_hs__a21oi_1_37/a_117_74#
+ sky130_fd_sc_hs__a21oi_1_37/a_29_368# sky130_fd_sc_hs__a21oi_1
Xsky130_fd_sc_hs__a21oi_1_26 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__a21oi_1_17/Y sky130_fd_sc_hs__o31ai_1_1/B1
+ sky130_fd_sc_hs__a21oi_1_19/Y fine_control_avg_window_select[1] sky130_fd_sc_hs__a21oi_1_27/a_117_74#
+ sky130_fd_sc_hs__a21oi_1_27/a_29_368# sky130_fd_sc_hs__a21oi_1
Xsky130_fd_sc_hs__a21oi_1_15 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_2_3/Y sky130_fd_sc_hs__a21oi_1_15/Y
+ sky130_fd_sc_hs__nor2_1_33/Y sky130_fd_sc_hs__o21a_1_3/A1 sky130_fd_sc_hs__a21oi_1_15/a_117_74#
+ sky130_fd_sc_hs__a21oi_1_15/a_29_368# sky130_fd_sc_hs__a21oi_1
Xsky130_fd_sc_hs__a21oi_1_59 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nor2_1_45/Y sky130_fd_sc_hs__dfrtn_1_17/D
+ sky130_fd_sc_hs__nor2_1_45/B sky130_fd_sc_hs__inv_4_63/Y sky130_fd_sc_hs__a21oi_1_59/a_117_74#
+ sky130_fd_sc_hs__a21oi_1_59/a_29_368# sky130_fd_sc_hs__a21oi_1
Xsky130_fd_sc_hs__a21oi_1_48 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nor2_1_27/Y sky130_fd_sc_hs__dfrtn_1_3/D
+ sky130_fd_sc_hs__nor2_1_27/B sky130_fd_sc_hs__inv_4_37/Y sky130_fd_sc_hs__a21oi_1_49/a_117_74#
+ sky130_fd_sc_hs__a21oi_1_49/a_29_368# sky130_fd_sc_hs__a21oi_1
Xsky130_fd_sc_hs__nor3_1_11 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__xnor2_1_7/B sky130_fd_sc_hs__xnor2_1_3/B
+ sky130_fd_sc_hs__nor3_1_11/B sky130_fd_sc_hs__xnor2_1_3/A sky130_fd_sc_hs__nor3_1_11/a_198_368#
+ sky130_fd_sc_hs__nor3_1_11/a_114_368# sky130_fd_sc_hs__nor3_1
Xsky130_fd_sc_hs__o21a_1_8 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__o21a_1_9/X sky130_fd_sc_hs__nor2_1_9/Y
+ sky130_fd_sc_hs__o21a_1_9/B1 sky130_fd_sc_hs__o21a_1_9/A1 sky130_fd_sc_hs__o21a_1_9/a_320_74#
+ sky130_fd_sc_hs__o21a_1_9/a_376_387# sky130_fd_sc_hs__o21a_1_9/a_83_244# sky130_fd_sc_hs__o21a_1
Xsky130_fd_sc_hs__nor2_1_100 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_121/Y sky130_fd_sc_hs__nor2_1_101/Y
+ sky130_fd_sc_hs__o21ai_1_7/Y sky130_fd_sc_hs__nor2_1_101/a_116_368# sky130_fd_sc_hs__nor2_1
Xsky130_fd_sc_hs__nor2_1_111 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__o21a_1_65/B1 sky130_fd_sc_hs__o21a_1_71/A2
+ sky130_fd_sc_hs__inv_4_99/Y sky130_fd_sc_hs__nor2_1_111/a_116_368# sky130_fd_sc_hs__nor2_1
Xsky130_fd_sc_hs__nor2_1_122 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__o21a_1_77/B1 sky130_fd_sc_hs__o21a_1_63/A2
+ sky130_fd_sc_hs__inv_4_137/Y sky130_fd_sc_hs__nor2_1_123/a_116_368# sky130_fd_sc_hs__nor2_1
Xsky130_fd_sc_hs__a22oi_1_20 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_33/Y sky130_fd_sc_hs__a22oi_1_21/Y
+ sky130_fd_sc_hs__a32oi_1_5/A1 sky130_fd_sc_hs__a222oi_1_1/Y fine_control_avg_window_select[0]
+ sky130_fd_sc_hs__a22oi_1_21/a_71_368# sky130_fd_sc_hs__a22oi_1_21/a_159_74# sky130_fd_sc_hs__a22oi_1_21/a_339_74#
+ sky130_fd_sc_hs__a22oi_1
Xsky130_fd_sc_hs__fa_2_16 DVSS DVDD sky130_fd_sc_hs__fa_2_9/B DVDD DVSS sky130_fd_sc_hs__fa_2_17/CIN
+ sky130_fd_sc_hs__fa_2_17/B sky130_fd_sc_hs__fa_2_19/CIN sky130_fd_sc_hs__fa_2_17/SUM
+ sky130_fd_sc_hs__fa_2_17/a_27_378# sky130_fd_sc_hs__fa_2_17/a_701_79# sky130_fd_sc_hs__fa_2_17/a_484_347#
+ sky130_fd_sc_hs__fa_2_17/a_1094_347# sky130_fd_sc_hs__fa_2_17/a_1205_79# sky130_fd_sc_hs__fa_2_17/a_27_79#
+ sky130_fd_sc_hs__fa_2_17/a_1202_368# sky130_fd_sc_hs__fa_2_17/a_336_347# sky130_fd_sc_hs__fa_2_17/a_992_347#
+ sky130_fd_sc_hs__fa_2_17/a_1119_79# sky130_fd_sc_hs__fa_2_17/a_487_79# sky130_fd_sc_hs__fa_2_17/a_683_347#
+ sky130_fd_sc_hs__fa_2
Xsky130_fd_sc_hs__dfsbp_2_0 DVSS DVDD sky130_fd_sc_hs__inv_4_49/Y DVDD DVSS sky130_fd_sc_hs__o21ai_1_1/Y
+ sky130_fd_sc_hs__dfstp_2_7/Q sky130_fd_sc_hs__inv_4_23/A sky130_fd_sc_hs__dfsbp_2_1/Q
+ sky130_fd_sc_hs__dfsbp_2_1/a_595_97# sky130_fd_sc_hs__dfsbp_2_1/a_731_97# sky130_fd_sc_hs__dfsbp_2_1/a_1521_508#
+ sky130_fd_sc_hs__dfsbp_2_1/a_2221_74# sky130_fd_sc_hs__dfsbp_2_1/a_1339_74# sky130_fd_sc_hs__dfsbp_2_1/a_1531_118#
+ sky130_fd_sc_hs__dfsbp_2_1/a_1453_118# sky130_fd_sc_hs__dfsbp_2_1/a_398_74# sky130_fd_sc_hs__dfsbp_2_1/a_27_74#
+ sky130_fd_sc_hs__dfsbp_2_1/a_225_74# sky130_fd_sc_hs__dfsbp_2_1/a_1501_92# sky130_fd_sc_hs__dfsbp_2_1/a_757_401#
+ sky130_fd_sc_hs__dfsbp_2_1/a_1258_341# sky130_fd_sc_hs__dfsbp_2_1/a_1001_74# sky130_fd_sc_hs__dfsbp_2_1/a_706_463#
+ sky130_fd_sc_hs__dfsbp_2_1/a_1261_74# sky130_fd_sc_hs__dfsbp_2
Xsky130_fd_sc_hs__nand2b_4_0 DVSS DVDD DVDD DVSS div_ratio_half[4] sky130_fd_sc_hs__xnor2_1_13/A
+ sky130_fd_sc_hs__inv_4_103/A sky130_fd_sc_hs__nand2b_4_1/a_31_74# sky130_fd_sc_hs__nand2b_4_1/a_243_74#
+ sky130_fd_sc_hs__nand2b_4
Xsky130_fd_sc_hs__o21a_1_23 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__o21a_1_23/X sky130_fd_sc_hs__nor2_1_17/Y
+ sky130_fd_sc_hs__xnor2_1_1/B sky130_fd_sc_hs__o21a_1_23/A1 sky130_fd_sc_hs__o21a_1_23/a_320_74#
+ sky130_fd_sc_hs__o21a_1_23/a_376_387# sky130_fd_sc_hs__o21a_1_23/a_83_244# sky130_fd_sc_hs__o21a_1
Xsky130_fd_sc_hs__o21a_1_12 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__o21a_1_13/X sky130_fd_sc_hs__nor2_1_11/Y
+ sky130_fd_sc_hs__nor2_1_31/B sky130_fd_sc_hs__o21a_1_13/A1 sky130_fd_sc_hs__o21a_1_13/a_320_74#
+ sky130_fd_sc_hs__o21a_1_13/a_376_387# sky130_fd_sc_hs__o21a_1_13/a_83_244# sky130_fd_sc_hs__o21a_1
Xsky130_fd_sc_hs__o21a_1_67 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__o21a_1_67/X sky130_fd_sc_hs__o21a_1_67/A2
+ sky130_fd_sc_hs__o21a_1_67/B1 sky130_fd_sc_hs__inv_4_133/A sky130_fd_sc_hs__o21a_1_67/a_320_74#
+ sky130_fd_sc_hs__o21a_1_67/a_376_387# sky130_fd_sc_hs__o21a_1_67/a_83_244# sky130_fd_sc_hs__o21a_1
Xsky130_fd_sc_hs__o21a_1_56 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__o21a_1_57/X sky130_fd_sc_hs__nor2_1_47/Y
+ sky130_fd_sc_hs__o21a_1_57/B1 sky130_fd_sc_hs__inv_4_93/A sky130_fd_sc_hs__o21a_1_57/a_320_74#
+ sky130_fd_sc_hs__o21a_1_57/a_376_387# sky130_fd_sc_hs__o21a_1_57/a_83_244# sky130_fd_sc_hs__o21a_1
Xsky130_fd_sc_hs__o21a_1_45 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__o21a_1_45/X sky130_fd_sc_hs__nor2_1_57/Y
+ sky130_fd_sc_hs__nor2_1_83/B sky130_fd_sc_hs__inv_4_69/A sky130_fd_sc_hs__o21a_1_45/a_320_74#
+ sky130_fd_sc_hs__o21a_1_45/a_376_387# sky130_fd_sc_hs__o21a_1_45/a_83_244# sky130_fd_sc_hs__o21a_1
Xsky130_fd_sc_hs__o21a_1_34 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__o21a_1_35/X sky130_fd_sc_hs__nor2_1_41/Y
+ sky130_fd_sc_hs__nor2_1_51/B sky130_fd_sc_hs__dfrbp_1_1/Q sky130_fd_sc_hs__o21a_1_35/a_320_74#
+ sky130_fd_sc_hs__o21a_1_35/a_376_387# sky130_fd_sc_hs__o21a_1_35/a_83_244# sky130_fd_sc_hs__o21a_1
Xsky130_fd_sc_hs__dfrtp_4_24 DVSS DVDD sky130_fd_sc_hs__clkbuf_8_1/X DVDD DVSS sky130_fd_sc_hs__dfrtp_4_25/D
+ sky130_fd_sc_hs__nand2_1_47/B sky130_fd_sc_hs__inv_4_13/A sky130_fd_sc_hs__dfrtp_4_25/a_37_78#
+ sky130_fd_sc_hs__dfrtp_4_25/a_494_366# sky130_fd_sc_hs__dfrtp_4_25/a_699_463# sky130_fd_sc_hs__dfrtp_4_25/a_313_74#
+ sky130_fd_sc_hs__dfrtp_4_25/a_1627_493# sky130_fd_sc_hs__dfrtp_4_25/a_1678_395#
+ sky130_fd_sc_hs__dfrtp_4_25/a_1827_81# sky130_fd_sc_hs__dfrtp_4_25/a_789_463# sky130_fd_sc_hs__dfrtp_4_25/a_1350_392#
+ sky130_fd_sc_hs__dfrtp_4_25/a_834_355# sky130_fd_sc_hs__dfrtp_4_25/a_812_138# sky130_fd_sc_hs__dfrtp_4_25/a_124_78#
+ sky130_fd_sc_hs__dfrtp_4_25/a_1647_81# sky130_fd_sc_hs__dfrtp_4_25/a_2010_409# sky130_fd_sc_hs__dfrtp_4_25/a_890_138#
+ sky130_fd_sc_hs__dfrtp_4
Xsky130_fd_sc_hs__dfrtp_4_13 DVSS DVDD sky130_fd_sc_hs__clkbuf_8_1/A DVDD DVSS sky130_fd_sc_hs__o21a_1_5/X
+ sky130_fd_sc_hs__nand2_1_47/B sky130_fd_sc_hs__o21a_1_5/A1 sky130_fd_sc_hs__dfrtp_4_13/a_37_78#
+ sky130_fd_sc_hs__dfrtp_4_13/a_494_366# sky130_fd_sc_hs__dfrtp_4_13/a_699_463# sky130_fd_sc_hs__dfrtp_4_13/a_313_74#
+ sky130_fd_sc_hs__dfrtp_4_13/a_1627_493# sky130_fd_sc_hs__dfrtp_4_13/a_1678_395#
+ sky130_fd_sc_hs__dfrtp_4_13/a_1827_81# sky130_fd_sc_hs__dfrtp_4_13/a_789_463# sky130_fd_sc_hs__dfrtp_4_13/a_1350_392#
+ sky130_fd_sc_hs__dfrtp_4_13/a_834_355# sky130_fd_sc_hs__dfrtp_4_13/a_812_138# sky130_fd_sc_hs__dfrtp_4_13/a_124_78#
+ sky130_fd_sc_hs__dfrtp_4_13/a_1647_81# sky130_fd_sc_hs__dfrtp_4_13/a_2010_409# sky130_fd_sc_hs__dfrtp_4_13/a_890_138#
+ sky130_fd_sc_hs__dfrtp_4
Xsky130_fd_sc_hs__dfrtp_4_68 DVSS DVDD sky130_fd_sc_hs__clkbuf_8_1/A DVDD DVSS sky130_fd_sc_hs__xnor2_1_1/Y
+ sky130_fd_sc_hs__nand2_1_47/B sky130_fd_sc_hs__xnor2_1_1/A sky130_fd_sc_hs__dfrtp_4_69/a_37_78#
+ sky130_fd_sc_hs__dfrtp_4_69/a_494_366# sky130_fd_sc_hs__dfrtp_4_69/a_699_463# sky130_fd_sc_hs__dfrtp_4_69/a_313_74#
+ sky130_fd_sc_hs__dfrtp_4_69/a_1627_493# sky130_fd_sc_hs__dfrtp_4_69/a_1678_395#
+ sky130_fd_sc_hs__dfrtp_4_69/a_1827_81# sky130_fd_sc_hs__dfrtp_4_69/a_789_463# sky130_fd_sc_hs__dfrtp_4_69/a_1350_392#
+ sky130_fd_sc_hs__dfrtp_4_69/a_834_355# sky130_fd_sc_hs__dfrtp_4_69/a_812_138# sky130_fd_sc_hs__dfrtp_4_69/a_124_78#
+ sky130_fd_sc_hs__dfrtp_4_69/a_1647_81# sky130_fd_sc_hs__dfrtp_4_69/a_2010_409# sky130_fd_sc_hs__dfrtp_4_69/a_890_138#
+ sky130_fd_sc_hs__dfrtp_4
Xsky130_fd_sc_hs__dfrtp_4_57 DVSS DVDD sky130_fd_sc_hs__clkbuf_8_1/X DVDD DVSS sky130_fd_sc_hs__dfrtp_4_57/D
+ sky130_fd_sc_hs__nand2_1_47/B sky130_fd_sc_hs__inv_4_29/A sky130_fd_sc_hs__dfrtp_4_57/a_37_78#
+ sky130_fd_sc_hs__dfrtp_4_57/a_494_366# sky130_fd_sc_hs__dfrtp_4_57/a_699_463# sky130_fd_sc_hs__dfrtp_4_57/a_313_74#
+ sky130_fd_sc_hs__dfrtp_4_57/a_1627_493# sky130_fd_sc_hs__dfrtp_4_57/a_1678_395#
+ sky130_fd_sc_hs__dfrtp_4_57/a_1827_81# sky130_fd_sc_hs__dfrtp_4_57/a_789_463# sky130_fd_sc_hs__dfrtp_4_57/a_1350_392#
+ sky130_fd_sc_hs__dfrtp_4_57/a_834_355# sky130_fd_sc_hs__dfrtp_4_57/a_812_138# sky130_fd_sc_hs__dfrtp_4_57/a_124_78#
+ sky130_fd_sc_hs__dfrtp_4_57/a_1647_81# sky130_fd_sc_hs__dfrtp_4_57/a_2010_409# sky130_fd_sc_hs__dfrtp_4_57/a_890_138#
+ sky130_fd_sc_hs__dfrtp_4
Xsky130_fd_sc_hs__dfrtp_4_46 DVSS DVDD sky130_fd_sc_hs__inv_4_49/Y DVDD DVSS sky130_fd_sc_hs__nor2b_1_11/Y
+ sky130_fd_sc_hs__dfstp_2_1/CLK sky130_fd_sc_hs__fa_2_9/A sky130_fd_sc_hs__dfrtp_4_47/a_37_78#
+ sky130_fd_sc_hs__dfrtp_4_47/a_494_366# sky130_fd_sc_hs__dfrtp_4_47/a_699_463# sky130_fd_sc_hs__dfrtp_4_47/a_313_74#
+ sky130_fd_sc_hs__dfrtp_4_47/a_1627_493# sky130_fd_sc_hs__dfrtp_4_47/a_1678_395#
+ sky130_fd_sc_hs__dfrtp_4_47/a_1827_81# sky130_fd_sc_hs__dfrtp_4_47/a_789_463# sky130_fd_sc_hs__dfrtp_4_47/a_1350_392#
+ sky130_fd_sc_hs__dfrtp_4_47/a_834_355# sky130_fd_sc_hs__dfrtp_4_47/a_812_138# sky130_fd_sc_hs__dfrtp_4_47/a_124_78#
+ sky130_fd_sc_hs__dfrtp_4_47/a_1647_81# sky130_fd_sc_hs__dfrtp_4_47/a_2010_409# sky130_fd_sc_hs__dfrtp_4_47/a_890_138#
+ sky130_fd_sc_hs__dfrtp_4
Xsky130_fd_sc_hs__dfrtp_4_35 DVSS DVDD sky130_fd_sc_hs__clkbuf_8_1/A DVDD DVSS sky130_fd_sc_hs__dfrtp_4_35/D
+ sky130_fd_sc_hs__nand2_1_47/B sky130_fd_sc_hs__inv_4_15/A sky130_fd_sc_hs__dfrtp_4_35/a_37_78#
+ sky130_fd_sc_hs__dfrtp_4_35/a_494_366# sky130_fd_sc_hs__dfrtp_4_35/a_699_463# sky130_fd_sc_hs__dfrtp_4_35/a_313_74#
+ sky130_fd_sc_hs__dfrtp_4_35/a_1627_493# sky130_fd_sc_hs__dfrtp_4_35/a_1678_395#
+ sky130_fd_sc_hs__dfrtp_4_35/a_1827_81# sky130_fd_sc_hs__dfrtp_4_35/a_789_463# sky130_fd_sc_hs__dfrtp_4_35/a_1350_392#
+ sky130_fd_sc_hs__dfrtp_4_35/a_834_355# sky130_fd_sc_hs__dfrtp_4_35/a_812_138# sky130_fd_sc_hs__dfrtp_4_35/a_124_78#
+ sky130_fd_sc_hs__dfrtp_4_35/a_1647_81# sky130_fd_sc_hs__dfrtp_4_35/a_2010_409# sky130_fd_sc_hs__dfrtp_4_35/a_890_138#
+ sky130_fd_sc_hs__dfrtp_4
Xsky130_fd_sc_hs__dfrtp_4_79 DVSS DVDD sky130_fd_sc_hs__clkbuf_8_1/X DVDD DVSS sky130_fd_sc_hs__dfrtp_4_79/D
+ sky130_fd_sc_hs__nand2_1_47/B sky130_fd_sc_hs__inv_4_41/A sky130_fd_sc_hs__dfrtp_4_79/a_37_78#
+ sky130_fd_sc_hs__dfrtp_4_79/a_494_366# sky130_fd_sc_hs__dfrtp_4_79/a_699_463# sky130_fd_sc_hs__dfrtp_4_79/a_313_74#
+ sky130_fd_sc_hs__dfrtp_4_79/a_1627_493# sky130_fd_sc_hs__dfrtp_4_79/a_1678_395#
+ sky130_fd_sc_hs__dfrtp_4_79/a_1827_81# sky130_fd_sc_hs__dfrtp_4_79/a_789_463# sky130_fd_sc_hs__dfrtp_4_79/a_1350_392#
+ sky130_fd_sc_hs__dfrtp_4_79/a_834_355# sky130_fd_sc_hs__dfrtp_4_79/a_812_138# sky130_fd_sc_hs__dfrtp_4_79/a_124_78#
+ sky130_fd_sc_hs__dfrtp_4_79/a_1647_81# sky130_fd_sc_hs__dfrtp_4_79/a_2010_409# sky130_fd_sc_hs__dfrtp_4_79/a_890_138#
+ sky130_fd_sc_hs__dfrtp_4
Xsky130_fd_sc_hs__nand2_1_70 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_95/Y sky130_fd_sc_hs__nand2_1_71/Y
+ sky130_fd_sc_hs__xnor2_1_9/A sky130_fd_sc_hs__nand2_1_71/a_117_74# sky130_fd_sc_hs__nand2_1
Xsky130_fd_sc_hs__nand2_1_92 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__o21a_1_63/A2 sky130_fd_sc_hs__nor2_1_63/B
+ sky130_fd_sc_hs__o21a_1_63/A1 sky130_fd_sc_hs__nand2_1_93/a_117_74# sky130_fd_sc_hs__nand2_1
Xsky130_fd_sc_hs__nand2_1_81 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_2_3/A sky130_fd_sc_hs__nand2_1_91/A
+ sky130_fd_sc_hs__inv_2_5/Y sky130_fd_sc_hs__nand2_1_81/a_117_74# sky130_fd_sc_hs__nand2_1
Xsky130_fd_sc_hs__nor2_1_8 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nor2_1_9/B sky130_fd_sc_hs__nor2_1_9/Y
+ sky130_fd_sc_hs__inv_4_9/Y sky130_fd_sc_hs__nor2_1_9/a_116_368# sky130_fd_sc_hs__nor2_1
Xsky130_fd_sc_hs__a21oi_1_38 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__a22oi_1_21/Y sky130_fd_sc_hs__o22ai_1_1/A1
+ sky130_fd_sc_hs__and2_2_1/X sky130_fd_sc_hs__xnor2_1_1/A sky130_fd_sc_hs__a21oi_1_39/a_117_74#
+ sky130_fd_sc_hs__a21oi_1_39/a_29_368# sky130_fd_sc_hs__a21oi_1
Xsky130_fd_sc_hs__a21oi_1_27 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__a21oi_1_17/Y sky130_fd_sc_hs__o31ai_1_1/B1
+ sky130_fd_sc_hs__a21oi_1_19/Y fine_control_avg_window_select[1] sky130_fd_sc_hs__a21oi_1_27/a_117_74#
+ sky130_fd_sc_hs__a21oi_1_27/a_29_368# sky130_fd_sc_hs__a21oi_1
Xsky130_fd_sc_hs__a21oi_1_16 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_1_15/Y sky130_fd_sc_hs__a21oi_1_17/Y
+ sky130_fd_sc_hs__a22oi_1_13/Y sky130_fd_sc_hs__a22oi_1_11/Y sky130_fd_sc_hs__a21oi_1_17/a_117_74#
+ sky130_fd_sc_hs__a21oi_1_17/a_29_368# sky130_fd_sc_hs__a21oi_1
Xsky130_fd_sc_hs__a21oi_1_49 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nor2_1_27/Y sky130_fd_sc_hs__dfrtn_1_3/D
+ sky130_fd_sc_hs__nor2_1_27/B sky130_fd_sc_hs__inv_4_37/Y sky130_fd_sc_hs__a21oi_1_49/a_117_74#
+ sky130_fd_sc_hs__a21oi_1_49/a_29_368# sky130_fd_sc_hs__a21oi_1
Xsky130_fd_sc_hs__nor3_1_12 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nor3_1_13/Y sky130_fd_sc_hs__nor3_1_13/C
+ sky130_fd_sc_hs__nor3_1_13/B sky130_fd_sc_hs__nor3_1_13/A sky130_fd_sc_hs__nor3_1_13/a_198_368#
+ sky130_fd_sc_hs__nor3_1_13/a_114_368# sky130_fd_sc_hs__nor3_1
Xsky130_fd_sc_hs__o21a_1_9 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__o21a_1_9/X sky130_fd_sc_hs__nor2_1_9/Y
+ sky130_fd_sc_hs__o21a_1_9/B1 sky130_fd_sc_hs__o21a_1_9/A1 sky130_fd_sc_hs__o21a_1_9/a_320_74#
+ sky130_fd_sc_hs__o21a_1_9/a_376_387# sky130_fd_sc_hs__o21a_1_9/a_83_244# sky130_fd_sc_hs__o21a_1
Xsky130_fd_sc_hs__nor2_1_101 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_121/Y sky130_fd_sc_hs__nor2_1_101/Y
+ sky130_fd_sc_hs__o21ai_1_7/Y sky130_fd_sc_hs__nor2_1_101/a_116_368# sky130_fd_sc_hs__nor2_1
Xsky130_fd_sc_hs__nor2_1_112 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__o21a_1_53/B1 sky130_fd_sc_hs__o21a_1_73/A2
+ sky130_fd_sc_hs__inv_4_117/Y sky130_fd_sc_hs__nor2_1_113/a_116_368# sky130_fd_sc_hs__nor2_1
Xsky130_fd_sc_hs__nor2_1_123 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__o21a_1_77/B1 sky130_fd_sc_hs__o21a_1_63/A2
+ sky130_fd_sc_hs__inv_4_137/Y sky130_fd_sc_hs__nor2_1_123/a_116_368# sky130_fd_sc_hs__nor2_1
Xsky130_fd_sc_hs__a22oi_1_10 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nor2b_1_25/Y sky130_fd_sc_hs__a22oi_1_11/Y
+ sky130_fd_sc_hs__inv_4_17/A sky130_fd_sc_hs__nor2b_1_23/Y sky130_fd_sc_hs__inv_4_11/A
+ sky130_fd_sc_hs__a22oi_1_11/a_71_368# sky130_fd_sc_hs__a22oi_1_11/a_159_74# sky130_fd_sc_hs__a22oi_1_11/a_339_74#
+ sky130_fd_sc_hs__a22oi_1
Xsky130_fd_sc_hs__a22oi_1_21 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_33/Y sky130_fd_sc_hs__a22oi_1_21/Y
+ sky130_fd_sc_hs__a32oi_1_5/A1 sky130_fd_sc_hs__a222oi_1_1/Y fine_control_avg_window_select[0]
+ sky130_fd_sc_hs__a22oi_1_21/a_71_368# sky130_fd_sc_hs__a22oi_1_21/a_159_74# sky130_fd_sc_hs__a22oi_1_21/a_339_74#
+ sky130_fd_sc_hs__a22oi_1
Xsky130_fd_sc_hs__fa_2_17 DVSS DVDD sky130_fd_sc_hs__fa_2_9/B DVDD DVSS sky130_fd_sc_hs__fa_2_17/CIN
+ sky130_fd_sc_hs__fa_2_17/B sky130_fd_sc_hs__fa_2_19/CIN sky130_fd_sc_hs__fa_2_17/SUM
+ sky130_fd_sc_hs__fa_2_17/a_27_378# sky130_fd_sc_hs__fa_2_17/a_701_79# sky130_fd_sc_hs__fa_2_17/a_484_347#
+ sky130_fd_sc_hs__fa_2_17/a_1094_347# sky130_fd_sc_hs__fa_2_17/a_1205_79# sky130_fd_sc_hs__fa_2_17/a_27_79#
+ sky130_fd_sc_hs__fa_2_17/a_1202_368# sky130_fd_sc_hs__fa_2_17/a_336_347# sky130_fd_sc_hs__fa_2_17/a_992_347#
+ sky130_fd_sc_hs__fa_2_17/a_1119_79# sky130_fd_sc_hs__fa_2_17/a_487_79# sky130_fd_sc_hs__fa_2_17/a_683_347#
+ sky130_fd_sc_hs__fa_2
Xsky130_fd_sc_hs__dfsbp_2_1 DVSS DVDD sky130_fd_sc_hs__inv_4_49/Y DVDD DVSS sky130_fd_sc_hs__o21ai_1_1/Y
+ sky130_fd_sc_hs__dfstp_2_7/Q sky130_fd_sc_hs__inv_4_23/A sky130_fd_sc_hs__dfsbp_2_1/Q
+ sky130_fd_sc_hs__dfsbp_2_1/a_595_97# sky130_fd_sc_hs__dfsbp_2_1/a_731_97# sky130_fd_sc_hs__dfsbp_2_1/a_1521_508#
+ sky130_fd_sc_hs__dfsbp_2_1/a_2221_74# sky130_fd_sc_hs__dfsbp_2_1/a_1339_74# sky130_fd_sc_hs__dfsbp_2_1/a_1531_118#
+ sky130_fd_sc_hs__dfsbp_2_1/a_1453_118# sky130_fd_sc_hs__dfsbp_2_1/a_398_74# sky130_fd_sc_hs__dfsbp_2_1/a_27_74#
+ sky130_fd_sc_hs__dfsbp_2_1/a_225_74# sky130_fd_sc_hs__dfsbp_2_1/a_1501_92# sky130_fd_sc_hs__dfsbp_2_1/a_757_401#
+ sky130_fd_sc_hs__dfsbp_2_1/a_1258_341# sky130_fd_sc_hs__dfsbp_2_1/a_1001_74# sky130_fd_sc_hs__dfsbp_2_1/a_706_463#
+ sky130_fd_sc_hs__dfsbp_2_1/a_1261_74# sky130_fd_sc_hs__dfsbp_2
Xsky130_fd_sc_hs__or3b_2_0 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__or3b_2_1/X rst sky130_fd_sc_hs__or3b_2_1/B
+ sky130_fd_sc_hs__or3b_2_1/C_N sky130_fd_sc_hs__or3b_2_1/a_542_368# sky130_fd_sc_hs__or3b_2_1/a_27_368#
+ sky130_fd_sc_hs__or3b_2_1/a_190_260# sky130_fd_sc_hs__or3b_2_1/a_458_368# sky130_fd_sc_hs__or3b_2
Xsky130_fd_sc_hs__nand2b_4_1 DVSS DVDD DVDD DVSS div_ratio_half[4] sky130_fd_sc_hs__xnor2_1_13/A
+ sky130_fd_sc_hs__inv_4_103/A sky130_fd_sc_hs__nand2b_4_1/a_31_74# sky130_fd_sc_hs__nand2b_4_1/a_243_74#
+ sky130_fd_sc_hs__nand2b_4
Xsky130_fd_sc_hs__o21a_1_24 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__o21a_1_25/X sky130_fd_sc_hs__nor2_1_25/Y
+ sky130_fd_sc_hs__nor2_1_19/B sky130_fd_sc_hs__o21a_1_25/A1 sky130_fd_sc_hs__o21a_1_25/a_320_74#
+ sky130_fd_sc_hs__o21a_1_25/a_376_387# sky130_fd_sc_hs__o21a_1_25/a_83_244# sky130_fd_sc_hs__o21a_1
Xsky130_fd_sc_hs__o21a_1_13 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__o21a_1_13/X sky130_fd_sc_hs__nor2_1_11/Y
+ sky130_fd_sc_hs__nor2_1_31/B sky130_fd_sc_hs__o21a_1_13/A1 sky130_fd_sc_hs__o21a_1_13/a_320_74#
+ sky130_fd_sc_hs__o21a_1_13/a_376_387# sky130_fd_sc_hs__o21a_1_13/a_83_244# sky130_fd_sc_hs__o21a_1
Xsky130_fd_sc_hs__o21a_1_57 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__o21a_1_57/X sky130_fd_sc_hs__nor2_1_47/Y
+ sky130_fd_sc_hs__o21a_1_57/B1 sky130_fd_sc_hs__inv_4_93/A sky130_fd_sc_hs__o21a_1_57/a_320_74#
+ sky130_fd_sc_hs__o21a_1_57/a_376_387# sky130_fd_sc_hs__o21a_1_57/a_83_244# sky130_fd_sc_hs__o21a_1
Xsky130_fd_sc_hs__o21a_1_46 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__o21a_1_47/X sky130_fd_sc_hs__nor2_1_51/Y
+ sky130_fd_sc_hs__nor2_1_57/B sky130_fd_sc_hs__nor2_1_59/A sky130_fd_sc_hs__o21a_1_47/a_320_74#
+ sky130_fd_sc_hs__o21a_1_47/a_376_387# sky130_fd_sc_hs__o21a_1_47/a_83_244# sky130_fd_sc_hs__o21a_1
Xsky130_fd_sc_hs__o21a_1_35 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__o21a_1_35/X sky130_fd_sc_hs__nor2_1_41/Y
+ sky130_fd_sc_hs__nor2_1_51/B sky130_fd_sc_hs__dfrbp_1_1/Q sky130_fd_sc_hs__o21a_1_35/a_320_74#
+ sky130_fd_sc_hs__o21a_1_35/a_376_387# sky130_fd_sc_hs__o21a_1_35/a_83_244# sky130_fd_sc_hs__o21a_1
Xsky130_fd_sc_hs__o21a_1_68 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__o21a_1_69/X sky130_fd_sc_hs__o21a_1_69/A2
+ sky130_fd_sc_hs__xnor2_1_9/B sky130_fd_sc_hs__inv_4_127/A sky130_fd_sc_hs__o21a_1_69/a_320_74#
+ sky130_fd_sc_hs__o21a_1_69/a_376_387# sky130_fd_sc_hs__o21a_1_69/a_83_244# sky130_fd_sc_hs__o21a_1
Xsky130_fd_sc_hs__dfrtp_4_25 DVSS DVDD sky130_fd_sc_hs__clkbuf_8_1/X DVDD DVSS sky130_fd_sc_hs__dfrtp_4_25/D
+ sky130_fd_sc_hs__nand2_1_47/B sky130_fd_sc_hs__inv_4_13/A sky130_fd_sc_hs__dfrtp_4_25/a_37_78#
+ sky130_fd_sc_hs__dfrtp_4_25/a_494_366# sky130_fd_sc_hs__dfrtp_4_25/a_699_463# sky130_fd_sc_hs__dfrtp_4_25/a_313_74#
+ sky130_fd_sc_hs__dfrtp_4_25/a_1627_493# sky130_fd_sc_hs__dfrtp_4_25/a_1678_395#
+ sky130_fd_sc_hs__dfrtp_4_25/a_1827_81# sky130_fd_sc_hs__dfrtp_4_25/a_789_463# sky130_fd_sc_hs__dfrtp_4_25/a_1350_392#
+ sky130_fd_sc_hs__dfrtp_4_25/a_834_355# sky130_fd_sc_hs__dfrtp_4_25/a_812_138# sky130_fd_sc_hs__dfrtp_4_25/a_124_78#
+ sky130_fd_sc_hs__dfrtp_4_25/a_1647_81# sky130_fd_sc_hs__dfrtp_4_25/a_2010_409# sky130_fd_sc_hs__dfrtp_4_25/a_890_138#
+ sky130_fd_sc_hs__dfrtp_4
Xsky130_fd_sc_hs__dfrtp_4_14 DVSS DVDD sky130_fd_sc_hs__inv_4_49/Y DVDD DVSS sky130_fd_sc_hs__nor2b_1_1/Y
+ sky130_fd_sc_hs__dfstp_2_1/CLK sky130_fd_sc_hs__fa_2_1/B sky130_fd_sc_hs__dfrtp_4_15/a_37_78#
+ sky130_fd_sc_hs__dfrtp_4_15/a_494_366# sky130_fd_sc_hs__dfrtp_4_15/a_699_463# sky130_fd_sc_hs__dfrtp_4_15/a_313_74#
+ sky130_fd_sc_hs__dfrtp_4_15/a_1627_493# sky130_fd_sc_hs__dfrtp_4_15/a_1678_395#
+ sky130_fd_sc_hs__dfrtp_4_15/a_1827_81# sky130_fd_sc_hs__dfrtp_4_15/a_789_463# sky130_fd_sc_hs__dfrtp_4_15/a_1350_392#
+ sky130_fd_sc_hs__dfrtp_4_15/a_834_355# sky130_fd_sc_hs__dfrtp_4_15/a_812_138# sky130_fd_sc_hs__dfrtp_4_15/a_124_78#
+ sky130_fd_sc_hs__dfrtp_4_15/a_1647_81# sky130_fd_sc_hs__dfrtp_4_15/a_2010_409# sky130_fd_sc_hs__dfrtp_4_15/a_890_138#
+ sky130_fd_sc_hs__dfrtp_4
Xsky130_fd_sc_hs__dfrtp_4_58 DVSS DVDD sky130_fd_sc_hs__clkbuf_8_1/X DVDD DVSS sky130_fd_sc_hs__dfrtp_4_59/D
+ sky130_fd_sc_hs__nand2_1_47/B sky130_fd_sc_hs__inv_4_31/A sky130_fd_sc_hs__dfrtp_4_59/a_37_78#
+ sky130_fd_sc_hs__dfrtp_4_59/a_494_366# sky130_fd_sc_hs__dfrtp_4_59/a_699_463# sky130_fd_sc_hs__dfrtp_4_59/a_313_74#
+ sky130_fd_sc_hs__dfrtp_4_59/a_1627_493# sky130_fd_sc_hs__dfrtp_4_59/a_1678_395#
+ sky130_fd_sc_hs__dfrtp_4_59/a_1827_81# sky130_fd_sc_hs__dfrtp_4_59/a_789_463# sky130_fd_sc_hs__dfrtp_4_59/a_1350_392#
+ sky130_fd_sc_hs__dfrtp_4_59/a_834_355# sky130_fd_sc_hs__dfrtp_4_59/a_812_138# sky130_fd_sc_hs__dfrtp_4_59/a_124_78#
+ sky130_fd_sc_hs__dfrtp_4_59/a_1647_81# sky130_fd_sc_hs__dfrtp_4_59/a_2010_409# sky130_fd_sc_hs__dfrtp_4_59/a_890_138#
+ sky130_fd_sc_hs__dfrtp_4
Xsky130_fd_sc_hs__dfrtp_4_47 DVSS DVDD sky130_fd_sc_hs__inv_4_49/Y DVDD DVSS sky130_fd_sc_hs__nor2b_1_11/Y
+ sky130_fd_sc_hs__dfstp_2_1/CLK sky130_fd_sc_hs__fa_2_9/A sky130_fd_sc_hs__dfrtp_4_47/a_37_78#
+ sky130_fd_sc_hs__dfrtp_4_47/a_494_366# sky130_fd_sc_hs__dfrtp_4_47/a_699_463# sky130_fd_sc_hs__dfrtp_4_47/a_313_74#
+ sky130_fd_sc_hs__dfrtp_4_47/a_1627_493# sky130_fd_sc_hs__dfrtp_4_47/a_1678_395#
+ sky130_fd_sc_hs__dfrtp_4_47/a_1827_81# sky130_fd_sc_hs__dfrtp_4_47/a_789_463# sky130_fd_sc_hs__dfrtp_4_47/a_1350_392#
+ sky130_fd_sc_hs__dfrtp_4_47/a_834_355# sky130_fd_sc_hs__dfrtp_4_47/a_812_138# sky130_fd_sc_hs__dfrtp_4_47/a_124_78#
+ sky130_fd_sc_hs__dfrtp_4_47/a_1647_81# sky130_fd_sc_hs__dfrtp_4_47/a_2010_409# sky130_fd_sc_hs__dfrtp_4_47/a_890_138#
+ sky130_fd_sc_hs__dfrtp_4
Xsky130_fd_sc_hs__dfrtp_4_36 DVSS DVDD sky130_fd_sc_hs__inv_4_49/Y DVDD DVSS sky130_fd_sc_hs__nor2b_1_5/Y
+ sky130_fd_sc_hs__dfstp_2_1/CLK sky130_fd_sc_hs__fa_2_5/B sky130_fd_sc_hs__dfrtp_4_37/a_37_78#
+ sky130_fd_sc_hs__dfrtp_4_37/a_494_366# sky130_fd_sc_hs__dfrtp_4_37/a_699_463# sky130_fd_sc_hs__dfrtp_4_37/a_313_74#
+ sky130_fd_sc_hs__dfrtp_4_37/a_1627_493# sky130_fd_sc_hs__dfrtp_4_37/a_1678_395#
+ sky130_fd_sc_hs__dfrtp_4_37/a_1827_81# sky130_fd_sc_hs__dfrtp_4_37/a_789_463# sky130_fd_sc_hs__dfrtp_4_37/a_1350_392#
+ sky130_fd_sc_hs__dfrtp_4_37/a_834_355# sky130_fd_sc_hs__dfrtp_4_37/a_812_138# sky130_fd_sc_hs__dfrtp_4_37/a_124_78#
+ sky130_fd_sc_hs__dfrtp_4_37/a_1647_81# sky130_fd_sc_hs__dfrtp_4_37/a_2010_409# sky130_fd_sc_hs__dfrtp_4_37/a_890_138#
+ sky130_fd_sc_hs__dfrtp_4
Xsky130_fd_sc_hs__dfrtp_4_69 DVSS DVDD sky130_fd_sc_hs__clkbuf_8_1/A DVDD DVSS sky130_fd_sc_hs__xnor2_1_1/Y
+ sky130_fd_sc_hs__nand2_1_47/B sky130_fd_sc_hs__xnor2_1_1/A sky130_fd_sc_hs__dfrtp_4_69/a_37_78#
+ sky130_fd_sc_hs__dfrtp_4_69/a_494_366# sky130_fd_sc_hs__dfrtp_4_69/a_699_463# sky130_fd_sc_hs__dfrtp_4_69/a_313_74#
+ sky130_fd_sc_hs__dfrtp_4_69/a_1627_493# sky130_fd_sc_hs__dfrtp_4_69/a_1678_395#
+ sky130_fd_sc_hs__dfrtp_4_69/a_1827_81# sky130_fd_sc_hs__dfrtp_4_69/a_789_463# sky130_fd_sc_hs__dfrtp_4_69/a_1350_392#
+ sky130_fd_sc_hs__dfrtp_4_69/a_834_355# sky130_fd_sc_hs__dfrtp_4_69/a_812_138# sky130_fd_sc_hs__dfrtp_4_69/a_124_78#
+ sky130_fd_sc_hs__dfrtp_4_69/a_1647_81# sky130_fd_sc_hs__dfrtp_4_69/a_2010_409# sky130_fd_sc_hs__dfrtp_4_69/a_890_138#
+ sky130_fd_sc_hs__dfrtp_4
Xsky130_fd_sc_hs__nand2_1_60 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nor2_1_87/Y sky130_fd_sc_hs__nor2_1_45/B
+ sky130_fd_sc_hs__inv_4_83/A sky130_fd_sc_hs__nand2_1_61/a_117_74# sky130_fd_sc_hs__nand2_1
Xsky130_fd_sc_hs__nand2_1_93 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__o21a_1_63/A2 sky130_fd_sc_hs__nor2_1_63/B
+ sky130_fd_sc_hs__o21a_1_63/A1 sky130_fd_sc_hs__nand2_1_93/a_117_74# sky130_fd_sc_hs__nand2_1
Xsky130_fd_sc_hs__nand2_1_82 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__o21a_1_61/A2 sky130_fd_sc_hs__xnor2_1_5/B
+ sky130_fd_sc_hs__maj3_1_3/A sky130_fd_sc_hs__nand2_1_83/a_117_74# sky130_fd_sc_hs__nand2_1
Xsky130_fd_sc_hs__nand2_1_71 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_95/Y sky130_fd_sc_hs__nand2_1_71/Y
+ sky130_fd_sc_hs__xnor2_1_9/A sky130_fd_sc_hs__nand2_1_71/a_117_74# sky130_fd_sc_hs__nand2_1
Xsky130_fd_sc_hs__nor2_1_9 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nor2_1_9/B sky130_fd_sc_hs__nor2_1_9/Y
+ sky130_fd_sc_hs__inv_4_9/Y sky130_fd_sc_hs__nor2_1_9/a_116_368# sky130_fd_sc_hs__nor2_1
Xsky130_fd_sc_hs__a21oi_1_28 DVSS DVDD DVDD DVSS fine_control_avg_window_select[2]
+ sky130_fd_sc_hs__nand2_2_3/B sky130_fd_sc_hs__and2_2_1/X sky130_fd_sc_hs__o21a_1_19/A1
+ sky130_fd_sc_hs__a21oi_1_29/a_117_74# sky130_fd_sc_hs__a21oi_1_29/a_29_368# sky130_fd_sc_hs__a21oi_1
Xsky130_fd_sc_hs__a21oi_1_17 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_1_15/Y sky130_fd_sc_hs__a21oi_1_17/Y
+ sky130_fd_sc_hs__a22oi_1_13/Y sky130_fd_sc_hs__a22oi_1_11/Y sky130_fd_sc_hs__a21oi_1_17/a_117_74#
+ sky130_fd_sc_hs__a21oi_1_17/a_29_368# sky130_fd_sc_hs__a21oi_1
Xsky130_fd_sc_hs__a21oi_1_39 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__a22oi_1_21/Y sky130_fd_sc_hs__o22ai_1_1/A1
+ sky130_fd_sc_hs__and2_2_1/X sky130_fd_sc_hs__xnor2_1_1/A sky130_fd_sc_hs__a21oi_1_39/a_117_74#
+ sky130_fd_sc_hs__a21oi_1_39/a_29_368# sky130_fd_sc_hs__a21oi_1
Xsky130_fd_sc_hs__nand2_4_0 DVSS DVDD DVDD DVSS aux_clk_out aux_osc_en sky130_fd_sc_hs__nand2_4_5/Y
+ sky130_fd_sc_hs__nand2_4_1/a_27_74# sky130_fd_sc_hs__nand2_4
Xsky130_fd_sc_hs__nor3_1_13 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nor3_1_13/Y sky130_fd_sc_hs__nor3_1_13/C
+ sky130_fd_sc_hs__nor3_1_13/B sky130_fd_sc_hs__nor3_1_13/A sky130_fd_sc_hs__nor3_1_13/a_198_368#
+ sky130_fd_sc_hs__nor3_1_13/a_114_368# sky130_fd_sc_hs__nor3_1
Xsky130_fd_sc_hs__nor2_1_102 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__o21a_1_57/B1 sky130_fd_sc_hs__o21a_1_67/A2
+ sky130_fd_sc_hs__nor2_1_95/B sky130_fd_sc_hs__nor2_1_103/a_116_368# sky130_fd_sc_hs__nor2_1
Xsky130_fd_sc_hs__nor2_1_113 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__o21a_1_53/B1 sky130_fd_sc_hs__o21a_1_73/A2
+ sky130_fd_sc_hs__inv_4_117/Y sky130_fd_sc_hs__nor2_1_113/a_116_368# sky130_fd_sc_hs__nor2_1
Xsky130_fd_sc_hs__a22oi_1_22 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nor4_1_3/C sky130_fd_sc_hs__a22oi_1_23/Y
+ sky130_fd_sc_hs__a21oi_1_97/Y sky130_fd_sc_hs__nand2_1_85/Y sky130_fd_sc_hs__nor3_1_5/C
+ sky130_fd_sc_hs__a22oi_1_23/a_71_368# sky130_fd_sc_hs__a22oi_1_23/a_159_74# sky130_fd_sc_hs__a22oi_1_23/a_339_74#
+ sky130_fd_sc_hs__a22oi_1
Xsky130_fd_sc_hs__a22oi_1_11 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nor2b_1_25/Y sky130_fd_sc_hs__a22oi_1_11/Y
+ sky130_fd_sc_hs__inv_4_17/A sky130_fd_sc_hs__nor2b_1_23/Y sky130_fd_sc_hs__inv_4_11/A
+ sky130_fd_sc_hs__a22oi_1_11/a_71_368# sky130_fd_sc_hs__a22oi_1_11/a_159_74# sky130_fd_sc_hs__a22oi_1_11/a_339_74#
+ sky130_fd_sc_hs__a22oi_1
Xsky130_fd_sc_hs__nor2_1_90 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nor2_1_91/B sky130_fd_sc_hs__nor2_1_91/Y
+ sky130_fd_sc_hs__xnor2_1_7/Y sky130_fd_sc_hs__nor2_1_91/a_116_368# sky130_fd_sc_hs__nor2_1
Xsky130_fd_sc_hs__fa_2_18 DVSS DVDD sky130_fd_sc_hs__fa_2_9/B DVDD DVSS sky130_fd_sc_hs__fa_2_19/CIN
+ sky130_fd_sc_hs__fa_2_19/B sky130_fd_sc_hs__fa_2_21/CIN sky130_fd_sc_hs__fa_2_19/SUM
+ sky130_fd_sc_hs__fa_2_19/a_27_378# sky130_fd_sc_hs__fa_2_19/a_701_79# sky130_fd_sc_hs__fa_2_19/a_484_347#
+ sky130_fd_sc_hs__fa_2_19/a_1094_347# sky130_fd_sc_hs__fa_2_19/a_1205_79# sky130_fd_sc_hs__fa_2_19/a_27_79#
+ sky130_fd_sc_hs__fa_2_19/a_1202_368# sky130_fd_sc_hs__fa_2_19/a_336_347# sky130_fd_sc_hs__fa_2_19/a_992_347#
+ sky130_fd_sc_hs__fa_2_19/a_1119_79# sky130_fd_sc_hs__fa_2_19/a_487_79# sky130_fd_sc_hs__fa_2_19/a_683_347#
+ sky130_fd_sc_hs__fa_2
Xsky130_fd_sc_hs__or3b_2_1 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__or3b_2_1/X rst sky130_fd_sc_hs__or3b_2_1/B
+ sky130_fd_sc_hs__or3b_2_1/C_N sky130_fd_sc_hs__or3b_2_1/a_542_368# sky130_fd_sc_hs__or3b_2_1/a_27_368#
+ sky130_fd_sc_hs__or3b_2_1/a_190_260# sky130_fd_sc_hs__or3b_2_1/a_458_368# sky130_fd_sc_hs__or3b_2
Xsky130_fd_sc_hs__o21a_1_14 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__o21a_1_15/X sky130_fd_sc_hs__nor2_1_7/Y
+ sky130_fd_sc_hs__nor2_1_35/B sky130_fd_sc_hs__o21a_1_15/A1 sky130_fd_sc_hs__o21a_1_15/a_320_74#
+ sky130_fd_sc_hs__o21a_1_15/a_376_387# sky130_fd_sc_hs__o21a_1_15/a_83_244# sky130_fd_sc_hs__o21a_1
Xsky130_fd_sc_hs__o21a_1_58 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__o21a_1_59/X sky130_fd_sc_hs__o21a_1_59/A2
+ sky130_fd_sc_hs__nor2_1_87/B sky130_fd_sc_hs__o21a_1_59/A1 sky130_fd_sc_hs__o21a_1_59/a_320_74#
+ sky130_fd_sc_hs__o21a_1_59/a_376_387# sky130_fd_sc_hs__o21a_1_59/a_83_244# sky130_fd_sc_hs__o21a_1
Xsky130_fd_sc_hs__o21a_1_47 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__o21a_1_47/X sky130_fd_sc_hs__nor2_1_51/Y
+ sky130_fd_sc_hs__nor2_1_57/B sky130_fd_sc_hs__nor2_1_59/A sky130_fd_sc_hs__o21a_1_47/a_320_74#
+ sky130_fd_sc_hs__o21a_1_47/a_376_387# sky130_fd_sc_hs__o21a_1_47/a_83_244# sky130_fd_sc_hs__o21a_1
Xsky130_fd_sc_hs__o21a_1_36 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__o21a_1_37/X sky130_fd_sc_hs__nor2_1_45/Y
+ sky130_fd_sc_hs__nor2_1_29/B sky130_fd_sc_hs__nor2_1_65/A sky130_fd_sc_hs__o21a_1_37/a_320_74#
+ sky130_fd_sc_hs__o21a_1_37/a_376_387# sky130_fd_sc_hs__o21a_1_37/a_83_244# sky130_fd_sc_hs__o21a_1
Xsky130_fd_sc_hs__o21a_1_25 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__o21a_1_25/X sky130_fd_sc_hs__nor2_1_25/Y
+ sky130_fd_sc_hs__nor2_1_19/B sky130_fd_sc_hs__o21a_1_25/A1 sky130_fd_sc_hs__o21a_1_25/a_320_74#
+ sky130_fd_sc_hs__o21a_1_25/a_376_387# sky130_fd_sc_hs__o21a_1_25/a_83_244# sky130_fd_sc_hs__o21a_1
Xsky130_fd_sc_hs__o21a_1_69 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__o21a_1_69/X sky130_fd_sc_hs__o21a_1_69/A2
+ sky130_fd_sc_hs__xnor2_1_9/B sky130_fd_sc_hs__inv_4_127/A sky130_fd_sc_hs__o21a_1_69/a_320_74#
+ sky130_fd_sc_hs__o21a_1_69/a_376_387# sky130_fd_sc_hs__o21a_1_69/a_83_244# sky130_fd_sc_hs__o21a_1
Xsky130_fd_sc_hs__dfrtp_4_15 DVSS DVDD sky130_fd_sc_hs__inv_4_49/Y DVDD DVSS sky130_fd_sc_hs__nor2b_1_1/Y
+ sky130_fd_sc_hs__dfstp_2_1/CLK sky130_fd_sc_hs__fa_2_1/B sky130_fd_sc_hs__dfrtp_4_15/a_37_78#
+ sky130_fd_sc_hs__dfrtp_4_15/a_494_366# sky130_fd_sc_hs__dfrtp_4_15/a_699_463# sky130_fd_sc_hs__dfrtp_4_15/a_313_74#
+ sky130_fd_sc_hs__dfrtp_4_15/a_1627_493# sky130_fd_sc_hs__dfrtp_4_15/a_1678_395#
+ sky130_fd_sc_hs__dfrtp_4_15/a_1827_81# sky130_fd_sc_hs__dfrtp_4_15/a_789_463# sky130_fd_sc_hs__dfrtp_4_15/a_1350_392#
+ sky130_fd_sc_hs__dfrtp_4_15/a_834_355# sky130_fd_sc_hs__dfrtp_4_15/a_812_138# sky130_fd_sc_hs__dfrtp_4_15/a_124_78#
+ sky130_fd_sc_hs__dfrtp_4_15/a_1647_81# sky130_fd_sc_hs__dfrtp_4_15/a_2010_409# sky130_fd_sc_hs__dfrtp_4_15/a_890_138#
+ sky130_fd_sc_hs__dfrtp_4
Xsky130_fd_sc_hs__dfrtp_4_59 DVSS DVDD sky130_fd_sc_hs__clkbuf_8_1/X DVDD DVSS sky130_fd_sc_hs__dfrtp_4_59/D
+ sky130_fd_sc_hs__nand2_1_47/B sky130_fd_sc_hs__inv_4_31/A sky130_fd_sc_hs__dfrtp_4_59/a_37_78#
+ sky130_fd_sc_hs__dfrtp_4_59/a_494_366# sky130_fd_sc_hs__dfrtp_4_59/a_699_463# sky130_fd_sc_hs__dfrtp_4_59/a_313_74#
+ sky130_fd_sc_hs__dfrtp_4_59/a_1627_493# sky130_fd_sc_hs__dfrtp_4_59/a_1678_395#
+ sky130_fd_sc_hs__dfrtp_4_59/a_1827_81# sky130_fd_sc_hs__dfrtp_4_59/a_789_463# sky130_fd_sc_hs__dfrtp_4_59/a_1350_392#
+ sky130_fd_sc_hs__dfrtp_4_59/a_834_355# sky130_fd_sc_hs__dfrtp_4_59/a_812_138# sky130_fd_sc_hs__dfrtp_4_59/a_124_78#
+ sky130_fd_sc_hs__dfrtp_4_59/a_1647_81# sky130_fd_sc_hs__dfrtp_4_59/a_2010_409# sky130_fd_sc_hs__dfrtp_4_59/a_890_138#
+ sky130_fd_sc_hs__dfrtp_4
Xsky130_fd_sc_hs__dfrtp_4_48 DVSS DVDD sky130_fd_sc_hs__clkbuf_8_1/X DVDD DVSS sky130_fd_sc_hs__o21a_1_21/X
+ sky130_fd_sc_hs__nand2_1_47/B sky130_fd_sc_hs__o21a_1_21/A1 sky130_fd_sc_hs__dfrtp_4_49/a_37_78#
+ sky130_fd_sc_hs__dfrtp_4_49/a_494_366# sky130_fd_sc_hs__dfrtp_4_49/a_699_463# sky130_fd_sc_hs__dfrtp_4_49/a_313_74#
+ sky130_fd_sc_hs__dfrtp_4_49/a_1627_493# sky130_fd_sc_hs__dfrtp_4_49/a_1678_395#
+ sky130_fd_sc_hs__dfrtp_4_49/a_1827_81# sky130_fd_sc_hs__dfrtp_4_49/a_789_463# sky130_fd_sc_hs__dfrtp_4_49/a_1350_392#
+ sky130_fd_sc_hs__dfrtp_4_49/a_834_355# sky130_fd_sc_hs__dfrtp_4_49/a_812_138# sky130_fd_sc_hs__dfrtp_4_49/a_124_78#
+ sky130_fd_sc_hs__dfrtp_4_49/a_1647_81# sky130_fd_sc_hs__dfrtp_4_49/a_2010_409# sky130_fd_sc_hs__dfrtp_4_49/a_890_138#
+ sky130_fd_sc_hs__dfrtp_4
Xsky130_fd_sc_hs__dfrtp_4_37 DVSS DVDD sky130_fd_sc_hs__inv_4_49/Y DVDD DVSS sky130_fd_sc_hs__nor2b_1_5/Y
+ sky130_fd_sc_hs__dfstp_2_1/CLK sky130_fd_sc_hs__fa_2_5/B sky130_fd_sc_hs__dfrtp_4_37/a_37_78#
+ sky130_fd_sc_hs__dfrtp_4_37/a_494_366# sky130_fd_sc_hs__dfrtp_4_37/a_699_463# sky130_fd_sc_hs__dfrtp_4_37/a_313_74#
+ sky130_fd_sc_hs__dfrtp_4_37/a_1627_493# sky130_fd_sc_hs__dfrtp_4_37/a_1678_395#
+ sky130_fd_sc_hs__dfrtp_4_37/a_1827_81# sky130_fd_sc_hs__dfrtp_4_37/a_789_463# sky130_fd_sc_hs__dfrtp_4_37/a_1350_392#
+ sky130_fd_sc_hs__dfrtp_4_37/a_834_355# sky130_fd_sc_hs__dfrtp_4_37/a_812_138# sky130_fd_sc_hs__dfrtp_4_37/a_124_78#
+ sky130_fd_sc_hs__dfrtp_4_37/a_1647_81# sky130_fd_sc_hs__dfrtp_4_37/a_2010_409# sky130_fd_sc_hs__dfrtp_4_37/a_890_138#
+ sky130_fd_sc_hs__dfrtp_4
Xsky130_fd_sc_hs__dfrtp_4_26 DVSS DVDD sky130_fd_sc_hs__clkbuf_8_1/A DVDD DVSS sky130_fd_sc_hs__o21a_1_9/X
+ sky130_fd_sc_hs__nand2_1_47/B sky130_fd_sc_hs__o21a_1_9/A1 sky130_fd_sc_hs__dfrtp_4_27/a_37_78#
+ sky130_fd_sc_hs__dfrtp_4_27/a_494_366# sky130_fd_sc_hs__dfrtp_4_27/a_699_463# sky130_fd_sc_hs__dfrtp_4_27/a_313_74#
+ sky130_fd_sc_hs__dfrtp_4_27/a_1627_493# sky130_fd_sc_hs__dfrtp_4_27/a_1678_395#
+ sky130_fd_sc_hs__dfrtp_4_27/a_1827_81# sky130_fd_sc_hs__dfrtp_4_27/a_789_463# sky130_fd_sc_hs__dfrtp_4_27/a_1350_392#
+ sky130_fd_sc_hs__dfrtp_4_27/a_834_355# sky130_fd_sc_hs__dfrtp_4_27/a_812_138# sky130_fd_sc_hs__dfrtp_4_27/a_124_78#
+ sky130_fd_sc_hs__dfrtp_4_27/a_1647_81# sky130_fd_sc_hs__dfrtp_4_27/a_2010_409# sky130_fd_sc_hs__dfrtp_4_27/a_890_138#
+ sky130_fd_sc_hs__dfrtp_4
Xsky130_fd_sc_hs__inv_4_0 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_1/Y sky130_fd_sc_hs__inv_4_1/A
+ sky130_fd_sc_hs__inv_4
Xsky130_fd_sc_hs__nand4_1_0 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand4_1_1/C sky130_fd_sc_hs__nand4_1_1/Y
+ sky130_fd_sc_hs__nand4_1_1/D sky130_fd_sc_hs__nor3_1_9/Y sky130_fd_sc_hs__nor3_1_1/Y
+ sky130_fd_sc_hs__nand4_1_1/a_259_74# sky130_fd_sc_hs__nand4_1_1/a_373_74# sky130_fd_sc_hs__nand4_1_1/a_181_74#
+ sky130_fd_sc_hs__nand4_1
Xsky130_fd_sc_hs__nand2_1_50 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_53/Y sky130_fd_sc_hs__nand2_1_51/Y
+ sky130_fd_sc_hs__inv_4_51/A sky130_fd_sc_hs__nand2_1_51/a_117_74# sky130_fd_sc_hs__nand2_1
Xsky130_fd_sc_hs__nand2_1_94 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_129/Y sky130_fd_sc_hs__nand4_1_5/D
+ sky130_fd_sc_hs__inv_4_137/A sky130_fd_sc_hs__nand2_1_95/a_117_74# sky130_fd_sc_hs__nand2_1
Xsky130_fd_sc_hs__nand2_1_83 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__o21a_1_61/A2 sky130_fd_sc_hs__xnor2_1_5/B
+ sky130_fd_sc_hs__maj3_1_3/A sky130_fd_sc_hs__nand2_1_83/a_117_74# sky130_fd_sc_hs__nand2_1
Xsky130_fd_sc_hs__nand2_1_72 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nor2_1_73/Y sky130_fd_sc_hs__o21a_1_53/B1
+ sky130_fd_sc_hs__o22ai_1_7/A1 sky130_fd_sc_hs__nand2_1_73/a_117_74# sky130_fd_sc_hs__nand2_1
Xsky130_fd_sc_hs__nand2_1_61 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nor2_1_87/Y sky130_fd_sc_hs__nor2_1_45/B
+ sky130_fd_sc_hs__inv_4_83/A sky130_fd_sc_hs__nand2_1_61/a_117_74# sky130_fd_sc_hs__nand2_1
Xsky130_fd_sc_hs__a21oi_1_29 DVSS DVDD DVDD DVSS fine_control_avg_window_select[2]
+ sky130_fd_sc_hs__nand2_2_3/B sky130_fd_sc_hs__and2_2_1/X sky130_fd_sc_hs__o21a_1_19/A1
+ sky130_fd_sc_hs__a21oi_1_29/a_117_74# sky130_fd_sc_hs__a21oi_1_29/a_29_368# sky130_fd_sc_hs__a21oi_1
Xsky130_fd_sc_hs__a21oi_1_18 DVSS DVDD DVDD DVSS fine_control_avg_window_select[2]
+ sky130_fd_sc_hs__a21oi_1_19/Y sky130_fd_sc_hs__a22oi_1_1/Y sky130_fd_sc_hs__a22oi_1_5/Y
+ sky130_fd_sc_hs__a21oi_1_19/a_117_74# sky130_fd_sc_hs__a21oi_1_19/a_29_368# sky130_fd_sc_hs__a21oi_1
Xsky130_fd_sc_hs__nand2_4_1 DVSS DVDD DVDD DVSS aux_clk_out aux_osc_en sky130_fd_sc_hs__nand2_4_5/Y
+ sky130_fd_sc_hs__nand2_4_1/a_27_74# sky130_fd_sc_hs__nand2_4
Xsky130_fd_sc_hs__nor3_1_14 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nor3_1_15/Y sky130_fd_sc_hs__inv_4_99/Y
+ sky130_fd_sc_hs__nor3_1_15/B sky130_fd_sc_hs__nor3_1_15/A sky130_fd_sc_hs__nor3_1_15/a_198_368#
+ sky130_fd_sc_hs__nor3_1_15/a_114_368# sky130_fd_sc_hs__nor3_1
Xsky130_fd_sc_hs__nor2_1_103 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__o21a_1_57/B1 sky130_fd_sc_hs__o21a_1_67/A2
+ sky130_fd_sc_hs__nor2_1_95/B sky130_fd_sc_hs__nor2_1_103/a_116_368# sky130_fd_sc_hs__nor2_1
Xsky130_fd_sc_hs__nor2_1_114 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__o21a_1_67/B1 sky130_fd_sc_hs__o21a_1_69/A2
+ sky130_fd_sc_hs__inv_4_125/Y sky130_fd_sc_hs__nor2_1_115/a_116_368# sky130_fd_sc_hs__nor2_1
Xsky130_fd_sc_hs__a22oi_1_23 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nor4_1_3/C sky130_fd_sc_hs__a22oi_1_23/Y
+ sky130_fd_sc_hs__a21oi_1_97/Y sky130_fd_sc_hs__nand2_1_85/Y sky130_fd_sc_hs__nor3_1_5/C
+ sky130_fd_sc_hs__a22oi_1_23/a_71_368# sky130_fd_sc_hs__a22oi_1_23/a_159_74# sky130_fd_sc_hs__a22oi_1_23/a_339_74#
+ sky130_fd_sc_hs__a22oi_1
Xsky130_fd_sc_hs__a22oi_1_12 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nor2_1_33/Y sky130_fd_sc_hs__a22oi_1_13/Y
+ sky130_fd_sc_hs__inv_4_13/A sky130_fd_sc_hs__and2_2_1/X sky130_fd_sc_hs__inv_4_15/A
+ sky130_fd_sc_hs__a22oi_1_13/a_71_368# sky130_fd_sc_hs__a22oi_1_13/a_159_74# sky130_fd_sc_hs__a22oi_1_13/a_339_74#
+ sky130_fd_sc_hs__a22oi_1
Xsky130_fd_sc_hs__nor2_1_91 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nor2_1_91/B sky130_fd_sc_hs__nor2_1_91/Y
+ sky130_fd_sc_hs__xnor2_1_7/Y sky130_fd_sc_hs__nor2_1_91/a_116_368# sky130_fd_sc_hs__nor2_1
Xsky130_fd_sc_hs__nor2_1_80 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_2_3/A sky130_fd_sc_hs__nor2_1_81/Y
+ sky130_fd_sc_hs__or3b_2_1/B sky130_fd_sc_hs__nor2_1_81/a_116_368# sky130_fd_sc_hs__nor2_1
Xsky130_fd_sc_hs__fa_2_19 DVSS DVDD sky130_fd_sc_hs__fa_2_9/B DVDD DVSS sky130_fd_sc_hs__fa_2_19/CIN
+ sky130_fd_sc_hs__fa_2_19/B sky130_fd_sc_hs__fa_2_21/CIN sky130_fd_sc_hs__fa_2_19/SUM
+ sky130_fd_sc_hs__fa_2_19/a_27_378# sky130_fd_sc_hs__fa_2_19/a_701_79# sky130_fd_sc_hs__fa_2_19/a_484_347#
+ sky130_fd_sc_hs__fa_2_19/a_1094_347# sky130_fd_sc_hs__fa_2_19/a_1205_79# sky130_fd_sc_hs__fa_2_19/a_27_79#
+ sky130_fd_sc_hs__fa_2_19/a_1202_368# sky130_fd_sc_hs__fa_2_19/a_336_347# sky130_fd_sc_hs__fa_2_19/a_992_347#
+ sky130_fd_sc_hs__fa_2_19/a_1119_79# sky130_fd_sc_hs__fa_2_19/a_487_79# sky130_fd_sc_hs__fa_2_19/a_683_347#
+ sky130_fd_sc_hs__fa_2
Xsky130_fd_sc_hs__xnor2_1_0 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__xnor2_1_1/A sky130_fd_sc_hs__xnor2_1_1/Y
+ sky130_fd_sc_hs__xnor2_1_1/B sky130_fd_sc_hs__xnor2_1_1/a_376_368# sky130_fd_sc_hs__xnor2_1_1/a_112_119#
+ sky130_fd_sc_hs__xnor2_1_1/a_138_385# sky130_fd_sc_hs__xnor2_1_1/a_293_74# sky130_fd_sc_hs__xnor2_1
Xsky130_fd_sc_hs__o21a_1_15 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__o21a_1_15/X sky130_fd_sc_hs__nor2_1_7/Y
+ sky130_fd_sc_hs__nor2_1_35/B sky130_fd_sc_hs__o21a_1_15/A1 sky130_fd_sc_hs__o21a_1_15/a_320_74#
+ sky130_fd_sc_hs__o21a_1_15/a_376_387# sky130_fd_sc_hs__o21a_1_15/a_83_244# sky130_fd_sc_hs__o21a_1
Xsky130_fd_sc_hs__o21a_1_48 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__o21a_1_49/X sky130_fd_sc_hs__nor2_1_87/Y
+ sky130_fd_sc_hs__nor2_1_45/B sky130_fd_sc_hs__inv_4_83/A sky130_fd_sc_hs__o21a_1_49/a_320_74#
+ sky130_fd_sc_hs__o21a_1_49/a_376_387# sky130_fd_sc_hs__o21a_1_49/a_83_244# sky130_fd_sc_hs__o21a_1
Xsky130_fd_sc_hs__o21a_1_37 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__o21a_1_37/X sky130_fd_sc_hs__nor2_1_45/Y
+ sky130_fd_sc_hs__nor2_1_29/B sky130_fd_sc_hs__nor2_1_65/A sky130_fd_sc_hs__o21a_1_37/a_320_74#
+ sky130_fd_sc_hs__o21a_1_37/a_376_387# sky130_fd_sc_hs__o21a_1_37/a_83_244# sky130_fd_sc_hs__o21a_1
Xsky130_fd_sc_hs__o21a_1_26 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__o21a_1_27/X sky130_fd_sc_hs__nor2_1_31/Y
+ sky130_fd_sc_hs__nor2_1_21/B sky130_fd_sc_hs__o21a_1_27/A1 sky130_fd_sc_hs__o21a_1_27/a_320_74#
+ sky130_fd_sc_hs__o21a_1_27/a_376_387# sky130_fd_sc_hs__o21a_1_27/a_83_244# sky130_fd_sc_hs__o21a_1
Xsky130_fd_sc_hs__o21a_1_59 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__o21a_1_59/X sky130_fd_sc_hs__o21a_1_59/A2
+ sky130_fd_sc_hs__nor2_1_87/B sky130_fd_sc_hs__o21a_1_59/A1 sky130_fd_sc_hs__o21a_1_59/a_320_74#
+ sky130_fd_sc_hs__o21a_1_59/a_376_387# sky130_fd_sc_hs__o21a_1_59/a_83_244# sky130_fd_sc_hs__o21a_1
Xsky130_fd_sc_hs__dfrtp_4_16 DVSS DVDD sky130_fd_sc_hs__clkbuf_8_1/X DVDD DVSS sky130_fd_sc_hs__o21a_1_7/X
+ sky130_fd_sc_hs__nand2_1_47/B sky130_fd_sc_hs__o21a_1_7/A1 sky130_fd_sc_hs__dfrtp_4_17/a_37_78#
+ sky130_fd_sc_hs__dfrtp_4_17/a_494_366# sky130_fd_sc_hs__dfrtp_4_17/a_699_463# sky130_fd_sc_hs__dfrtp_4_17/a_313_74#
+ sky130_fd_sc_hs__dfrtp_4_17/a_1627_493# sky130_fd_sc_hs__dfrtp_4_17/a_1678_395#
+ sky130_fd_sc_hs__dfrtp_4_17/a_1827_81# sky130_fd_sc_hs__dfrtp_4_17/a_789_463# sky130_fd_sc_hs__dfrtp_4_17/a_1350_392#
+ sky130_fd_sc_hs__dfrtp_4_17/a_834_355# sky130_fd_sc_hs__dfrtp_4_17/a_812_138# sky130_fd_sc_hs__dfrtp_4_17/a_124_78#
+ sky130_fd_sc_hs__dfrtp_4_17/a_1647_81# sky130_fd_sc_hs__dfrtp_4_17/a_2010_409# sky130_fd_sc_hs__dfrtp_4_17/a_890_138#
+ sky130_fd_sc_hs__dfrtp_4
Xsky130_fd_sc_hs__dfrtp_4_49 DVSS DVDD sky130_fd_sc_hs__clkbuf_8_1/X DVDD DVSS sky130_fd_sc_hs__o21a_1_21/X
+ sky130_fd_sc_hs__nand2_1_47/B sky130_fd_sc_hs__o21a_1_21/A1 sky130_fd_sc_hs__dfrtp_4_49/a_37_78#
+ sky130_fd_sc_hs__dfrtp_4_49/a_494_366# sky130_fd_sc_hs__dfrtp_4_49/a_699_463# sky130_fd_sc_hs__dfrtp_4_49/a_313_74#
+ sky130_fd_sc_hs__dfrtp_4_49/a_1627_493# sky130_fd_sc_hs__dfrtp_4_49/a_1678_395#
+ sky130_fd_sc_hs__dfrtp_4_49/a_1827_81# sky130_fd_sc_hs__dfrtp_4_49/a_789_463# sky130_fd_sc_hs__dfrtp_4_49/a_1350_392#
+ sky130_fd_sc_hs__dfrtp_4_49/a_834_355# sky130_fd_sc_hs__dfrtp_4_49/a_812_138# sky130_fd_sc_hs__dfrtp_4_49/a_124_78#
+ sky130_fd_sc_hs__dfrtp_4_49/a_1647_81# sky130_fd_sc_hs__dfrtp_4_49/a_2010_409# sky130_fd_sc_hs__dfrtp_4_49/a_890_138#
+ sky130_fd_sc_hs__dfrtp_4
Xsky130_fd_sc_hs__dfrtp_4_38 DVSS DVDD sky130_fd_sc_hs__clkbuf_8_1/X DVDD DVSS sky130_fd_sc_hs__o21a_1_15/X
+ sky130_fd_sc_hs__nand2_1_47/B sky130_fd_sc_hs__o21a_1_15/A1 sky130_fd_sc_hs__dfrtp_4_39/a_37_78#
+ sky130_fd_sc_hs__dfrtp_4_39/a_494_366# sky130_fd_sc_hs__dfrtp_4_39/a_699_463# sky130_fd_sc_hs__dfrtp_4_39/a_313_74#
+ sky130_fd_sc_hs__dfrtp_4_39/a_1627_493# sky130_fd_sc_hs__dfrtp_4_39/a_1678_395#
+ sky130_fd_sc_hs__dfrtp_4_39/a_1827_81# sky130_fd_sc_hs__dfrtp_4_39/a_789_463# sky130_fd_sc_hs__dfrtp_4_39/a_1350_392#
+ sky130_fd_sc_hs__dfrtp_4_39/a_834_355# sky130_fd_sc_hs__dfrtp_4_39/a_812_138# sky130_fd_sc_hs__dfrtp_4_39/a_124_78#
+ sky130_fd_sc_hs__dfrtp_4_39/a_1647_81# sky130_fd_sc_hs__dfrtp_4_39/a_2010_409# sky130_fd_sc_hs__dfrtp_4_39/a_890_138#
+ sky130_fd_sc_hs__dfrtp_4
Xsky130_fd_sc_hs__dfrtp_4_27 DVSS DVDD sky130_fd_sc_hs__clkbuf_8_1/A DVDD DVSS sky130_fd_sc_hs__o21a_1_9/X
+ sky130_fd_sc_hs__nand2_1_47/B sky130_fd_sc_hs__o21a_1_9/A1 sky130_fd_sc_hs__dfrtp_4_27/a_37_78#
+ sky130_fd_sc_hs__dfrtp_4_27/a_494_366# sky130_fd_sc_hs__dfrtp_4_27/a_699_463# sky130_fd_sc_hs__dfrtp_4_27/a_313_74#
+ sky130_fd_sc_hs__dfrtp_4_27/a_1627_493# sky130_fd_sc_hs__dfrtp_4_27/a_1678_395#
+ sky130_fd_sc_hs__dfrtp_4_27/a_1827_81# sky130_fd_sc_hs__dfrtp_4_27/a_789_463# sky130_fd_sc_hs__dfrtp_4_27/a_1350_392#
+ sky130_fd_sc_hs__dfrtp_4_27/a_834_355# sky130_fd_sc_hs__dfrtp_4_27/a_812_138# sky130_fd_sc_hs__dfrtp_4_27/a_124_78#
+ sky130_fd_sc_hs__dfrtp_4_27/a_1647_81# sky130_fd_sc_hs__dfrtp_4_27/a_2010_409# sky130_fd_sc_hs__dfrtp_4_27/a_890_138#
+ sky130_fd_sc_hs__dfrtp_4
Xsky130_fd_sc_hs__inv_4_1 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_1/Y sky130_fd_sc_hs__inv_4_1/A
+ sky130_fd_sc_hs__inv_4
Xsky130_fd_sc_hs__nand4_1_1 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand4_1_1/C sky130_fd_sc_hs__nand4_1_1/Y
+ sky130_fd_sc_hs__nand4_1_1/D sky130_fd_sc_hs__nor3_1_9/Y sky130_fd_sc_hs__nor3_1_1/Y
+ sky130_fd_sc_hs__nand4_1_1/a_259_74# sky130_fd_sc_hs__nand4_1_1/a_373_74# sky130_fd_sc_hs__nand4_1_1/a_181_74#
+ sky130_fd_sc_hs__nand4_1
Xsky130_fd_sc_hs__nand2_1_51 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_53/Y sky130_fd_sc_hs__nand2_1_51/Y
+ sky130_fd_sc_hs__inv_4_51/A sky130_fd_sc_hs__nand2_1_51/a_117_74# sky130_fd_sc_hs__nand2_1
Xsky130_fd_sc_hs__nand2_1_40 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nor2_1_41/Y sky130_fd_sc_hs__nor2_1_51/B
+ sky130_fd_sc_hs__dfrbp_1_1/Q sky130_fd_sc_hs__nand2_1_41/a_117_74# sky130_fd_sc_hs__nand2_1
Xsky130_fd_sc_hs__nand2_1_84 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__or2_1_3/B sky130_fd_sc_hs__nand2_1_85/Y
+ sky130_fd_sc_hs__or2_1_3/A sky130_fd_sc_hs__nand2_1_85/a_117_74# sky130_fd_sc_hs__nand2_1
Xsky130_fd_sc_hs__nand2_1_73 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nor2_1_73/Y sky130_fd_sc_hs__o21a_1_53/B1
+ sky130_fd_sc_hs__o22ai_1_7/A1 sky130_fd_sc_hs__nand2_1_73/a_117_74# sky130_fd_sc_hs__nand2_1
Xsky130_fd_sc_hs__nand2_1_62 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nor2_1_57/Y sky130_fd_sc_hs__nor2_1_83/B
+ sky130_fd_sc_hs__inv_4_69/A sky130_fd_sc_hs__nand2_1_63/a_117_74# sky130_fd_sc_hs__nand2_1
Xsky130_fd_sc_hs__nand2_1_95 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_129/Y sky130_fd_sc_hs__nand4_1_5/D
+ sky130_fd_sc_hs__inv_4_137/A sky130_fd_sc_hs__nand2_1_95/a_117_74# sky130_fd_sc_hs__nand2_1
Xsky130_fd_sc_hs__a21oi_1_19 DVSS DVDD DVDD DVSS fine_control_avg_window_select[2]
+ sky130_fd_sc_hs__a21oi_1_19/Y sky130_fd_sc_hs__a22oi_1_1/Y sky130_fd_sc_hs__a22oi_1_5/Y
+ sky130_fd_sc_hs__a21oi_1_19/a_117_74# sky130_fd_sc_hs__a21oi_1_19/a_29_368# sky130_fd_sc_hs__a21oi_1
Xsky130_fd_sc_hs__nand2_4_2 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_4_7/A aux_osc_en
+ aux_clk_out sky130_fd_sc_hs__nand2_4_3/a_27_74# sky130_fd_sc_hs__nand2_4
Xsky130_fd_sc_hs__nor3_1_15 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nor3_1_15/Y sky130_fd_sc_hs__inv_4_99/Y
+ sky130_fd_sc_hs__nor3_1_15/B sky130_fd_sc_hs__nor3_1_15/A sky130_fd_sc_hs__nor3_1_15/a_198_368#
+ sky130_fd_sc_hs__nor3_1_15/a_114_368# sky130_fd_sc_hs__nor3_1
Xsky130_fd_sc_hs__nor2_1_104 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__o21a_1_51/B1 sky130_fd_sc_hs__o21a_1_75/A2
+ sky130_fd_sc_hs__inv_4_107/Y sky130_fd_sc_hs__nor2_1_105/a_116_368# sky130_fd_sc_hs__nor2_1
Xsky130_fd_sc_hs__nor2_1_115 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__o21a_1_67/B1 sky130_fd_sc_hs__o21a_1_69/A2
+ sky130_fd_sc_hs__inv_4_125/Y sky130_fd_sc_hs__nor2_1_115/a_116_368# sky130_fd_sc_hs__nor2_1
Xsky130_fd_sc_hs__a22oi_1_24 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__maj3_1_3/B sky130_fd_sc_hs__inv_4_109/A
+ sky130_fd_sc_hs__maj3_1_3/A sky130_fd_sc_hs__inv_4_125/Y sky130_fd_sc_hs__inv_4_135/A
+ sky130_fd_sc_hs__a22oi_1_25/a_71_368# sky130_fd_sc_hs__a22oi_1_25/a_159_74# sky130_fd_sc_hs__a22oi_1_25/a_339_74#
+ sky130_fd_sc_hs__a22oi_1
Xsky130_fd_sc_hs__a22oi_1_13 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nor2_1_33/Y sky130_fd_sc_hs__a22oi_1_13/Y
+ sky130_fd_sc_hs__inv_4_13/A sky130_fd_sc_hs__and2_2_1/X sky130_fd_sc_hs__inv_4_15/A
+ sky130_fd_sc_hs__a22oi_1_13/a_71_368# sky130_fd_sc_hs__a22oi_1_13/a_159_74# sky130_fd_sc_hs__a22oi_1_13/a_339_74#
+ sky130_fd_sc_hs__a22oi_1
Xsky130_fd_sc_hs__nor2_1_92 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_99/Y sky130_fd_sc_hs__nor3_1_13/B
+ sky130_fd_sc_hs__nor3_1_15/A sky130_fd_sc_hs__nor2_1_93/a_116_368# sky130_fd_sc_hs__nor2_1
Xsky130_fd_sc_hs__nor2_1_81 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_2_3/A sky130_fd_sc_hs__nor2_1_81/Y
+ sky130_fd_sc_hs__or3b_2_1/B sky130_fd_sc_hs__nor2_1_81/a_116_368# sky130_fd_sc_hs__nor2_1
Xsky130_fd_sc_hs__nor2_1_70 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_63/Y sky130_fd_sc_hs__nor3_1_5/A
+ sky130_fd_sc_hs__inv_4_67/A sky130_fd_sc_hs__nor2_1_71/a_116_368# sky130_fd_sc_hs__nor2_1
Xsky130_fd_sc_hs__xnor2_1_1 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__xnor2_1_1/A sky130_fd_sc_hs__xnor2_1_1/Y
+ sky130_fd_sc_hs__xnor2_1_1/B sky130_fd_sc_hs__xnor2_1_1/a_376_368# sky130_fd_sc_hs__xnor2_1_1/a_112_119#
+ sky130_fd_sc_hs__xnor2_1_1/a_138_385# sky130_fd_sc_hs__xnor2_1_1/a_293_74# sky130_fd_sc_hs__xnor2_1
Xsky130_fd_sc_hs__or2_1_0 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__or2_1_1/B sky130_fd_sc_hs__or2_1_1/A
+ sky130_fd_sc_hs__or2_1_1/X sky130_fd_sc_hs__or2_1_1/a_152_368# sky130_fd_sc_hs__or2_1_1/a_63_368#
+ sky130_fd_sc_hs__or2_1
Xsky130_fd_sc_hs__o21a_1_49 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__o21a_1_49/X sky130_fd_sc_hs__nor2_1_87/Y
+ sky130_fd_sc_hs__nor2_1_45/B sky130_fd_sc_hs__inv_4_83/A sky130_fd_sc_hs__o21a_1_49/a_320_74#
+ sky130_fd_sc_hs__o21a_1_49/a_376_387# sky130_fd_sc_hs__o21a_1_49/a_83_244# sky130_fd_sc_hs__o21a_1
Xsky130_fd_sc_hs__o21a_1_38 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__o21a_1_39/X sky130_fd_sc_hs__nor2_1_49/Y
+ sky130_fd_sc_hs__nor2_1_47/B sky130_fd_sc_hs__nor2_1_69/B sky130_fd_sc_hs__o21a_1_39/a_320_74#
+ sky130_fd_sc_hs__o21a_1_39/a_376_387# sky130_fd_sc_hs__o21a_1_39/a_83_244# sky130_fd_sc_hs__o21a_1
Xsky130_fd_sc_hs__o21a_1_27 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__o21a_1_27/X sky130_fd_sc_hs__nor2_1_31/Y
+ sky130_fd_sc_hs__nor2_1_21/B sky130_fd_sc_hs__o21a_1_27/A1 sky130_fd_sc_hs__o21a_1_27/a_320_74#
+ sky130_fd_sc_hs__o21a_1_27/a_376_387# sky130_fd_sc_hs__o21a_1_27/a_83_244# sky130_fd_sc_hs__o21a_1
Xsky130_fd_sc_hs__o21a_1_16 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__o21a_1_17/X sky130_fd_sc_hs__nor2_1_21/Y
+ sky130_fd_sc_hs__nor2_1_15/B sky130_fd_sc_hs__o21a_1_17/A1 sky130_fd_sc_hs__o21a_1_17/a_320_74#
+ sky130_fd_sc_hs__o21a_1_17/a_376_387# sky130_fd_sc_hs__o21a_1_17/a_83_244# sky130_fd_sc_hs__o21a_1
Xsky130_fd_sc_hs__dfrtp_4_39 DVSS DVDD sky130_fd_sc_hs__clkbuf_8_1/X DVDD DVSS sky130_fd_sc_hs__o21a_1_15/X
+ sky130_fd_sc_hs__nand2_1_47/B sky130_fd_sc_hs__o21a_1_15/A1 sky130_fd_sc_hs__dfrtp_4_39/a_37_78#
+ sky130_fd_sc_hs__dfrtp_4_39/a_494_366# sky130_fd_sc_hs__dfrtp_4_39/a_699_463# sky130_fd_sc_hs__dfrtp_4_39/a_313_74#
+ sky130_fd_sc_hs__dfrtp_4_39/a_1627_493# sky130_fd_sc_hs__dfrtp_4_39/a_1678_395#
+ sky130_fd_sc_hs__dfrtp_4_39/a_1827_81# sky130_fd_sc_hs__dfrtp_4_39/a_789_463# sky130_fd_sc_hs__dfrtp_4_39/a_1350_392#
+ sky130_fd_sc_hs__dfrtp_4_39/a_834_355# sky130_fd_sc_hs__dfrtp_4_39/a_812_138# sky130_fd_sc_hs__dfrtp_4_39/a_124_78#
+ sky130_fd_sc_hs__dfrtp_4_39/a_1647_81# sky130_fd_sc_hs__dfrtp_4_39/a_2010_409# sky130_fd_sc_hs__dfrtp_4_39/a_890_138#
+ sky130_fd_sc_hs__dfrtp_4
Xsky130_fd_sc_hs__dfrtp_4_28 DVSS DVDD sky130_fd_sc_hs__inv_4_49/Y DVDD DVSS sky130_fd_sc_hs__nor2b_1_7/Y
+ sky130_fd_sc_hs__dfstp_2_1/CLK sky130_fd_sc_hs__fa_2_7/B sky130_fd_sc_hs__dfrtp_4_29/a_37_78#
+ sky130_fd_sc_hs__dfrtp_4_29/a_494_366# sky130_fd_sc_hs__dfrtp_4_29/a_699_463# sky130_fd_sc_hs__dfrtp_4_29/a_313_74#
+ sky130_fd_sc_hs__dfrtp_4_29/a_1627_493# sky130_fd_sc_hs__dfrtp_4_29/a_1678_395#
+ sky130_fd_sc_hs__dfrtp_4_29/a_1827_81# sky130_fd_sc_hs__dfrtp_4_29/a_789_463# sky130_fd_sc_hs__dfrtp_4_29/a_1350_392#
+ sky130_fd_sc_hs__dfrtp_4_29/a_834_355# sky130_fd_sc_hs__dfrtp_4_29/a_812_138# sky130_fd_sc_hs__dfrtp_4_29/a_124_78#
+ sky130_fd_sc_hs__dfrtp_4_29/a_1647_81# sky130_fd_sc_hs__dfrtp_4_29/a_2010_409# sky130_fd_sc_hs__dfrtp_4_29/a_890_138#
+ sky130_fd_sc_hs__dfrtp_4
Xsky130_fd_sc_hs__dfrtp_4_17 DVSS DVDD sky130_fd_sc_hs__clkbuf_8_1/X DVDD DVSS sky130_fd_sc_hs__o21a_1_7/X
+ sky130_fd_sc_hs__nand2_1_47/B sky130_fd_sc_hs__o21a_1_7/A1 sky130_fd_sc_hs__dfrtp_4_17/a_37_78#
+ sky130_fd_sc_hs__dfrtp_4_17/a_494_366# sky130_fd_sc_hs__dfrtp_4_17/a_699_463# sky130_fd_sc_hs__dfrtp_4_17/a_313_74#
+ sky130_fd_sc_hs__dfrtp_4_17/a_1627_493# sky130_fd_sc_hs__dfrtp_4_17/a_1678_395#
+ sky130_fd_sc_hs__dfrtp_4_17/a_1827_81# sky130_fd_sc_hs__dfrtp_4_17/a_789_463# sky130_fd_sc_hs__dfrtp_4_17/a_1350_392#
+ sky130_fd_sc_hs__dfrtp_4_17/a_834_355# sky130_fd_sc_hs__dfrtp_4_17/a_812_138# sky130_fd_sc_hs__dfrtp_4_17/a_124_78#
+ sky130_fd_sc_hs__dfrtp_4_17/a_1647_81# sky130_fd_sc_hs__dfrtp_4_17/a_2010_409# sky130_fd_sc_hs__dfrtp_4_17/a_890_138#
+ sky130_fd_sc_hs__dfrtp_4
Xsky130_fd_sc_hs__inv_4_2 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_3/Y sky130_fd_sc_hs__inv_4_3/A
+ sky130_fd_sc_hs__inv_4
Xsky130_fd_sc_hs__nand4_1_2 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nor4_1_3/Y sky130_fd_sc_hs__nor3_1_3/B
+ sky130_fd_sc_hs__or2_1_3/X sky130_fd_sc_hs__nor3_1_5/Y sky130_fd_sc_hs__nor4_1_1/Y
+ sky130_fd_sc_hs__nand4_1_3/a_259_74# sky130_fd_sc_hs__nand4_1_3/a_373_74# sky130_fd_sc_hs__nand4_1_3/a_181_74#
+ sky130_fd_sc_hs__nand4_1
Xsky130_fd_sc_hs__nand2_1_41 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nor2_1_41/Y sky130_fd_sc_hs__nor2_1_51/B
+ sky130_fd_sc_hs__dfrbp_1_1/Q sky130_fd_sc_hs__nand2_1_41/a_117_74# sky130_fd_sc_hs__nand2_1
Xsky130_fd_sc_hs__nand2_1_30 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nor2_1_17/Y sky130_fd_sc_hs__xnor2_1_1/B
+ sky130_fd_sc_hs__o21a_1_23/A1 sky130_fd_sc_hs__nand2_1_31/a_117_74# sky130_fd_sc_hs__nand2_1
Xsky130_fd_sc_hs__nand2_1_85 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__or2_1_3/B sky130_fd_sc_hs__nand2_1_85/Y
+ sky130_fd_sc_hs__or2_1_3/A sky130_fd_sc_hs__nand2_1_85/a_117_74# sky130_fd_sc_hs__nand2_1
Xsky130_fd_sc_hs__nand2_1_74 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nor2_1_83/Y sky130_fd_sc_hs__o21a_1_51/B1
+ sky130_fd_sc_hs__maj3_1_1/A sky130_fd_sc_hs__nand2_1_75/a_117_74# sky130_fd_sc_hs__nand2_1
Xsky130_fd_sc_hs__nand2_1_63 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nor2_1_57/Y sky130_fd_sc_hs__nor2_1_83/B
+ sky130_fd_sc_hs__inv_4_69/A sky130_fd_sc_hs__nand2_1_63/a_117_74# sky130_fd_sc_hs__nand2_1
Xsky130_fd_sc_hs__nand2_1_52 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nor2_1_43/Y sky130_fd_sc_hs__nor2_1_41/B
+ sky130_fd_sc_hs__inv_4_73/A sky130_fd_sc_hs__nand2_1_53/a_117_74# sky130_fd_sc_hs__nand2_1
Xsky130_fd_sc_hs__nand2_1_96 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nor2_1_99/Y sky130_fd_sc_hs__o21a_1_65/B1
+ sky130_fd_sc_hs__inv_4_101/A sky130_fd_sc_hs__nand2_1_97/a_117_74# sky130_fd_sc_hs__nand2_1
Xsky130_fd_sc_hs__nand2_4_3 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_4_7/A aux_osc_en
+ aux_clk_out sky130_fd_sc_hs__nand2_4_3/a_27_74# sky130_fd_sc_hs__nand2_4
Xsky130_fd_sc_hs__nand2_2_0 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_2_1/Y sky130_fd_sc_hs__nand2_2_1/B
+ sky130_fd_sc_hs__nand2_2_1/A sky130_fd_sc_hs__nand2_2_1/a_27_74# sky130_fd_sc_hs__nand2_2
Xsky130_fd_sc_hs__nor2_1_105 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__o21a_1_51/B1 sky130_fd_sc_hs__o21a_1_75/A2
+ sky130_fd_sc_hs__inv_4_107/Y sky130_fd_sc_hs__nor2_1_105/a_116_368# sky130_fd_sc_hs__nor2_1
Xsky130_fd_sc_hs__nor2_1_116 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_133/Y sky130_fd_sc_hs__nor3_1_9/C
+ sky130_fd_sc_hs__o21a_1_75/A1 sky130_fd_sc_hs__nor2_1_117/a_116_368# sky130_fd_sc_hs__nor2_1
Xsky130_fd_sc_hs__a22oi_1_25 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__maj3_1_3/B sky130_fd_sc_hs__inv_4_109/A
+ sky130_fd_sc_hs__maj3_1_3/A sky130_fd_sc_hs__inv_4_125/Y sky130_fd_sc_hs__inv_4_135/A
+ sky130_fd_sc_hs__a22oi_1_25/a_71_368# sky130_fd_sc_hs__a22oi_1_25/a_159_74# sky130_fd_sc_hs__a22oi_1_25/a_339_74#
+ sky130_fd_sc_hs__a22oi_1
Xsky130_fd_sc_hs__a22oi_1_14 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nor2_1_33/Y sky130_fd_sc_hs__a22oi_1_15/Y
+ sky130_fd_sc_hs__o21a_1_13/A1 sky130_fd_sc_hs__nor2b_1_25/Y sky130_fd_sc_hs__o21a_1_21/A1
+ sky130_fd_sc_hs__a22oi_1_15/a_71_368# sky130_fd_sc_hs__a22oi_1_15/a_159_74# sky130_fd_sc_hs__a22oi_1_15/a_339_74#
+ sky130_fd_sc_hs__a22oi_1
Xsky130_fd_sc_hs__nor2_1_82 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nor2_1_83/B sky130_fd_sc_hs__nor2_1_83/Y
+ sky130_fd_sc_hs__inv_4_89/Y sky130_fd_sc_hs__nor2_1_83/a_116_368# sky130_fd_sc_hs__nor2_1
Xsky130_fd_sc_hs__nor2_1_71 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_63/Y sky130_fd_sc_hs__nor3_1_5/A
+ sky130_fd_sc_hs__inv_4_67/A sky130_fd_sc_hs__nor2_1_71/a_116_368# sky130_fd_sc_hs__nor2_1
Xsky130_fd_sc_hs__nor2_1_60 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nor2_1_61/B sky130_fd_sc_hs__nor2_1_61/Y
+ sky130_fd_sc_hs__o22ai_1_3/Y sky130_fd_sc_hs__nor2_1_61/a_116_368# sky130_fd_sc_hs__nor2_1
Xsky130_fd_sc_hs__nor2_1_93 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_99/Y sky130_fd_sc_hs__nor3_1_13/B
+ sky130_fd_sc_hs__nor3_1_15/A sky130_fd_sc_hs__nor2_1_93/a_116_368# sky130_fd_sc_hs__nor2_1
Xsky130_fd_sc_hs__xnor2_1_2 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__xnor2_1_3/A sky130_fd_sc_hs__xnor2_1_3/Y
+ sky130_fd_sc_hs__xnor2_1_3/B sky130_fd_sc_hs__xnor2_1_3/a_376_368# sky130_fd_sc_hs__xnor2_1_3/a_112_119#
+ sky130_fd_sc_hs__xnor2_1_3/a_138_385# sky130_fd_sc_hs__xnor2_1_3/a_293_74# sky130_fd_sc_hs__xnor2_1
Xsky130_fd_sc_hs__inv_4_130 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_2_7/B div_ratio_half[2]
+ sky130_fd_sc_hs__inv_4
Xsky130_fd_sc_hs__or2_1_1 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__or2_1_1/B sky130_fd_sc_hs__or2_1_1/A
+ sky130_fd_sc_hs__or2_1_1/X sky130_fd_sc_hs__or2_1_1/a_152_368# sky130_fd_sc_hs__or2_1_1/a_63_368#
+ sky130_fd_sc_hs__or2_1
Xsky130_fd_sc_hs__o21a_1_39 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__o21a_1_39/X sky130_fd_sc_hs__nor2_1_49/Y
+ sky130_fd_sc_hs__nor2_1_47/B sky130_fd_sc_hs__nor2_1_69/B sky130_fd_sc_hs__o21a_1_39/a_320_74#
+ sky130_fd_sc_hs__o21a_1_39/a_376_387# sky130_fd_sc_hs__o21a_1_39/a_83_244# sky130_fd_sc_hs__o21a_1
Xsky130_fd_sc_hs__o21a_1_28 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__o21a_1_29/X sky130_fd_sc_hs__nor2_1_29/Y
+ sky130_fd_sc_hs__nor2_1_27/B sky130_fd_sc_hs__inv_4_39/A sky130_fd_sc_hs__o21a_1_29/a_320_74#
+ sky130_fd_sc_hs__o21a_1_29/a_376_387# sky130_fd_sc_hs__o21a_1_29/a_83_244# sky130_fd_sc_hs__o21a_1
Xsky130_fd_sc_hs__o21a_1_17 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__o21a_1_17/X sky130_fd_sc_hs__nor2_1_21/Y
+ sky130_fd_sc_hs__nor2_1_15/B sky130_fd_sc_hs__o21a_1_17/A1 sky130_fd_sc_hs__o21a_1_17/a_320_74#
+ sky130_fd_sc_hs__o21a_1_17/a_376_387# sky130_fd_sc_hs__o21a_1_17/a_83_244# sky130_fd_sc_hs__o21a_1
Xsky130_fd_sc_hs__dfrtp_4_29 DVSS DVDD sky130_fd_sc_hs__inv_4_49/Y DVDD DVSS sky130_fd_sc_hs__nor2b_1_7/Y
+ sky130_fd_sc_hs__dfstp_2_1/CLK sky130_fd_sc_hs__fa_2_7/B sky130_fd_sc_hs__dfrtp_4_29/a_37_78#
+ sky130_fd_sc_hs__dfrtp_4_29/a_494_366# sky130_fd_sc_hs__dfrtp_4_29/a_699_463# sky130_fd_sc_hs__dfrtp_4_29/a_313_74#
+ sky130_fd_sc_hs__dfrtp_4_29/a_1627_493# sky130_fd_sc_hs__dfrtp_4_29/a_1678_395#
+ sky130_fd_sc_hs__dfrtp_4_29/a_1827_81# sky130_fd_sc_hs__dfrtp_4_29/a_789_463# sky130_fd_sc_hs__dfrtp_4_29/a_1350_392#
+ sky130_fd_sc_hs__dfrtp_4_29/a_834_355# sky130_fd_sc_hs__dfrtp_4_29/a_812_138# sky130_fd_sc_hs__dfrtp_4_29/a_124_78#
+ sky130_fd_sc_hs__dfrtp_4_29/a_1647_81# sky130_fd_sc_hs__dfrtp_4_29/a_2010_409# sky130_fd_sc_hs__dfrtp_4_29/a_890_138#
+ sky130_fd_sc_hs__dfrtp_4
Xsky130_fd_sc_hs__dfrtp_4_18 DVSS DVDD sky130_fd_sc_hs__inv_4_49/Y DVDD DVSS sky130_fd_sc_hs__nor2b_1_3/Y
+ sky130_fd_sc_hs__dfstp_2_1/CLK sky130_fd_sc_hs__fa_2_3/B sky130_fd_sc_hs__dfrtp_4_19/a_37_78#
+ sky130_fd_sc_hs__dfrtp_4_19/a_494_366# sky130_fd_sc_hs__dfrtp_4_19/a_699_463# sky130_fd_sc_hs__dfrtp_4_19/a_313_74#
+ sky130_fd_sc_hs__dfrtp_4_19/a_1627_493# sky130_fd_sc_hs__dfrtp_4_19/a_1678_395#
+ sky130_fd_sc_hs__dfrtp_4_19/a_1827_81# sky130_fd_sc_hs__dfrtp_4_19/a_789_463# sky130_fd_sc_hs__dfrtp_4_19/a_1350_392#
+ sky130_fd_sc_hs__dfrtp_4_19/a_834_355# sky130_fd_sc_hs__dfrtp_4_19/a_812_138# sky130_fd_sc_hs__dfrtp_4_19/a_124_78#
+ sky130_fd_sc_hs__dfrtp_4_19/a_1647_81# sky130_fd_sc_hs__dfrtp_4_19/a_2010_409# sky130_fd_sc_hs__dfrtp_4_19/a_890_138#
+ sky130_fd_sc_hs__dfrtp_4
Xsky130_fd_sc_hs__inv_4_3 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_3/Y sky130_fd_sc_hs__inv_4_3/A
+ sky130_fd_sc_hs__inv_4
Xsky130_fd_sc_hs__a22o_1_20 DVSS DVDD DVDD DVSS osc_fine_con_final[8] manual_control_osc[8]
+ sky130_fd_sc_hs__inv_4_43/Y sky130_fd_sc_hs__fa_2_19/B fftl_en sky130_fd_sc_hs__a22o_1_21/a_222_392#
+ sky130_fd_sc_hs__a22o_1_21/a_230_79# sky130_fd_sc_hs__a22o_1_21/a_52_123# sky130_fd_sc_hs__a22o_1_21/a_132_392#
+ sky130_fd_sc_hs__a22o_1
Xsky130_fd_sc_hs__nand4_1_3 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nor4_1_3/Y sky130_fd_sc_hs__nor3_1_3/B
+ sky130_fd_sc_hs__or2_1_3/X sky130_fd_sc_hs__nor3_1_5/Y sky130_fd_sc_hs__nor4_1_1/Y
+ sky130_fd_sc_hs__nand4_1_3/a_259_74# sky130_fd_sc_hs__nand4_1_3/a_373_74# sky130_fd_sc_hs__nand4_1_3/a_181_74#
+ sky130_fd_sc_hs__nand4_1
Xsky130_fd_sc_hs__nand2_1_42 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nor2_1_45/Y sky130_fd_sc_hs__nor2_1_29/B
+ sky130_fd_sc_hs__nor2_1_65/A sky130_fd_sc_hs__nand2_1_43/a_117_74# sky130_fd_sc_hs__nand2_1
Xsky130_fd_sc_hs__nand2_1_31 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nor2_1_17/Y sky130_fd_sc_hs__xnor2_1_1/B
+ sky130_fd_sc_hs__o21a_1_23/A1 sky130_fd_sc_hs__nand2_1_31/a_117_74# sky130_fd_sc_hs__nand2_1
Xsky130_fd_sc_hs__nand2_1_20 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nor2_1_37/Y sky130_fd_sc_hs__nor2_1_9/B
+ sky130_fd_sc_hs__o21a_1_19/A1 sky130_fd_sc_hs__nand2_1_21/a_117_74# sky130_fd_sc_hs__nand2_1
Xsky130_fd_sc_hs__nand2_1_75 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nor2_1_83/Y sky130_fd_sc_hs__o21a_1_51/B1
+ sky130_fd_sc_hs__maj3_1_1/A sky130_fd_sc_hs__nand2_1_75/a_117_74# sky130_fd_sc_hs__nand2_1
Xsky130_fd_sc_hs__nand2_1_64 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nor2_1_51/Y sky130_fd_sc_hs__nor2_1_57/B
+ sky130_fd_sc_hs__nor2_1_59/A sky130_fd_sc_hs__nand2_1_65/a_117_74# sky130_fd_sc_hs__nand2_1
Xsky130_fd_sc_hs__nand2_1_53 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nor2_1_43/Y sky130_fd_sc_hs__nor2_1_41/B
+ sky130_fd_sc_hs__inv_4_73/A sky130_fd_sc_hs__nand2_1_53/a_117_74# sky130_fd_sc_hs__nand2_1
Xsky130_fd_sc_hs__nand2_1_97 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nor2_1_99/Y sky130_fd_sc_hs__o21a_1_65/B1
+ sky130_fd_sc_hs__inv_4_101/A sky130_fd_sc_hs__nand2_1_97/a_117_74# sky130_fd_sc_hs__nand2_1
Xsky130_fd_sc_hs__nand2_1_86 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nor2_1_75/Y sky130_fd_sc_hs__nor2_1_99/B
+ sky130_fd_sc_hs__inv_4_97/A sky130_fd_sc_hs__nand2_1_87/a_117_74# sky130_fd_sc_hs__nand2_1
Xsky130_fd_sc_hs__inv_2_0 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_2_1/A sky130_fd_sc_hs__inv_2_1/Y
+ sky130_fd_sc_hs__inv_2
Xsky130_fd_sc_hs__a31oi_2_0 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__a32oi_1_9/Y sky130_fd_sc_hs__a31oi_2_1/A1
+ sky130_fd_sc_hs__o211ai_1_3/Y sky130_fd_sc_hs__a31oi_2_1/Y sky130_fd_sc_hs__nor2_1_61/B
+ sky130_fd_sc_hs__a31oi_2_1/a_114_74# sky130_fd_sc_hs__a31oi_2_1/a_27_368# sky130_fd_sc_hs__a31oi_2_1/a_200_74#
+ sky130_fd_sc_hs__a31oi_2
Xsky130_fd_sc_hs__o21ai_1_10 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__o21ai_1_11/Y sky130_fd_sc_hs__nand2_2_13/Y
+ sky130_fd_sc_hs__xnor2_1_3/A div_ratio_half[3] sky130_fd_sc_hs__o21ai_1_11/a_162_368#
+ sky130_fd_sc_hs__o21ai_1_11/a_27_74# sky130_fd_sc_hs__o21ai_1
Xsky130_fd_sc_hs__nand2_4_4 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_4_5/Y aux_osc_en
+ sky130_fd_sc_hs__nand2_4_9/Y sky130_fd_sc_hs__nand2_4_5/a_27_74# sky130_fd_sc_hs__nand2_4
Xsky130_fd_sc_hs__o211ai_1_10 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__a2bb2oi_1_1/Y sky130_fd_sc_hs__nor2_2_3/B
+ sky130_fd_sc_hs__nand2_2_11/Y sky130_fd_sc_hs__nand2_1_89/Y div_ratio_half[1] sky130_fd_sc_hs__o211ai_1_11/a_31_74#
+ sky130_fd_sc_hs__o211ai_1_11/a_311_74# sky130_fd_sc_hs__o211ai_1_11/a_116_368# sky130_fd_sc_hs__o211ai_1
Xsky130_fd_sc_hs__nor2_4_0 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__fa_2_9/B sky130_fd_sc_hs__or2_1_1/A
+ sky130_fd_sc_hs__nor2_4_1/B sky130_fd_sc_hs__nor2_4_1/a_27_368# sky130_fd_sc_hs__nor2_4
Xsky130_fd_sc_hs__a21oi_1_120 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__o21a_1_61/A2 sky130_fd_sc_hs__dfrbp_1_41/D
+ sky130_fd_sc_hs__o21a_1_75/B1 sky130_fd_sc_hs__inv_4_135/Y sky130_fd_sc_hs__a21oi_1_121/a_117_74#
+ sky130_fd_sc_hs__a21oi_1_121/a_29_368# sky130_fd_sc_hs__a21oi_1
Xsky130_fd_sc_hs__nand2_2_1 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_2_1/Y sky130_fd_sc_hs__nand2_2_1/B
+ sky130_fd_sc_hs__nand2_2_1/A sky130_fd_sc_hs__nand2_2_1/a_27_74# sky130_fd_sc_hs__nand2_2
Xsky130_fd_sc_hs__nor2_1_106 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__o21a_1_71/B1 sky130_fd_sc_hs__o21a_1_59/A2
+ sky130_fd_sc_hs__inv_4_129/Y sky130_fd_sc_hs__nor2_1_107/a_116_368# sky130_fd_sc_hs__nor2_1
Xsky130_fd_sc_hs__nor2_1_117 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_133/Y sky130_fd_sc_hs__nor3_1_9/C
+ sky130_fd_sc_hs__o21a_1_75/A1 sky130_fd_sc_hs__nor2_1_117/a_116_368# sky130_fd_sc_hs__nor2_1
Xsky130_fd_sc_hs__a22oi_1_15 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nor2_1_33/Y sky130_fd_sc_hs__a22oi_1_15/Y
+ sky130_fd_sc_hs__o21a_1_13/A1 sky130_fd_sc_hs__nor2b_1_25/Y sky130_fd_sc_hs__o21a_1_21/A1
+ sky130_fd_sc_hs__a22oi_1_15/a_71_368# sky130_fd_sc_hs__a22oi_1_15/a_159_74# sky130_fd_sc_hs__a22oi_1_15/a_339_74#
+ sky130_fd_sc_hs__a22oi_1
Xsky130_fd_sc_hs__nor2_1_83 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nor2_1_83/B sky130_fd_sc_hs__nor2_1_83/Y
+ sky130_fd_sc_hs__inv_4_89/Y sky130_fd_sc_hs__nor2_1_83/a_116_368# sky130_fd_sc_hs__nor2_1
Xsky130_fd_sc_hs__nor2_1_72 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nor2_1_73/B sky130_fd_sc_hs__nor2_1_73/Y
+ sky130_fd_sc_hs__inv_4_85/Y sky130_fd_sc_hs__nor2_1_73/a_116_368# sky130_fd_sc_hs__nor2_1
Xsky130_fd_sc_hs__nor2_1_61 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nor2_1_61/B sky130_fd_sc_hs__nor2_1_61/Y
+ sky130_fd_sc_hs__o22ai_1_3/Y sky130_fd_sc_hs__nor2_1_61/a_116_368# sky130_fd_sc_hs__nor2_1
Xsky130_fd_sc_hs__nor2_1_50 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nor2_1_51/B sky130_fd_sc_hs__nor2_1_51/Y
+ sky130_fd_sc_hs__inv_4_61/Y sky130_fd_sc_hs__nor2_1_51/a_116_368# sky130_fd_sc_hs__nor2_1
Xsky130_fd_sc_hs__nor2_1_94 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nor2_1_95/B sky130_fd_sc_hs__nor3_1_9/B
+ sky130_fd_sc_hs__nor2_1_95/A sky130_fd_sc_hs__nor2_1_95/a_116_368# sky130_fd_sc_hs__nor2_1
Xsky130_fd_sc_hs__xnor2_1_3 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__xnor2_1_3/A sky130_fd_sc_hs__xnor2_1_3/Y
+ sky130_fd_sc_hs__xnor2_1_3/B sky130_fd_sc_hs__xnor2_1_3/a_376_368# sky130_fd_sc_hs__xnor2_1_3/a_112_119#
+ sky130_fd_sc_hs__xnor2_1_3/a_138_385# sky130_fd_sc_hs__xnor2_1_3/a_293_74# sky130_fd_sc_hs__xnor2_1
Xsky130_fd_sc_hs__inv_4_120 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_121/Y sky130_fd_sc_hs__xnor2_1_3/B
+ sky130_fd_sc_hs__inv_4
Xsky130_fd_sc_hs__inv_4_131 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_2_7/B div_ratio_half[2]
+ sky130_fd_sc_hs__inv_4
Xsky130_fd_sc_hs__or2_1_2 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__or2_1_3/B sky130_fd_sc_hs__or2_1_3/A
+ sky130_fd_sc_hs__or2_1_3/X sky130_fd_sc_hs__or2_1_3/a_152_368# sky130_fd_sc_hs__or2_1_3/a_63_368#
+ sky130_fd_sc_hs__or2_1
Xsky130_fd_sc_hs__o21a_1_29 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__o21a_1_29/X sky130_fd_sc_hs__nor2_1_29/Y
+ sky130_fd_sc_hs__nor2_1_27/B sky130_fd_sc_hs__inv_4_39/A sky130_fd_sc_hs__o21a_1_29/a_320_74#
+ sky130_fd_sc_hs__o21a_1_29/a_376_387# sky130_fd_sc_hs__o21a_1_29/a_83_244# sky130_fd_sc_hs__o21a_1
Xsky130_fd_sc_hs__o21a_1_18 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__o21a_1_19/X sky130_fd_sc_hs__nor2_1_37/Y
+ sky130_fd_sc_hs__nor2_1_9/B sky130_fd_sc_hs__o21a_1_19/A1 sky130_fd_sc_hs__o21a_1_19/a_320_74#
+ sky130_fd_sc_hs__o21a_1_19/a_376_387# sky130_fd_sc_hs__o21a_1_19/a_83_244# sky130_fd_sc_hs__o21a_1
Xsky130_fd_sc_hs__dfrtp_4_19 DVSS DVDD sky130_fd_sc_hs__inv_4_49/Y DVDD DVSS sky130_fd_sc_hs__nor2b_1_3/Y
+ sky130_fd_sc_hs__dfstp_2_1/CLK sky130_fd_sc_hs__fa_2_3/B sky130_fd_sc_hs__dfrtp_4_19/a_37_78#
+ sky130_fd_sc_hs__dfrtp_4_19/a_494_366# sky130_fd_sc_hs__dfrtp_4_19/a_699_463# sky130_fd_sc_hs__dfrtp_4_19/a_313_74#
+ sky130_fd_sc_hs__dfrtp_4_19/a_1627_493# sky130_fd_sc_hs__dfrtp_4_19/a_1678_395#
+ sky130_fd_sc_hs__dfrtp_4_19/a_1827_81# sky130_fd_sc_hs__dfrtp_4_19/a_789_463# sky130_fd_sc_hs__dfrtp_4_19/a_1350_392#
+ sky130_fd_sc_hs__dfrtp_4_19/a_834_355# sky130_fd_sc_hs__dfrtp_4_19/a_812_138# sky130_fd_sc_hs__dfrtp_4_19/a_124_78#
+ sky130_fd_sc_hs__dfrtp_4_19/a_1647_81# sky130_fd_sc_hs__dfrtp_4_19/a_2010_409# sky130_fd_sc_hs__dfrtp_4_19/a_890_138#
+ sky130_fd_sc_hs__dfrtp_4
Xsky130_fd_sc_hs__inv_4_4 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_5/Y sky130_fd_sc_hs__inv_4_5/A
+ sky130_fd_sc_hs__inv_4
Xsky130_fd_sc_hs__a22o_1_21 DVSS DVDD DVDD DVSS osc_fine_con_final[8] manual_control_osc[8]
+ sky130_fd_sc_hs__inv_4_43/Y sky130_fd_sc_hs__fa_2_19/B fftl_en sky130_fd_sc_hs__a22o_1_21/a_222_392#
+ sky130_fd_sc_hs__a22o_1_21/a_230_79# sky130_fd_sc_hs__a22o_1_21/a_52_123# sky130_fd_sc_hs__a22o_1_21/a_132_392#
+ sky130_fd_sc_hs__a22o_1
Xsky130_fd_sc_hs__a22o_1_10 DVSS DVDD DVDD DVSS osc_fine_con_final[5] manual_control_osc[5]
+ sky130_fd_sc_hs__inv_4_43/Y sky130_fd_sc_hs__fa_2_11/B fftl_en sky130_fd_sc_hs__a22o_1_11/a_222_392#
+ sky130_fd_sc_hs__a22o_1_11/a_230_79# sky130_fd_sc_hs__a22o_1_11/a_52_123# sky130_fd_sc_hs__a22o_1_11/a_132_392#
+ sky130_fd_sc_hs__a22o_1
Xsky130_fd_sc_hs__nand4_1_4 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand4_1_5/C sky130_fd_sc_hs__nor3_1_3/C
+ sky130_fd_sc_hs__nand4_1_5/D sky130_fd_sc_hs__nor3_1_13/Y sky130_fd_sc_hs__nand4_1_5/A
+ sky130_fd_sc_hs__nand4_1_5/a_259_74# sky130_fd_sc_hs__nand4_1_5/a_373_74# sky130_fd_sc_hs__nand4_1_5/a_181_74#
+ sky130_fd_sc_hs__nand4_1
Xsky130_fd_sc_hs__nor4_1_0 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nor4_1_1/Y sky130_fd_sc_hs__nor4_1_1/D
+ sky130_fd_sc_hs__nor4_1_1/C sky130_fd_sc_hs__nor4_1_1/B sky130_fd_sc_hs__nor4_1_1/A
+ sky130_fd_sc_hs__nor4_1_1/a_144_368# sky130_fd_sc_hs__nor4_1_1/a_342_368# sky130_fd_sc_hs__nor4_1_1/a_228_368#
+ sky130_fd_sc_hs__nor4_1
Xsky130_fd_sc_hs__nand2_1_32 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nor2_1_25/Y sky130_fd_sc_hs__nor2_1_19/B
+ sky130_fd_sc_hs__o21a_1_25/A1 sky130_fd_sc_hs__nand2_1_33/a_117_74# sky130_fd_sc_hs__nand2_1
Xsky130_fd_sc_hs__nand2_1_21 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nor2_1_37/Y sky130_fd_sc_hs__nor2_1_9/B
+ sky130_fd_sc_hs__o21a_1_19/A1 sky130_fd_sc_hs__nand2_1_21/a_117_74# sky130_fd_sc_hs__nand2_1
Xsky130_fd_sc_hs__nand2_1_10 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__o21a_1_7/A2 sky130_fd_sc_hs__nor2_1_5/B
+ sky130_fd_sc_hs__o21a_1_7/A1 sky130_fd_sc_hs__nand2_1_11/a_117_74# sky130_fd_sc_hs__nand2_1
Xsky130_fd_sc_hs__nand2_1_76 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__o21a_1_59/A2 sky130_fd_sc_hs__nor2_1_87/B
+ sky130_fd_sc_hs__o21a_1_59/A1 sky130_fd_sc_hs__nand2_1_77/a_117_74# sky130_fd_sc_hs__nand2_1
Xsky130_fd_sc_hs__nand2_1_65 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nor2_1_51/Y sky130_fd_sc_hs__nor2_1_57/B
+ sky130_fd_sc_hs__nor2_1_59/A sky130_fd_sc_hs__nand2_1_65/a_117_74# sky130_fd_sc_hs__nand2_1
Xsky130_fd_sc_hs__nand2_1_54 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nor2_1_63/Y sky130_fd_sc_hs__nor2_1_43/B
+ sky130_fd_sc_hs__dfrbp_1_7/Q sky130_fd_sc_hs__nand2_1_55/a_117_74# sky130_fd_sc_hs__nand2_1
Xsky130_fd_sc_hs__nand2_1_43 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nor2_1_45/Y sky130_fd_sc_hs__nor2_1_29/B
+ sky130_fd_sc_hs__nor2_1_65/A sky130_fd_sc_hs__nand2_1_43/a_117_74# sky130_fd_sc_hs__nand2_1
Xsky130_fd_sc_hs__nand2_1_98 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__xnor2_1_11/Y sky130_fd_sc_hs__nor2_2_3/A
+ sky130_fd_sc_hs__nand2_1_99/A sky130_fd_sc_hs__nand2_1_99/a_117_74# sky130_fd_sc_hs__nand2_1
Xsky130_fd_sc_hs__nand2_1_87 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nor2_1_75/Y sky130_fd_sc_hs__nor2_1_99/B
+ sky130_fd_sc_hs__inv_4_97/A sky130_fd_sc_hs__nand2_1_87/a_117_74# sky130_fd_sc_hs__nand2_1
Xsky130_fd_sc_hs__dfxtp_4_0 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__dfxtp_4_2/Q sky130_fd_sc_hs__dfxtp_4_2/D
+ out_star sky130_fd_sc_hs__dfxtp_4_2/a_1226_296# sky130_fd_sc_hs__dfxtp_4_2/a_735_102#
+ sky130_fd_sc_hs__dfxtp_4_2/a_1141_508# sky130_fd_sc_hs__dfxtp_4_2/a_206_368# sky130_fd_sc_hs__dfxtp_4_2/a_437_503#
+ sky130_fd_sc_hs__dfxtp_4_2/a_27_74# sky130_fd_sc_hs__dfxtp_4_2/a_651_503# sky130_fd_sc_hs__dfxtp_4_2/a_696_458#
+ sky130_fd_sc_hs__dfxtp_4_2/a_544_485# sky130_fd_sc_hs__dfxtp_4_2/a_1178_124# sky130_fd_sc_hs__dfxtp_4_2/a_1034_424#
+ sky130_fd_sc_hs__dfxtp_4
Xsky130_fd_sc_hs__inv_2_1 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_2_1/A sky130_fd_sc_hs__inv_2_1/Y
+ sky130_fd_sc_hs__inv_2
Xsky130_fd_sc_hs__a31oi_2_1 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__a32oi_1_9/Y sky130_fd_sc_hs__a31oi_2_1/A1
+ sky130_fd_sc_hs__o211ai_1_3/Y sky130_fd_sc_hs__a31oi_2_1/Y sky130_fd_sc_hs__nor2_1_61/B
+ sky130_fd_sc_hs__a31oi_2_1/a_114_74# sky130_fd_sc_hs__a31oi_2_1/a_27_368# sky130_fd_sc_hs__a31oi_2_1/a_200_74#
+ sky130_fd_sc_hs__a31oi_2
Xsky130_fd_sc_hs__o21ai_1_11 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__o21ai_1_11/Y sky130_fd_sc_hs__nand2_2_13/Y
+ sky130_fd_sc_hs__xnor2_1_3/A div_ratio_half[3] sky130_fd_sc_hs__o21ai_1_11/a_162_368#
+ sky130_fd_sc_hs__o21ai_1_11/a_27_74# sky130_fd_sc_hs__o21ai_1
Xsky130_fd_sc_hs__nand2_4_5 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_4_5/Y aux_osc_en
+ sky130_fd_sc_hs__nand2_4_9/Y sky130_fd_sc_hs__nand2_4_5/a_27_74# sky130_fd_sc_hs__nand2_4
Xsky130_fd_sc_hs__o211ai_1_11 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__a2bb2oi_1_1/Y sky130_fd_sc_hs__nor2_2_3/B
+ sky130_fd_sc_hs__nand2_2_11/Y sky130_fd_sc_hs__nand2_1_89/Y div_ratio_half[1] sky130_fd_sc_hs__o211ai_1_11/a_31_74#
+ sky130_fd_sc_hs__o211ai_1_11/a_311_74# sky130_fd_sc_hs__o211ai_1_11/a_116_368# sky130_fd_sc_hs__o211ai_1
Xsky130_fd_sc_hs__nor2_4_1 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__fa_2_9/B sky130_fd_sc_hs__or2_1_1/A
+ sky130_fd_sc_hs__nor2_4_1/B sky130_fd_sc_hs__nor2_4_1/a_27_368# sky130_fd_sc_hs__nor2_4
Xsky130_fd_sc_hs__a21oi_1_110 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__o21a_1_71/A2 sky130_fd_sc_hs__dfrtn_1_31/D
+ sky130_fd_sc_hs__o21a_1_65/B1 sky130_fd_sc_hs__inv_4_99/Y sky130_fd_sc_hs__a21oi_1_111/a_117_74#
+ sky130_fd_sc_hs__a21oi_1_111/a_29_368# sky130_fd_sc_hs__a21oi_1
Xsky130_fd_sc_hs__a21oi_1_121 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__o21a_1_61/A2 sky130_fd_sc_hs__dfrbp_1_41/D
+ sky130_fd_sc_hs__o21a_1_75/B1 sky130_fd_sc_hs__inv_4_135/Y sky130_fd_sc_hs__a21oi_1_121/a_117_74#
+ sky130_fd_sc_hs__a21oi_1_121/a_29_368# sky130_fd_sc_hs__a21oi_1
Xsky130_fd_sc_hs__nor2b_2_0 DVSS DVDD DVDD DVSS rst sky130_fd_sc_hs__nor2b_1_43/Y
+ sky130_fd_sc_hs__nor2b_2_1/Y sky130_fd_sc_hs__nor2b_2_1/a_27_392# sky130_fd_sc_hs__nor2b_2_1/a_228_368#
+ sky130_fd_sc_hs__nor2b_2
Xsky130_fd_sc_hs__nand2_2_2 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_2_3/Y sky130_fd_sc_hs__nand2_2_3/B
+ sky130_fd_sc_hs__nand2_2_3/A sky130_fd_sc_hs__nand2_2_3/a_27_74# sky130_fd_sc_hs__nand2_2
Xsky130_fd_sc_hs__nor2_1_107 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__o21a_1_71/B1 sky130_fd_sc_hs__o21a_1_59/A2
+ sky130_fd_sc_hs__inv_4_129/Y sky130_fd_sc_hs__nor2_1_107/a_116_368# sky130_fd_sc_hs__nor2_1
Xsky130_fd_sc_hs__nor2_1_118 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__o21a_1_73/B1 sky130_fd_sc_hs__o21a_1_77/A2
+ sky130_fd_sc_hs__inv_4_115/Y sky130_fd_sc_hs__nor2_1_119/a_116_368# sky130_fd_sc_hs__nor2_1
Xsky130_fd_sc_hs__a22oi_1_16 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__a32oi_1_7/Y sky130_fd_sc_hs__o21ai_1_1/B1
+ sky130_fd_sc_hs__nor2_1_23/Y sky130_fd_sc_hs__a32oi_1_5/Y fine_control_avg_window_select[0]
+ sky130_fd_sc_hs__a22oi_1_17/a_71_368# sky130_fd_sc_hs__a22oi_1_17/a_159_74# sky130_fd_sc_hs__a22oi_1_17/a_339_74#
+ sky130_fd_sc_hs__a22oi_1
Xsky130_fd_sc_hs__nor2_1_40 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nor2_1_41/B sky130_fd_sc_hs__nor2_1_41/Y
+ sky130_fd_sc_hs__inv_4_51/Y sky130_fd_sc_hs__nor2_1_41/a_116_368# sky130_fd_sc_hs__nor2_1
Xsky130_fd_sc_hs__nor2_1_73 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nor2_1_73/B sky130_fd_sc_hs__nor2_1_73/Y
+ sky130_fd_sc_hs__inv_4_85/Y sky130_fd_sc_hs__nor2_1_73/a_116_368# sky130_fd_sc_hs__nor2_1
Xsky130_fd_sc_hs__nor2_1_62 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nor2_1_63/B sky130_fd_sc_hs__nor2_1_63/Y
+ sky130_fd_sc_hs__inv_4_71/Y sky130_fd_sc_hs__nor2_1_63/a_116_368# sky130_fd_sc_hs__nor2_1
Xsky130_fd_sc_hs__nor2_1_51 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nor2_1_51/B sky130_fd_sc_hs__nor2_1_51/Y
+ sky130_fd_sc_hs__inv_4_61/Y sky130_fd_sc_hs__nor2_1_51/a_116_368# sky130_fd_sc_hs__nor2_1
Xsky130_fd_sc_hs__nor2_1_95 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nor2_1_95/B sky130_fd_sc_hs__nor3_1_9/B
+ sky130_fd_sc_hs__nor2_1_95/A sky130_fd_sc_hs__nor2_1_95/a_116_368# sky130_fd_sc_hs__nor2_1
Xsky130_fd_sc_hs__nor2_1_84 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_59/Y sky130_fd_sc_hs__nor3_1_9/A
+ sky130_fd_sc_hs__inv_4_79/A sky130_fd_sc_hs__nor2_1_85/a_116_368# sky130_fd_sc_hs__nor2_1
Xsky130_fd_sc_hs__xnor2_1_4 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_95/A sky130_fd_sc_hs__xnor2_1_5/Y
+ sky130_fd_sc_hs__xnor2_1_5/B sky130_fd_sc_hs__xnor2_1_5/a_376_368# sky130_fd_sc_hs__xnor2_1_5/a_112_119#
+ sky130_fd_sc_hs__xnor2_1_5/a_138_385# sky130_fd_sc_hs__xnor2_1_5/a_293_74# sky130_fd_sc_hs__xnor2_1
Xsky130_fd_sc_hs__nor2b_1_40 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_87/Y sky130_fd_sc_hs__dfxtp_2_5/D
+ sky130_fd_sc_hs__nor2b_1_41/A sky130_fd_sc_hs__nor2b_1_41/a_278_368# sky130_fd_sc_hs__nor2b_1_41/a_27_112#
+ sky130_fd_sc_hs__nor2b_1
Xsky130_fd_sc_hs__inv_4_110 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nor2_1_99/A sky130_fd_sc_hs__inv_4_111/A
+ sky130_fd_sc_hs__inv_4
Xsky130_fd_sc_hs__inv_4_121 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_121/Y sky130_fd_sc_hs__xnor2_1_3/B
+ sky130_fd_sc_hs__inv_4
Xsky130_fd_sc_hs__inv_4_132 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_133/Y sky130_fd_sc_hs__inv_4_133/A
+ sky130_fd_sc_hs__inv_4
Xsky130_fd_sc_hs__nand2_4_10 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_4_9/A aux_osc_en
+ sky130_fd_sc_hs__nand2_4_13/Y sky130_fd_sc_hs__nand2_4_11/a_27_74# sky130_fd_sc_hs__nand2_4
Xsky130_fd_sc_hs__or2_1_3 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__or2_1_3/B sky130_fd_sc_hs__or2_1_3/A
+ sky130_fd_sc_hs__or2_1_3/X sky130_fd_sc_hs__or2_1_3/a_152_368# sky130_fd_sc_hs__or2_1_3/a_63_368#
+ sky130_fd_sc_hs__or2_1
Xsky130_fd_sc_hs__o21a_1_19 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__o21a_1_19/X sky130_fd_sc_hs__nor2_1_37/Y
+ sky130_fd_sc_hs__nor2_1_9/B sky130_fd_sc_hs__o21a_1_19/A1 sky130_fd_sc_hs__o21a_1_19/a_320_74#
+ sky130_fd_sc_hs__o21a_1_19/a_376_387# sky130_fd_sc_hs__o21a_1_19/a_83_244# sky130_fd_sc_hs__o21a_1
Xsky130_fd_sc_hs__inv_4_5 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_5/Y sky130_fd_sc_hs__inv_4_5/A
+ sky130_fd_sc_hs__inv_4
Xsky130_fd_sc_hs__clkbuf_2_0 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__clkbuf_2_1/X ref_clk
+ sky130_fd_sc_hs__clkbuf_2_1/a_43_192# sky130_fd_sc_hs__clkbuf_2
Xsky130_fd_sc_hs__a22o_1_22 DVSS DVDD DVDD DVSS osc_fine_con_final[9] manual_control_osc[9]
+ sky130_fd_sc_hs__inv_4_43/Y sky130_fd_sc_hs__fa_2_21/B fftl_en sky130_fd_sc_hs__a22o_1_23/a_222_392#
+ sky130_fd_sc_hs__a22o_1_23/a_230_79# sky130_fd_sc_hs__a22o_1_23/a_52_123# sky130_fd_sc_hs__a22o_1_23/a_132_392#
+ sky130_fd_sc_hs__a22o_1
Xsky130_fd_sc_hs__a22o_1_11 DVSS DVDD DVDD DVSS osc_fine_con_final[5] manual_control_osc[5]
+ sky130_fd_sc_hs__inv_4_43/Y sky130_fd_sc_hs__fa_2_11/B fftl_en sky130_fd_sc_hs__a22o_1_11/a_222_392#
+ sky130_fd_sc_hs__a22o_1_11/a_230_79# sky130_fd_sc_hs__a22o_1_11/a_52_123# sky130_fd_sc_hs__a22o_1_11/a_132_392#
+ sky130_fd_sc_hs__a22o_1
Xsky130_fd_sc_hs__nand4_1_5 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand4_1_5/C sky130_fd_sc_hs__nor3_1_3/C
+ sky130_fd_sc_hs__nand4_1_5/D sky130_fd_sc_hs__nor3_1_13/Y sky130_fd_sc_hs__nand4_1_5/A
+ sky130_fd_sc_hs__nand4_1_5/a_259_74# sky130_fd_sc_hs__nand4_1_5/a_373_74# sky130_fd_sc_hs__nand4_1_5/a_181_74#
+ sky130_fd_sc_hs__nand4_1
Xsky130_fd_sc_hs__sdlclkp_1_0 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__dfxtp_4_9/CLK clk_out
+ sky130_fd_sc_hs__nand2b_1_3/Y sky130_fd_sc_hs__conb_1_3/LO sky130_fd_sc_hs__sdlclkp_1_1/a_114_112#
+ sky130_fd_sc_hs__sdlclkp_1_1/a_667_80# sky130_fd_sc_hs__sdlclkp_1_1/a_1166_94# sky130_fd_sc_hs__sdlclkp_1_1/a_288_48#
+ sky130_fd_sc_hs__sdlclkp_1_1/a_722_492# sky130_fd_sc_hs__sdlclkp_1_1/a_1238_94#
+ sky130_fd_sc_hs__sdlclkp_1_1/a_116_424# sky130_fd_sc_hs__sdlclkp_1_1/a_709_54# sky130_fd_sc_hs__sdlclkp_1_1/a_566_74#
+ sky130_fd_sc_hs__sdlclkp_1_1/a_318_74# sky130_fd_sc_hs__sdlclkp_1
Xsky130_fd_sc_hs__nor4_1_1 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nor4_1_1/Y sky130_fd_sc_hs__nor4_1_1/D
+ sky130_fd_sc_hs__nor4_1_1/C sky130_fd_sc_hs__nor4_1_1/B sky130_fd_sc_hs__nor4_1_1/A
+ sky130_fd_sc_hs__nor4_1_1/a_144_368# sky130_fd_sc_hs__nor4_1_1/a_342_368# sky130_fd_sc_hs__nor4_1_1/a_228_368#
+ sky130_fd_sc_hs__nor4_1
Xsky130_fd_sc_hs__nand2_1_33 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nor2_1_25/Y sky130_fd_sc_hs__nor2_1_19/B
+ sky130_fd_sc_hs__o21a_1_25/A1 sky130_fd_sc_hs__nand2_1_33/a_117_74# sky130_fd_sc_hs__nand2_1
Xsky130_fd_sc_hs__nand2_1_22 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_23/A sky130_fd_sc_hs__nand2_1_23/Y
+ sky130_fd_sc_hs__or2_1_1/A sky130_fd_sc_hs__nand2_1_23/a_117_74# sky130_fd_sc_hs__nand2_1
Xsky130_fd_sc_hs__nand2_1_11 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__o21a_1_7/A2 sky130_fd_sc_hs__nor2_1_5/B
+ sky130_fd_sc_hs__o21a_1_7/A1 sky130_fd_sc_hs__nand2_1_11/a_117_74# sky130_fd_sc_hs__nand2_1
Xsky130_fd_sc_hs__nand2_1_66 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_65/Y sky130_fd_sc_hs__nand2_1_67/Y
+ sky130_fd_sc_hs__inv_4_89/A sky130_fd_sc_hs__nand2_1_67/a_117_74# sky130_fd_sc_hs__nand2_1
Xsky130_fd_sc_hs__nand2_1_55 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nor2_1_63/Y sky130_fd_sc_hs__nor2_1_43/B
+ sky130_fd_sc_hs__dfrbp_1_7/Q sky130_fd_sc_hs__nand2_1_55/a_117_74# sky130_fd_sc_hs__nand2_1
Xsky130_fd_sc_hs__nand2_1_44 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nor2_1_35/Y sky130_fd_sc_hs__nor2_1_37/B
+ sky130_fd_sc_hs__o21ai_1_3/B1 sky130_fd_sc_hs__nand2_1_45/a_117_74# sky130_fd_sc_hs__nand2_1
Xsky130_fd_sc_hs__nand2_1_99 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__xnor2_1_11/Y sky130_fd_sc_hs__nor2_2_3/A
+ sky130_fd_sc_hs__nand2_1_99/A sky130_fd_sc_hs__nand2_1_99/a_117_74# sky130_fd_sc_hs__nand2_1
Xsky130_fd_sc_hs__nand2_1_88 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_2_5/A sky130_fd_sc_hs__nand2_1_89/Y
+ sky130_fd_sc_hs__inv_2_3/Y sky130_fd_sc_hs__nand2_1_89/a_117_74# sky130_fd_sc_hs__nand2_1
Xsky130_fd_sc_hs__nand2_1_77 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__o21a_1_59/A2 sky130_fd_sc_hs__nor2_1_87/B
+ sky130_fd_sc_hs__o21a_1_59/A1 sky130_fd_sc_hs__nand2_1_77/a_117_74# sky130_fd_sc_hs__nand2_1
Xsky130_fd_sc_hs__inv_2_2 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_2_3/A sky130_fd_sc_hs__inv_2_3/Y
+ sky130_fd_sc_hs__inv_2
Xsky130_fd_sc_hs__dfxtp_4_1 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_91/A sky130_fd_sc_hs__inv_4_49/Y
+ ref_clk sky130_fd_sc_hs__dfxtp_4_3/a_1226_296# sky130_fd_sc_hs__dfxtp_4_3/a_735_102#
+ sky130_fd_sc_hs__dfxtp_4_3/a_1141_508# sky130_fd_sc_hs__dfxtp_4_3/a_206_368# sky130_fd_sc_hs__dfxtp_4_3/a_437_503#
+ sky130_fd_sc_hs__dfxtp_4_3/a_27_74# sky130_fd_sc_hs__dfxtp_4_3/a_651_503# sky130_fd_sc_hs__dfxtp_4_3/a_696_458#
+ sky130_fd_sc_hs__dfxtp_4_3/a_544_485# sky130_fd_sc_hs__dfxtp_4_3/a_1178_124# sky130_fd_sc_hs__dfxtp_4_3/a_1034_424#
+ sky130_fd_sc_hs__dfxtp_4
Xsky130_fd_sc_hs__nand2_4_6 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_4_7/Y aux_osc_en
+ sky130_fd_sc_hs__nand2_4_7/A sky130_fd_sc_hs__nand2_4_7/a_27_74# sky130_fd_sc_hs__nand2_4
Xsky130_fd_sc_hs__nor2_4_2 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_2_9/A div_ratio_half[0]
+ div_ratio_half[1] sky130_fd_sc_hs__nor2_4_3/a_27_368# sky130_fd_sc_hs__nor2_4
Xsky130_fd_sc_hs__a21oi_1_100 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nor2_1_99/Y sky130_fd_sc_hs__dfrtn_1_37/D
+ sky130_fd_sc_hs__nor2_1_99/B sky130_fd_sc_hs__nor2_1_99/A sky130_fd_sc_hs__a21oi_1_101/a_117_74#
+ sky130_fd_sc_hs__a21oi_1_101/a_29_368# sky130_fd_sc_hs__a21oi_1
Xsky130_fd_sc_hs__a21oi_1_111 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__o21a_1_71/A2 sky130_fd_sc_hs__dfrtn_1_31/D
+ sky130_fd_sc_hs__o21a_1_65/B1 sky130_fd_sc_hs__inv_4_99/Y sky130_fd_sc_hs__a21oi_1_111/a_117_74#
+ sky130_fd_sc_hs__a21oi_1_111/a_29_368# sky130_fd_sc_hs__a21oi_1
Xsky130_fd_sc_hs__a21oi_1_122 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__o21a_1_63/A2 sky130_fd_sc_hs__dfrbp_1_43/D
+ sky130_fd_sc_hs__o21a_1_77/B1 sky130_fd_sc_hs__inv_4_137/Y sky130_fd_sc_hs__a21oi_1_123/a_117_74#
+ sky130_fd_sc_hs__a21oi_1_123/a_29_368# sky130_fd_sc_hs__a21oi_1
Xsky130_fd_sc_hs__nor2b_2_1 DVSS DVDD DVDD DVSS rst sky130_fd_sc_hs__nor2b_1_43/Y
+ sky130_fd_sc_hs__nor2b_2_1/Y sky130_fd_sc_hs__nor2b_2_1/a_27_392# sky130_fd_sc_hs__nor2b_2_1/a_228_368#
+ sky130_fd_sc_hs__nor2b_2
Xsky130_fd_sc_hs__nand2_2_3 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_2_3/Y sky130_fd_sc_hs__nand2_2_3/B
+ sky130_fd_sc_hs__nand2_2_3/A sky130_fd_sc_hs__nand2_2_3/a_27_74# sky130_fd_sc_hs__nand2_2
Xsky130_fd_sc_hs__nor2_1_108 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_113/Y sky130_fd_sc_hs__nor3_1_15/B
+ sky130_fd_sc_hs__o21a_1_71/A1 sky130_fd_sc_hs__nor2_1_109/a_116_368# sky130_fd_sc_hs__nor2_1
Xsky130_fd_sc_hs__nor2_1_119 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__o21a_1_73/B1 sky130_fd_sc_hs__o21a_1_77/A2
+ sky130_fd_sc_hs__inv_4_115/Y sky130_fd_sc_hs__nor2_1_119/a_116_368# sky130_fd_sc_hs__nor2_1
Xsky130_fd_sc_hs__a22oi_1_17 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__a32oi_1_7/Y sky130_fd_sc_hs__o21ai_1_1/B1
+ sky130_fd_sc_hs__nor2_1_23/Y sky130_fd_sc_hs__a32oi_1_5/Y fine_control_avg_window_select[0]
+ sky130_fd_sc_hs__a22oi_1_17/a_71_368# sky130_fd_sc_hs__a22oi_1_17/a_159_74# sky130_fd_sc_hs__a22oi_1_17/a_339_74#
+ sky130_fd_sc_hs__a22oi_1
Xsky130_fd_sc_hs__nor2_1_30 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nor2_1_31/B sky130_fd_sc_hs__nor2_1_31/Y
+ sky130_fd_sc_hs__inv_4_45/Y sky130_fd_sc_hs__nor2_1_31/a_116_368# sky130_fd_sc_hs__nor2_1
Xsky130_fd_sc_hs__nor2_1_74 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nor2_1_75/B sky130_fd_sc_hs__nor2_1_75/Y
+ sky130_fd_sc_hs__inv_4_75/Y sky130_fd_sc_hs__nor2_1_75/a_116_368# sky130_fd_sc_hs__nor2_1
Xsky130_fd_sc_hs__nor2_1_63 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nor2_1_63/B sky130_fd_sc_hs__nor2_1_63/Y
+ sky130_fd_sc_hs__inv_4_71/Y sky130_fd_sc_hs__nor2_1_63/a_116_368# sky130_fd_sc_hs__nor2_1
Xsky130_fd_sc_hs__nor2_1_52 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_91/A sky130_fd_sc_hs__nor2_1_53/Y
+ rst sky130_fd_sc_hs__nor2_1_53/a_116_368# sky130_fd_sc_hs__nor2_1
Xsky130_fd_sc_hs__nor2_1_41 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nor2_1_41/B sky130_fd_sc_hs__nor2_1_41/Y
+ sky130_fd_sc_hs__inv_4_51/Y sky130_fd_sc_hs__nor2_1_41/a_116_368# sky130_fd_sc_hs__nor2_1
Xsky130_fd_sc_hs__nor2_1_96 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nor2_1_99/A sky130_fd_sc_hs__nor3_1_5/C
+ sky130_fd_sc_hs__nor2_1_97/A sky130_fd_sc_hs__nor2_1_97/a_116_368# sky130_fd_sc_hs__nor2_1
Xsky130_fd_sc_hs__nor2_1_85 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_59/Y sky130_fd_sc_hs__nor3_1_9/A
+ sky130_fd_sc_hs__inv_4_79/A sky130_fd_sc_hs__nor2_1_85/a_116_368# sky130_fd_sc_hs__nor2_1
Xsky130_fd_sc_hs__xnor2_1_5 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_95/A sky130_fd_sc_hs__xnor2_1_5/Y
+ sky130_fd_sc_hs__xnor2_1_5/B sky130_fd_sc_hs__xnor2_1_5/a_376_368# sky130_fd_sc_hs__xnor2_1_5/a_112_119#
+ sky130_fd_sc_hs__xnor2_1_5/a_138_385# sky130_fd_sc_hs__xnor2_1_5/a_293_74# sky130_fd_sc_hs__xnor2_1
Xsky130_fd_sc_hs__nor2b_1_41 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_87/Y sky130_fd_sc_hs__dfxtp_2_5/D
+ sky130_fd_sc_hs__nor2b_1_41/A sky130_fd_sc_hs__nor2b_1_41/a_278_368# sky130_fd_sc_hs__nor2b_1_41/a_27_112#
+ sky130_fd_sc_hs__nor2b_1
Xsky130_fd_sc_hs__nor2b_1_30 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_87/A sky130_fd_sc_hs__dfxtp_4_5/D
+ rst sky130_fd_sc_hs__nor2b_1_31/a_278_368# sky130_fd_sc_hs__nor2b_1_31/a_27_112#
+ sky130_fd_sc_hs__nor2b_1
Xsky130_fd_sc_hs__inv_4_100 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__or2_1_3/B sky130_fd_sc_hs__inv_4_101/A
+ sky130_fd_sc_hs__inv_4
Xsky130_fd_sc_hs__inv_4_111 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nor2_1_99/A sky130_fd_sc_hs__inv_4_111/A
+ sky130_fd_sc_hs__inv_4
Xsky130_fd_sc_hs__inv_4_122 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_123/Y div_ratio_half[1]
+ sky130_fd_sc_hs__inv_4
Xsky130_fd_sc_hs__inv_4_133 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_133/Y sky130_fd_sc_hs__inv_4_133/A
+ sky130_fd_sc_hs__inv_4
Xsky130_fd_sc_hs__o22ai_1_0 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_33/Y sky130_fd_sc_hs__a32oi_1_3/Y
+ sky130_fd_sc_hs__o22ai_1_1/Y sky130_fd_sc_hs__o22ai_1_1/A2 sky130_fd_sc_hs__o22ai_1_1/A1
+ sky130_fd_sc_hs__o22ai_1_1/a_340_368# sky130_fd_sc_hs__o22ai_1_1/a_142_368# sky130_fd_sc_hs__o22ai_1_1/a_27_74#
+ sky130_fd_sc_hs__o22ai_1
Xsky130_fd_sc_hs__nand2_4_11 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_4_9/A aux_osc_en
+ sky130_fd_sc_hs__nand2_4_13/Y sky130_fd_sc_hs__nand2_4_11/a_27_74# sky130_fd_sc_hs__nand2_4
Xsky130_fd_sc_hs__inv_4_6 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_7/Y sky130_fd_sc_hs__inv_4_7/A
+ sky130_fd_sc_hs__inv_4
Xsky130_fd_sc_hs__clkbuf_2_1 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__clkbuf_2_1/X ref_clk
+ sky130_fd_sc_hs__clkbuf_2_1/a_43_192# sky130_fd_sc_hs__clkbuf_2
Xsky130_fd_sc_hs__a22o_1_23 DVSS DVDD DVDD DVSS osc_fine_con_final[9] manual_control_osc[9]
+ sky130_fd_sc_hs__inv_4_43/Y sky130_fd_sc_hs__fa_2_21/B fftl_en sky130_fd_sc_hs__a22o_1_23/a_222_392#
+ sky130_fd_sc_hs__a22o_1_23/a_230_79# sky130_fd_sc_hs__a22o_1_23/a_52_123# sky130_fd_sc_hs__a22o_1_23/a_132_392#
+ sky130_fd_sc_hs__a22o_1
Xsky130_fd_sc_hs__a22o_1_12 DVSS DVDD DVDD DVSS osc_fine_con_final[11] manual_control_osc[11]
+ sky130_fd_sc_hs__inv_4_43/Y sky130_fd_sc_hs__fa_2_15/B fftl_en sky130_fd_sc_hs__a22o_1_13/a_222_392#
+ sky130_fd_sc_hs__a22o_1_13/a_230_79# sky130_fd_sc_hs__a22o_1_13/a_52_123# sky130_fd_sc_hs__a22o_1_13/a_132_392#
+ sky130_fd_sc_hs__a22o_1
Xsky130_fd_sc_hs__sdlclkp_1_1 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__dfxtp_4_9/CLK clk_out
+ sky130_fd_sc_hs__nand2b_1_3/Y sky130_fd_sc_hs__conb_1_3/LO sky130_fd_sc_hs__sdlclkp_1_1/a_114_112#
+ sky130_fd_sc_hs__sdlclkp_1_1/a_667_80# sky130_fd_sc_hs__sdlclkp_1_1/a_1166_94# sky130_fd_sc_hs__sdlclkp_1_1/a_288_48#
+ sky130_fd_sc_hs__sdlclkp_1_1/a_722_492# sky130_fd_sc_hs__sdlclkp_1_1/a_1238_94#
+ sky130_fd_sc_hs__sdlclkp_1_1/a_116_424# sky130_fd_sc_hs__sdlclkp_1_1/a_709_54# sky130_fd_sc_hs__sdlclkp_1_1/a_566_74#
+ sky130_fd_sc_hs__sdlclkp_1_1/a_318_74# sky130_fd_sc_hs__sdlclkp_1
Xsky130_fd_sc_hs__nor4_1_2 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nor4_1_3/Y sky130_fd_sc_hs__nor4_1_3/D
+ sky130_fd_sc_hs__nor4_1_3/C sky130_fd_sc_hs__nor4_1_3/B sky130_fd_sc_hs__nor4_1_3/A
+ sky130_fd_sc_hs__nor4_1_3/a_144_368# sky130_fd_sc_hs__nor4_1_3/a_342_368# sky130_fd_sc_hs__nor4_1_3/a_228_368#
+ sky130_fd_sc_hs__nor4_1
Xsky130_fd_sc_hs__nand2_1_23 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_23/A sky130_fd_sc_hs__nand2_1_23/Y
+ sky130_fd_sc_hs__or2_1_1/A sky130_fd_sc_hs__nand2_1_23/a_117_74# sky130_fd_sc_hs__nand2_1
Xsky130_fd_sc_hs__nand2_1_12 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nor2_1_11/Y sky130_fd_sc_hs__nor2_1_31/B
+ sky130_fd_sc_hs__o21a_1_13/A1 sky130_fd_sc_hs__nand2_1_13/a_117_74# sky130_fd_sc_hs__nand2_1
Xsky130_fd_sc_hs__nand2_1_67 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_65/Y sky130_fd_sc_hs__nand2_1_67/Y
+ sky130_fd_sc_hs__inv_4_89/A sky130_fd_sc_hs__nand2_1_67/a_117_74# sky130_fd_sc_hs__nand2_1
Xsky130_fd_sc_hs__nand2_1_56 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_69/Y sky130_fd_sc_hs__nand4_1_1/D
+ sky130_fd_sc_hs__nor2_1_69/B sky130_fd_sc_hs__nand2_1_57/a_117_74# sky130_fd_sc_hs__nand2_1
Xsky130_fd_sc_hs__nand2_1_45 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nor2_1_35/Y sky130_fd_sc_hs__nor2_1_37/B
+ sky130_fd_sc_hs__o21ai_1_3/B1 sky130_fd_sc_hs__nand2_1_45/a_117_74# sky130_fd_sc_hs__nand2_1
Xsky130_fd_sc_hs__nand2_1_34 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nor2_1_31/Y sky130_fd_sc_hs__nor2_1_21/B
+ sky130_fd_sc_hs__o21a_1_27/A1 sky130_fd_sc_hs__nand2_1_35/a_117_74# sky130_fd_sc_hs__nand2_1
Xsky130_fd_sc_hs__nand2_1_89 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_2_5/A sky130_fd_sc_hs__nand2_1_89/Y
+ sky130_fd_sc_hs__inv_2_3/Y sky130_fd_sc_hs__nand2_1_89/a_117_74# sky130_fd_sc_hs__nand2_1
Xsky130_fd_sc_hs__nand2_1_78 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_1_91/A sky130_fd_sc_hs__or3b_2_1/C_N
+ sky130_fd_sc_hs__nand2_1_89/Y sky130_fd_sc_hs__nand2_1_79/a_117_74# sky130_fd_sc_hs__nand2_1
Xsky130_fd_sc_hs__inv_2_3 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_2_3/A sky130_fd_sc_hs__inv_2_3/Y
+ sky130_fd_sc_hs__inv_2
Xsky130_fd_sc_hs__dfxtp_4_2 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__dfxtp_4_2/Q sky130_fd_sc_hs__dfxtp_4_2/D
+ out_star sky130_fd_sc_hs__dfxtp_4_2/a_1226_296# sky130_fd_sc_hs__dfxtp_4_2/a_735_102#
+ sky130_fd_sc_hs__dfxtp_4_2/a_1141_508# sky130_fd_sc_hs__dfxtp_4_2/a_206_368# sky130_fd_sc_hs__dfxtp_4_2/a_437_503#
+ sky130_fd_sc_hs__dfxtp_4_2/a_27_74# sky130_fd_sc_hs__dfxtp_4_2/a_651_503# sky130_fd_sc_hs__dfxtp_4_2/a_696_458#
+ sky130_fd_sc_hs__dfxtp_4_2/a_544_485# sky130_fd_sc_hs__dfxtp_4_2/a_1178_124# sky130_fd_sc_hs__dfxtp_4_2/a_1034_424#
+ sky130_fd_sc_hs__dfxtp_4
Xsky130_fd_sc_hs__nand2_4_7 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_4_7/Y aux_osc_en
+ sky130_fd_sc_hs__nand2_4_7/A sky130_fd_sc_hs__nand2_4_7/a_27_74# sky130_fd_sc_hs__nand2_4
Xsky130_fd_sc_hs__nor2_4_3 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_2_9/A div_ratio_half[0]
+ div_ratio_half[1] sky130_fd_sc_hs__nor2_4_3/a_27_368# sky130_fd_sc_hs__nor2_4
Xsky130_fd_sc_hs__a21oi_1_101 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nor2_1_99/Y sky130_fd_sc_hs__dfrtn_1_37/D
+ sky130_fd_sc_hs__nor2_1_99/B sky130_fd_sc_hs__nor2_1_99/A sky130_fd_sc_hs__a21oi_1_101/a_117_74#
+ sky130_fd_sc_hs__a21oi_1_101/a_29_368# sky130_fd_sc_hs__a21oi_1
Xsky130_fd_sc_hs__a21oi_1_112 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__o21a_1_73/A2 sky130_fd_sc_hs__dfrbp_1_29/D
+ sky130_fd_sc_hs__o21a_1_53/B1 sky130_fd_sc_hs__inv_4_117/Y sky130_fd_sc_hs__a21oi_1_113/a_117_74#
+ sky130_fd_sc_hs__a21oi_1_113/a_29_368# sky130_fd_sc_hs__a21oi_1
Xsky130_fd_sc_hs__a21oi_1_123 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__o21a_1_63/A2 sky130_fd_sc_hs__dfrbp_1_43/D
+ sky130_fd_sc_hs__o21a_1_77/B1 sky130_fd_sc_hs__inv_4_137/Y sky130_fd_sc_hs__a21oi_1_123/a_117_74#
+ sky130_fd_sc_hs__a21oi_1_123/a_29_368# sky130_fd_sc_hs__a21oi_1
Xsky130_fd_sc_hs__nand2_2_4 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__xnor2_1_3/B sky130_fd_sc_hs__nand2_2_5/B
+ sky130_fd_sc_hs__and2_2_5/X sky130_fd_sc_hs__nand2_2_5/a_27_74# sky130_fd_sc_hs__nand2_2
Xsky130_fd_sc_hs__nor2_2_0 DVSS DVDD DVDD DVSS rst sky130_fd_sc_hs__nor2_2_1/Y sky130_fd_sc_hs__nor2_2_1/A
+ sky130_fd_sc_hs__nor2_2_1/a_35_368# sky130_fd_sc_hs__nor2_2
Xsky130_fd_sc_hs__nor2_1_109 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_113/Y sky130_fd_sc_hs__nor3_1_15/B
+ sky130_fd_sc_hs__o21a_1_71/A1 sky130_fd_sc_hs__nor2_1_109/a_116_368# sky130_fd_sc_hs__nor2_1
Xsky130_fd_sc_hs__a22oi_1_18 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nor2b_1_25/Y sky130_fd_sc_hs__a32oi_1_7/A1
+ sky130_fd_sc_hs__o21a_1_27/A1 sky130_fd_sc_hs__nor2b_1_23/Y sky130_fd_sc_hs__o21a_1_25/A1
+ sky130_fd_sc_hs__a22oi_1_19/a_71_368# sky130_fd_sc_hs__a22oi_1_19/a_159_74# sky130_fd_sc_hs__a22oi_1_19/a_339_74#
+ sky130_fd_sc_hs__a22oi_1
Xsky130_fd_sc_hs__nor2_1_31 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nor2_1_31/B sky130_fd_sc_hs__nor2_1_31/Y
+ sky130_fd_sc_hs__inv_4_45/Y sky130_fd_sc_hs__nor2_1_31/a_116_368# sky130_fd_sc_hs__nor2_1
Xsky130_fd_sc_hs__nor2_1_20 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nor2_1_21/B sky130_fd_sc_hs__nor2_1_21/Y
+ sky130_fd_sc_hs__inv_4_31/Y sky130_fd_sc_hs__nor2_1_21/a_116_368# sky130_fd_sc_hs__nor2_1
Xsky130_fd_sc_hs__nor2_1_64 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_73/Y sky130_fd_sc_hs__nor2_1_65/Y
+ sky130_fd_sc_hs__nor2_1_65/A sky130_fd_sc_hs__nor2_1_65/a_116_368# sky130_fd_sc_hs__nor2_1
Xsky130_fd_sc_hs__nor2_1_53 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_91/A sky130_fd_sc_hs__nor2_1_53/Y
+ rst sky130_fd_sc_hs__nor2_1_53/a_116_368# sky130_fd_sc_hs__nor2_1
Xsky130_fd_sc_hs__nor2_1_42 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nor2_1_43/B sky130_fd_sc_hs__nor2_1_43/Y
+ sky130_fd_sc_hs__inv_4_67/Y sky130_fd_sc_hs__nor2_1_43/a_116_368# sky130_fd_sc_hs__nor2_1
Xsky130_fd_sc_hs__nor2_1_97 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nor2_1_99/A sky130_fd_sc_hs__nor3_1_5/C
+ sky130_fd_sc_hs__nor2_1_97/A sky130_fd_sc_hs__nor2_1_97/a_116_368# sky130_fd_sc_hs__nor2_1
Xsky130_fd_sc_hs__nor2_1_86 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nor2_1_87/B sky130_fd_sc_hs__nor2_1_87/Y
+ sky130_fd_sc_hs__inv_4_81/Y sky130_fd_sc_hs__nor2_1_87/a_116_368# sky130_fd_sc_hs__nor2_1
Xsky130_fd_sc_hs__nor2_1_75 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nor2_1_75/B sky130_fd_sc_hs__nor2_1_75/Y
+ sky130_fd_sc_hs__inv_4_75/Y sky130_fd_sc_hs__nor2_1_75/a_116_368# sky130_fd_sc_hs__nor2_1
Xsky130_fd_sc_hs__xnor2_1_6 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__xnor2_1_7/A sky130_fd_sc_hs__xnor2_1_7/Y
+ sky130_fd_sc_hs__xnor2_1_7/B sky130_fd_sc_hs__xnor2_1_7/a_376_368# sky130_fd_sc_hs__xnor2_1_7/a_112_119#
+ sky130_fd_sc_hs__xnor2_1_7/a_138_385# sky130_fd_sc_hs__xnor2_1_7/a_293_74# sky130_fd_sc_hs__xnor2_1
Xsky130_fd_sc_hs__nor2b_1_31 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_87/A sky130_fd_sc_hs__dfxtp_4_5/D
+ rst sky130_fd_sc_hs__nor2b_1_31/a_278_368# sky130_fd_sc_hs__nor2b_1_31/a_27_112#
+ sky130_fd_sc_hs__nor2b_1
Xsky130_fd_sc_hs__nor2b_1_20 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__fa_2_23/SUM sky130_fd_sc_hs__nor2b_1_21/Y
+ sky130_fd_sc_hs__or2_1_1/A sky130_fd_sc_hs__nor2b_1_21/a_278_368# sky130_fd_sc_hs__nor2b_1_21/a_27_112#
+ sky130_fd_sc_hs__nor2b_1
Xsky130_fd_sc_hs__nor2b_1_42 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nor2_1_101/Y sky130_fd_sc_hs__nor2b_1_43/Y
+ sky130_fd_sc_hs__inv_4_87/A sky130_fd_sc_hs__nor2b_1_43/a_278_368# sky130_fd_sc_hs__nor2b_1_43/a_27_112#
+ sky130_fd_sc_hs__nor2b_1
Xsky130_fd_sc_hs__inv_4_101 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__or2_1_3/B sky130_fd_sc_hs__inv_4_101/A
+ sky130_fd_sc_hs__inv_4
Xsky130_fd_sc_hs__inv_4_112 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_113/Y sky130_fd_sc_hs__inv_4_113/A
+ sky130_fd_sc_hs__inv_4
Xsky130_fd_sc_hs__inv_4_123 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_123/Y div_ratio_half[1]
+ sky130_fd_sc_hs__inv_4
Xsky130_fd_sc_hs__inv_4_134 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_135/Y sky130_fd_sc_hs__inv_4_135/A
+ sky130_fd_sc_hs__inv_4
Xsky130_fd_sc_hs__o22ai_1_1 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_33/Y sky130_fd_sc_hs__a32oi_1_3/Y
+ sky130_fd_sc_hs__o22ai_1_1/Y sky130_fd_sc_hs__o22ai_1_1/A2 sky130_fd_sc_hs__o22ai_1_1/A1
+ sky130_fd_sc_hs__o22ai_1_1/a_340_368# sky130_fd_sc_hs__o22ai_1_1/a_142_368# sky130_fd_sc_hs__o22ai_1_1/a_27_74#
+ sky130_fd_sc_hs__o22ai_1
Xsky130_fd_sc_hs__nand2_4_12 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_4_13/Y aux_osc_en
+ sky130_fd_sc_hs__nand2_4_7/Y sky130_fd_sc_hs__nand2_4_13/a_27_74# sky130_fd_sc_hs__nand2_4
Xsky130_fd_sc_hs__inv_4_7 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_7/Y sky130_fd_sc_hs__inv_4_7/A
+ sky130_fd_sc_hs__inv_4
Xsky130_fd_sc_hs__a22o_1_13 DVSS DVDD DVDD DVSS osc_fine_con_final[11] manual_control_osc[11]
+ sky130_fd_sc_hs__inv_4_43/Y sky130_fd_sc_hs__fa_2_15/B fftl_en sky130_fd_sc_hs__a22o_1_13/a_222_392#
+ sky130_fd_sc_hs__a22o_1_13/a_230_79# sky130_fd_sc_hs__a22o_1_13/a_52_123# sky130_fd_sc_hs__a22o_1_13/a_132_392#
+ sky130_fd_sc_hs__a22o_1
Xsky130_fd_sc_hs__a22o_1_24 DVSS DVDD DVDD DVSS osc_fine_con_final[10] manual_control_osc[10]
+ sky130_fd_sc_hs__inv_4_43/Y sky130_fd_sc_hs__fa_2_23/B fftl_en sky130_fd_sc_hs__a22o_1_25/a_222_392#
+ sky130_fd_sc_hs__a22o_1_25/a_230_79# sky130_fd_sc_hs__a22o_1_25/a_52_123# sky130_fd_sc_hs__a22o_1_25/a_132_392#
+ sky130_fd_sc_hs__a22o_1
Xsky130_fd_sc_hs__o21ai_1_0 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__o21ai_1_1/Y sky130_fd_sc_hs__o21ai_1_1/B1
+ sky130_fd_sc_hs__a32oi_1_1/Y fine_control_avg_window_select[0] sky130_fd_sc_hs__o21ai_1_1/a_162_368#
+ sky130_fd_sc_hs__o21ai_1_1/a_27_74# sky130_fd_sc_hs__o21ai_1
Xsky130_fd_sc_hs__nor4_1_3 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nor4_1_3/Y sky130_fd_sc_hs__nor4_1_3/D
+ sky130_fd_sc_hs__nor4_1_3/C sky130_fd_sc_hs__nor4_1_3/B sky130_fd_sc_hs__nor4_1_3/A
+ sky130_fd_sc_hs__nor4_1_3/a_144_368# sky130_fd_sc_hs__nor4_1_3/a_342_368# sky130_fd_sc_hs__nor4_1_3/a_228_368#
+ sky130_fd_sc_hs__nor4_1
Xsky130_fd_sc_hs__nand2_1_24 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nor2_1_13/Y sky130_fd_sc_hs__nor2_1_25/B
+ sky130_fd_sc_hs__o21a_1_21/A1 sky130_fd_sc_hs__nand2_1_25/a_117_74# sky130_fd_sc_hs__nand2_1
Xsky130_fd_sc_hs__nand2_1_13 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nor2_1_11/Y sky130_fd_sc_hs__nor2_1_31/B
+ sky130_fd_sc_hs__o21a_1_13/A1 sky130_fd_sc_hs__nand2_1_13/a_117_74# sky130_fd_sc_hs__nand2_1
Xsky130_fd_sc_hs__nand2_1_57 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_69/Y sky130_fd_sc_hs__nand4_1_1/D
+ sky130_fd_sc_hs__nor2_1_69/B sky130_fd_sc_hs__nand2_1_57/a_117_74# sky130_fd_sc_hs__nand2_1
Xsky130_fd_sc_hs__nand2_1_46 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_1_47/B sky130_fd_sc_hs__nor2_1_75/B
+ sky130_fd_sc_hs__nor2b_1_33/Y sky130_fd_sc_hs__nand2_1_47/a_117_74# sky130_fd_sc_hs__nand2_1
Xsky130_fd_sc_hs__nand2_1_35 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nor2_1_31/Y sky130_fd_sc_hs__nor2_1_21/B
+ sky130_fd_sc_hs__o21a_1_27/A1 sky130_fd_sc_hs__nand2_1_35/a_117_74# sky130_fd_sc_hs__nand2_1
Xsky130_fd_sc_hs__nand2_1_79 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_1_91/A sky130_fd_sc_hs__or3b_2_1/C_N
+ sky130_fd_sc_hs__nand2_1_89/Y sky130_fd_sc_hs__nand2_1_79/a_117_74# sky130_fd_sc_hs__nand2_1
Xsky130_fd_sc_hs__nand2_1_68 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nor2_1_47/Y sky130_fd_sc_hs__o21a_1_57/B1
+ sky130_fd_sc_hs__inv_4_93/A sky130_fd_sc_hs__nand2_1_69/a_117_74# sky130_fd_sc_hs__nand2_1
Xsky130_fd_sc_hs__inv_2_4 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_2_5/A sky130_fd_sc_hs__inv_2_5/Y
+ sky130_fd_sc_hs__inv_2
Xsky130_fd_sc_hs__dfxtp_4_3 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_91/A sky130_fd_sc_hs__inv_4_49/Y
+ ref_clk sky130_fd_sc_hs__dfxtp_4_3/a_1226_296# sky130_fd_sc_hs__dfxtp_4_3/a_735_102#
+ sky130_fd_sc_hs__dfxtp_4_3/a_1141_508# sky130_fd_sc_hs__dfxtp_4_3/a_206_368# sky130_fd_sc_hs__dfxtp_4_3/a_437_503#
+ sky130_fd_sc_hs__dfxtp_4_3/a_27_74# sky130_fd_sc_hs__dfxtp_4_3/a_651_503# sky130_fd_sc_hs__dfxtp_4_3/a_696_458#
+ sky130_fd_sc_hs__dfxtp_4_3/a_544_485# sky130_fd_sc_hs__dfxtp_4_3/a_1178_124# sky130_fd_sc_hs__dfxtp_4_3/a_1034_424#
+ sky130_fd_sc_hs__dfxtp_4
Xsky130_fd_sc_hs__nand2_4_8 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_4_9/Y aux_osc_en
+ sky130_fd_sc_hs__nand2_4_9/A sky130_fd_sc_hs__nand2_4_9/a_27_74# sky130_fd_sc_hs__nand2_4
Xsky130_fd_sc_hs__dfxtp_2_0 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__xnor2_1_3/A sky130_fd_sc_hs__dfxtp_4_9/CLK
+ sky130_fd_sc_hs__inv_2_1/Y sky130_fd_sc_hs__dfxtp_2_1/a_431_508# sky130_fd_sc_hs__dfxtp_2_1/a_1125_508#
+ sky130_fd_sc_hs__dfxtp_2_1/a_206_368# sky130_fd_sc_hs__dfxtp_2_1/a_27_74# sky130_fd_sc_hs__dfxtp_2_1/a_708_101#
+ sky130_fd_sc_hs__dfxtp_2_1/a_1019_424# sky130_fd_sc_hs__dfxtp_2_1/a_1172_124# sky130_fd_sc_hs__dfxtp_2_1/a_644_504#
+ sky130_fd_sc_hs__dfxtp_2_1/a_1217_314# sky130_fd_sc_hs__dfxtp_2_1/a_538_429# sky130_fd_sc_hs__dfxtp_2_1/a_695_459#
+ sky130_fd_sc_hs__dfxtp_2
Xsky130_fd_sc_hs__a21oi_1_102 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_123/Y sky130_fd_sc_hs__nand2_1_91/B
+ div_ratio_half[0] sky130_fd_sc_hs__inv_2_5/A sky130_fd_sc_hs__a21oi_1_103/a_117_74#
+ sky130_fd_sc_hs__a21oi_1_103/a_29_368# sky130_fd_sc_hs__a21oi_1
Xsky130_fd_sc_hs__a21oi_1_113 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__o21a_1_73/A2 sky130_fd_sc_hs__dfrbp_1_29/D
+ sky130_fd_sc_hs__o21a_1_53/B1 sky130_fd_sc_hs__inv_4_117/Y sky130_fd_sc_hs__a21oi_1_113/a_117_74#
+ sky130_fd_sc_hs__a21oi_1_113/a_29_368# sky130_fd_sc_hs__a21oi_1
Xsky130_fd_sc_hs__maj3_1_0 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__maj3_1_1/A sky130_fd_sc_hs__maj3_1_1/B
+ sky130_fd_sc_hs__maj3_1_1/X sky130_fd_sc_hs__maj3_1_1/C sky130_fd_sc_hs__maj3_1_1/a_598_384#
+ sky130_fd_sc_hs__maj3_1_1/a_226_384# sky130_fd_sc_hs__maj3_1_1/a_84_74# sky130_fd_sc_hs__maj3_1_1/a_403_136#
+ sky130_fd_sc_hs__maj3_1_1/a_406_384# sky130_fd_sc_hs__maj3_1_1/a_595_136# sky130_fd_sc_hs__maj3_1_1/a_223_120#
+ sky130_fd_sc_hs__maj3_1
Xsky130_fd_sc_hs__nand2_2_5 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__xnor2_1_3/B sky130_fd_sc_hs__nand2_2_5/B
+ sky130_fd_sc_hs__and2_2_5/X sky130_fd_sc_hs__nand2_2_5/a_27_74# sky130_fd_sc_hs__nand2_2
Xsky130_fd_sc_hs__nor2_2_1 DVSS DVDD DVDD DVSS rst sky130_fd_sc_hs__nor2_2_1/Y sky130_fd_sc_hs__nor2_2_1/A
+ sky130_fd_sc_hs__nor2_2_1/a_35_368# sky130_fd_sc_hs__nor2_2
Xsky130_fd_sc_hs__a22oi_1_19 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nor2b_1_25/Y sky130_fd_sc_hs__a32oi_1_7/A1
+ sky130_fd_sc_hs__o21a_1_27/A1 sky130_fd_sc_hs__nor2b_1_23/Y sky130_fd_sc_hs__o21a_1_25/A1
+ sky130_fd_sc_hs__a22oi_1_19/a_71_368# sky130_fd_sc_hs__a22oi_1_19/a_159_74# sky130_fd_sc_hs__a22oi_1_19/a_339_74#
+ sky130_fd_sc_hs__a22oi_1
Xsky130_fd_sc_hs__nor2_1_21 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nor2_1_21/B sky130_fd_sc_hs__nor2_1_21/Y
+ sky130_fd_sc_hs__inv_4_31/Y sky130_fd_sc_hs__nor2_1_21/a_116_368# sky130_fd_sc_hs__nor2_1
Xsky130_fd_sc_hs__nor2_1_10 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__o21a_1_5/B1 sky130_fd_sc_hs__nor2_1_11/Y
+ sky130_fd_sc_hs__inv_4_13/Y sky130_fd_sc_hs__nor2_1_11/a_116_368# sky130_fd_sc_hs__nor2_1
Xsky130_fd_sc_hs__nor2_1_65 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_73/Y sky130_fd_sc_hs__nor2_1_65/Y
+ sky130_fd_sc_hs__nor2_1_65/A sky130_fd_sc_hs__nor2_1_65/a_116_368# sky130_fd_sc_hs__nor2_1
Xsky130_fd_sc_hs__nor2_1_54 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_67/Y sky130_fd_sc_hs__nor4_1_1/B
+ sky130_fd_sc_hs__inv_4_63/A sky130_fd_sc_hs__nor2_1_55/a_116_368# sky130_fd_sc_hs__nor2_1
Xsky130_fd_sc_hs__nor2_1_43 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nor2_1_43/B sky130_fd_sc_hs__nor2_1_43/Y
+ sky130_fd_sc_hs__inv_4_67/Y sky130_fd_sc_hs__nor2_1_43/a_116_368# sky130_fd_sc_hs__nor2_1
Xsky130_fd_sc_hs__nor2_1_32 DVSS DVDD DVDD DVSS fine_control_avg_window_select[4]
+ sky130_fd_sc_hs__nor2_1_33/Y fine_control_avg_window_select[3] sky130_fd_sc_hs__nor2_1_33/a_116_368#
+ sky130_fd_sc_hs__nor2_1
Xsky130_fd_sc_hs__nor2_1_98 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nor2_1_99/B sky130_fd_sc_hs__nor2_1_99/Y
+ sky130_fd_sc_hs__nor2_1_99/A sky130_fd_sc_hs__nor2_1_99/a_116_368# sky130_fd_sc_hs__nor2_1
Xsky130_fd_sc_hs__nor2_1_87 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nor2_1_87/B sky130_fd_sc_hs__nor2_1_87/Y
+ sky130_fd_sc_hs__inv_4_81/Y sky130_fd_sc_hs__nor2_1_87/a_116_368# sky130_fd_sc_hs__nor2_1
Xsky130_fd_sc_hs__nor2_1_76 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_87/A sky130_fd_sc_hs__nor2_1_77/Y
+ sky130_fd_sc_hs__or3b_2_1/X sky130_fd_sc_hs__nor2_1_77/a_116_368# sky130_fd_sc_hs__nor2_1
.ends

.subckt sky130_fd_sc_hs__clkdlyinv5sd2_1 VNB VPB VGND VPWR A Y a_28_74# a_682_74#
+ a_549_74# a_288_74#
X0 Y a_682_74# VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X1 VGND a_549_74# a_682_74# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=420000u l=180000u
X2 VPWR a_549_74# a_682_74# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=250000u
X3 VGND A a_28_74# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4 a_549_74# a_288_74# VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=420000u l=180000u
X5 Y a_682_74# VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 VPWR A a_28_74# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X7 a_549_74# a_288_74# VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=250000u
X8 a_288_74# a_28_74# VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=250000u
X9 a_288_74# a_28_74# VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=420000u l=180000u
.ends

.subckt sky130_fd_sc_hs__o21ai_4 VNB VPB VPWR VGND Y A1 A2 B1 a_116_368# a_27_74#
X0 Y B1 a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X1 Y A2 a_116_368# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X2 Y B1 a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X3 VGND A2 a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X4 VGND A1 a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X5 a_27_74# B1 Y VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X6 a_27_74# A2 VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X7 a_27_74# B1 Y VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X8 VGND A2 a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X9 VPWR B1 Y VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X10 Y B1 VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X11 a_27_74# A1 VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X12 VPWR A1 a_116_368# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X13 a_27_74# A2 VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X14 a_116_368# A1 VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X15 VPWR A1 a_116_368# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X16 a_27_74# A1 VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X17 Y A2 a_116_368# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X18 a_116_368# A2 Y VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X19 a_116_368# A2 Y VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X20 VGND A1 a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X21 a_116_368# A1 VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
.ends

.subckt sky130_fd_sc_hs__nor4_2 VNB VPB VPWR VGND C A B D Y a_116_368# a_490_368#
+ a_27_368#
X0 VPWR A a_490_368# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X1 Y D a_116_368# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X2 VGND C Y VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X3 Y D VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X4 VGND A Y VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X5 a_490_368# B a_27_368# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X6 a_27_368# C a_116_368# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X7 a_116_368# D Y VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X8 a_27_368# B a_490_368# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X9 Y B VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X10 a_490_368# A VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X11 a_116_368# C a_27_368# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
.ends

.subckt sky130_fd_sc_hs__einvn_8 VNB VPB VPWR VGND A TE_B Z a_126_74# a_239_368# a_293_74#
X0 a_239_368# A Z VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X1 Z A a_239_368# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X2 VPWR TE_B a_239_368# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X3 a_239_368# A Z VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X4 VGND a_126_74# a_293_74# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X5 VPWR TE_B a_239_368# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X6 a_239_368# TE_B VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X7 Z A a_293_74# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X8 Z A a_239_368# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X9 a_239_368# A Z VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X10 Z A a_293_74# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X11 a_126_74# TE_B VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X12 a_293_74# a_126_74# VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X13 a_293_74# a_126_74# VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X14 a_293_74# A Z VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X15 VPWR TE_B a_239_368# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X16 a_239_368# TE_B VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X17 a_293_74# A Z VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X18 Z A a_239_368# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X19 a_239_368# TE_B VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X20 a_239_368# A Z VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X21 Z A a_239_368# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X22 a_293_74# A Z VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X23 VGND a_126_74# a_293_74# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X24 VGND a_126_74# a_293_74# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X25 a_126_74# TE_B VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X26 Z A a_293_74# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X27 VPWR TE_B a_239_368# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X28 VGND a_126_74# a_293_74# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X29 a_293_74# a_126_74# VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X30 a_239_368# TE_B VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X31 Z A a_293_74# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X32 a_293_74# A Z VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X33 a_293_74# a_126_74# VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
.ends

.subckt sky130_fd_sc_hs__mux4_4 VNB VPB VPWR VGND S1 A0 A1 A2 A3 S0 X a_1278_121#
+ a_1465_377# a_2489_347# a_114_126# a_509_392# a_296_392# a_2199_74# a_116_392# a_1285_377#
+ a_299_126# a_758_306# a_1191_121# a_1450_121#
X0 a_1191_121# a_758_306# a_1285_377# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_509_392# a_2489_347# a_2199_74# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X2 a_116_392# A1 VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 a_2199_74# a_2489_347# a_1191_121# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 a_1285_377# a_758_306# a_1191_121# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 a_1278_121# a_758_306# a_1191_121# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X6 a_2199_74# S1 a_1191_121# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X7 VGND A3 a_1450_121# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X8 a_509_392# a_758_306# a_116_392# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 a_1450_121# A3 VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X10 X a_2199_74# VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X11 a_116_392# a_758_306# a_509_392# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 VPWR A3 a_1285_377# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13 X a_2199_74# VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X14 a_1278_121# A2 VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X15 VPWR A0 a_296_392# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16 VPWR A2 a_1465_377# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17 a_1465_377# A2 VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X18 a_1191_121# a_758_306# a_1278_121# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X19 VGND S1 a_2489_347# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X20 a_1191_121# a_2489_347# a_2199_74# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X21 a_299_126# A0 VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X22 a_509_392# S0 a_114_126# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X23 a_509_392# S0 a_296_392# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X24 VGND a_2199_74# X VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X25 a_1285_377# A3 VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X26 VPWR a_2199_74# X VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X27 a_296_392# S0 a_509_392# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X28 a_114_126# S0 a_509_392# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X29 VGND a_2199_74# X VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X30 a_296_392# A0 VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X31 a_1450_121# S0 a_1191_121# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X32 X a_2199_74# VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X33 X a_2199_74# VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X34 VGND A0 a_299_126# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X35 VPWR A1 a_116_392# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X36 a_2199_74# S1 a_509_392# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X37 a_299_126# a_758_306# a_509_392# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X38 a_2199_74# a_2489_347# a_509_392# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X39 VGND A1 a_114_126# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X40 a_1191_121# S0 a_1450_121# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X41 VPWR a_2199_74# X VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X42 a_509_392# a_758_306# a_299_126# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X43 a_1191_121# S1 a_2199_74# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X44 a_114_126# A1 VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X45 VGND S0 a_758_306# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X46 VPWR S1 a_2489_347# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X47 VPWR S0 a_758_306# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X48 a_1191_121# S0 a_1465_377# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X49 a_509_392# S1 a_2199_74# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X50 a_1465_377# S0 a_1191_121# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X51 VGND A2 a_1278_121# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
.ends

.subckt sky130_fd_sc_hs__clkbuf_1 VNB VPB VPWR VGND A X a_27_74#
X0 VGND A a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1 X a_27_74# VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X2 X a_27_74# VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3 VPWR A a_27_74# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
.ends

.subckt sky130_fd_sc_hs__mux4_1 VNB VPB VPWR VGND S0 A3 A2 A1 A0 S1 X a_450_74# a_1396_99#
+ a_768_74# a_1338_125# a_763_341# a_846_74# a_27_74# a_979_74# a_264_74# a_342_74#
+ a_255_341# a_537_341# a_1065_387#
X0 a_342_74# a_27_74# a_264_74# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1 a_450_74# S0 a_342_74# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X2 VGND A1 a_450_74# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X3 a_768_74# A2 VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X4 VGND A3 a_979_74# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X5 a_1338_125# S1 a_846_74# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X6 a_846_74# S0 a_763_341# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 a_846_74# a_1396_99# a_1338_125# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 VGND S0 a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X9 VPWR S1 a_1396_99# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 X a_1338_125# VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X11 X a_1338_125# VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X12 a_763_341# A2 VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13 a_1338_125# S1 a_342_74# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14 a_342_74# a_1396_99# a_1338_125# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X15 a_264_74# A0 VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X16 VGND S1 a_1396_99# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X17 a_537_341# a_27_74# a_342_74# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X18 a_846_74# a_27_74# a_768_74# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X19 a_255_341# A0 VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X20 a_342_74# S0 a_255_341# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X21 VPWR A1 a_537_341# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X22 VPWR S0 a_27_74# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X23 a_979_74# S0 a_846_74# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X24 VPWR A3 a_1065_387# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X25 a_1065_387# a_27_74# a_846_74# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt qr_4t1_mux_top clk_Q clk_QB clk_I clk_IB din[3] din[2] din[1] din[0] rst din_2_dummy
+ din_3_dummy D1DQB_dummy D1DIB_dummy data mux_out_dummy DVSS DVDD sky130_fd_sc_hs__dfxtp_2_1/a_1172_124#
+ sky130_fd_sc_hs__dfxtp_2_3/a_1217_314# sky130_fd_sc_hs__dfxtp_4_1/a_1141_508# sky130_fd_sc_hs__dfxtp_2_3/a_695_459#
+ sky130_fd_sc_hs__dfxtp_4_3/a_651_503# sky130_fd_sc_hs__dfxtp_2_1/a_538_429# sky130_fd_sc_hs__mux4_1_1/A0
+ sky130_fd_sc_hs__mux4_1_1/a_264_74# sky130_fd_sc_hs__dfxtp_2_1/a_1217_314# sky130_fd_sc_hs__mux4_1_1/a_1338_125#
+ sky130_fd_sc_hs__mux4_4_1/a_758_306# sky130_fd_sc_hs__mux4_1_1/A2 sky130_fd_sc_hs__dfxtp_2_7/a_206_368#
+ sky130_fd_sc_hs__dfxtp_2_5/a_431_508# sky130_fd_sc_hs__mux4_1_1/A1 sky130_fd_sc_hs__dfxtp_2_7/D
+ sky130_fd_sc_hs__dfxtp_4_1/a_206_368# sky130_fd_sc_hs__dfxtp_2_7/a_708_101# sky130_fd_sc_hs__dfxtp_4_3/a_696_458#
+ sky130_fd_sc_hs__dfxtp_2_9/a_644_504# sky130_fd_sc_hs__mux4_1_1/X sky130_fd_sc_hs__dfxtp_2_11/a_206_368#
+ sky130_fd_sc_hs__dfxtp_4_1/a_437_503# sky130_fd_sc_hs__clkbuf_1_1/a_27_74# sky130_fd_sc_hs__dfxtp_2_3/a_431_508#
+ sky130_fd_sc_hs__dfxtp_4_3/a_544_485# sky130_fd_sc_hs__dfxtp_2_9/a_538_429# sky130_fd_sc_hs__dfxtp_2_11/a_708_101#
+ sky130_fd_sc_hs__dfxtp_2_11/a_1125_508# sky130_fd_sc_hs__mux4_1_1/a_27_74# sky130_fd_sc_hs__mux4_1_1/a_342_74#
+ sky130_fd_sc_hs__dfxtp_2_11/a_27_74# sky130_fd_sc_hs__dfxtp_2_1/a_695_459# sky130_fd_sc_hs__dfxtp_4_1/a_651_503#
+ sky130_fd_sc_hs__dfxtp_4_1/D sky130_fd_sc_hs__dfxtp_2_7/a_644_504# sky130_fd_sc_hs__dfxtp_4_3/a_1178_124#
+ sky130_fd_sc_hs__clkbuf_2_1/a_43_192# sky130_fd_sc_hs__dfxtp_2_5/a_206_368# sky130_fd_sc_hs__clkbuf_1_5/X
+ sky130_fd_sc_hs__dfxtp_2_9/a_1125_508# sky130_fd_sc_hs__clkbuf_2_3/X sky130_fd_sc_hs__dfxtp_2_7/a_538_429#
+ sky130_fd_sc_hs__dfxtp_2_9/Q sky130_fd_sc_hs__dfxtp_4_1/a_1178_124# sky130_fd_sc_hs__dfxtp_2_11/a_644_504#
+ sky130_fd_sc_hs__dfxtp_4_1/a_696_458# sky130_fd_sc_hs__dfxtp_2_5/a_27_74# sky130_fd_sc_hs__dfxtp_2_5/a_708_101#
+ sky130_fd_sc_hs__dfxtp_4_1/a_27_74# sky130_fd_sc_hs__mux4_4_1/a_1285_377# sky130_fd_sc_hs__dfxtp_2_7/a_1125_508#
+ sky130_fd_sc_hs__mux4_1_1/a_537_341# sky130_fd_sc_hs__mux4_1_1/a_255_341# sky130_fd_sc_hs__mux4_4_1/A0
+ sky130_fd_sc_hs__clkbuf_1_3/X sky130_fd_sc_hs__mux4_1_1/A3 sky130_fd_sc_hs__dfxtp_2_11/a_538_429#
+ sky130_fd_sc_hs__dfxtp_2_3/a_206_368# sky130_fd_sc_hs__dfxtp_2_1/a_431_508# sky130_fd_sc_hs__clkbuf_1_1/X
+ sky130_fd_sc_hs__dfxtp_2_9/a_695_459# sky130_fd_sc_hs__dfxtp_4_1/a_544_485# sky130_fd_sc_hs__dfxtp_2_5/a_1125_508#
+ sky130_fd_sc_hs__mux4_4_1/A2 sky130_fd_sc_hs__dfxtp_2_7/a_27_74# sky130_fd_sc_hs__dfxtp_2_3/a_708_101#
+ sky130_fd_sc_hs__dfxtp_2_3/a_1125_508# sky130_fd_sc_hs__dfxtp_4_3/a_27_74# sky130_fd_sc_hs__dfxtp_2_11/a_1019_424#
+ sky130_fd_sc_hs__mux4_1_1/a_450_74# sky130_fd_sc_hs__dfxtp_4_3/a_1034_424# sky130_fd_sc_hs__clkbuf_1_3/a_27_74#
+ sky130_fd_sc_hs__dfxtp_2_1/a_1125_508# sky130_fd_sc_hs__mux4_4_1/a_114_126# sky130_fd_sc_hs__dfxtp_2_1/a_27_74#
+ sky130_fd_sc_hs__dfxtp_2_5/a_644_504# sky130_fd_sc_hs__dfxtp_4_1/a_1034_424# sky130_fd_sc_hs__dfxtp_2_11/a_1172_124#
+ sky130_fd_sc_hs__mux4_4_1/a_1450_121# sky130_fd_sc_hs__dfxtp_2_9/a_431_508# sky130_fd_sc_hs__dfxtp_2_7/a_695_459#
+ sky130_fd_sc_hs__mux4_4_1/a_1191_121# sky130_fd_sc_hs__mux4_1_1/a_768_74# sky130_fd_sc_hs__dfxtp_2_5/a_538_429#
+ sky130_fd_sc_hs__dfxtp_2_9/a_1019_424# sky130_fd_sc_hs__mux4_1_1/a_1396_99# sky130_fd_sc_hs__dfxtp_2_3/a_644_504#
+ sky130_fd_sc_hs__mux4_1_1/a_1065_387# sky130_fd_sc_hs__dfxtp_4_3/a_735_102# sky130_fd_sc_hs__dfxtp_2_3/a_27_74#
+ sky130_fd_sc_hs__dfxtp_2_11/a_695_459# sky130_fd_sc_hs__dfxtp_2_11/a_1217_314# sky130_fd_sc_hs__dfxtp_2_7/a_1019_424#
+ sky130_fd_sc_hs__dfxtp_2_1/a_206_368# sky130_fd_sc_hs__mux4_4_1/a_1278_121# sky130_fd_sc_hs__dfxtp_2_3/a_538_429#
+ sky130_fd_sc_hs__dfxtp_4_3/a_1226_296# sky130_fd_sc_hs__dfxtp_2_1/a_708_101# sky130_fd_sc_hs__dfxtp_2_9/a_1172_124#
+ sky130_fd_sc_hs__mux4_4_1/a_509_392# sky130_fd_sc_hs__dfxtp_2_5/a_1019_424# sky130_fd_sc_hs__dfxtp_2_3/a_1019_424#
+ sky130_fd_sc_hs__dfxtp_2_7/a_431_508# sky130_fd_sc_hs__dfxtp_2_7/a_1172_124# sky130_fd_sc_hs__dfxtp_4_1/a_1226_296#
+ sky130_fd_sc_hs__mux4_4_1/a_1465_377# sky130_fd_sc_hs__mux4_1_1/a_846_74# sky130_fd_sc_hs__mux4_4_1/a_2199_74#
+ sky130_fd_sc_hs__dfxtp_2_9/a_1217_314# sky130_fd_sc_hs__dfxtp_4_3/a_206_368# sky130_fd_sc_hs__clkbuf_2_3/a_43_192#
+ sky130_fd_sc_hs__mux4_4_1/a_296_392# sky130_fd_sc_hs__dfxtp_2_1/a_1019_424# sky130_fd_sc_hs__dfxtp_4_3/a_437_503#
+ sky130_fd_sc_hs__dfxtp_2_11/a_431_508# sky130_fd_sc_hs__dfxtp_2_5/a_1172_124# sky130_fd_sc_hs__dfxtp_2_9/a_27_74#
+ sky130_fd_sc_hs__dfxtp_2_7/a_1217_314# sky130_fd_sc_hs__dfxtp_2_9/a_206_368# sky130_fd_sc_hs__dfxtp_2_3/a_1172_124#
+ sky130_fd_sc_hs__dfxtp_2_5/a_695_459# sky130_fd_sc_hs__mux4_4_1/a_2489_347# sky130_fd_sc_hs__mux4_1_1/a_763_341#
+ sky130_fd_sc_hs__dfxtp_4_3/a_1141_508# sky130_fd_sc_hs__mux4_4_1/a_299_126# sky130_fd_sc_hs__dfxtp_2_9/a_708_101#
+ sky130_fd_sc_hs__mux4_4_1/a_116_392# sky130_fd_sc_hs__dfxtp_2_1/a_644_504# sky130_fd_sc_hs__mux4_1_1/a_979_74#
+ sky130_fd_sc_hs__dfxtp_2_5/a_1217_314# sky130_fd_sc_hs__dfxtp_4_1/a_735_102# sky130_fd_sc_hs__clkbuf_1_5/a_27_74#
Xsky130_fd_sc_hs__clkbuf_2_3 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__clkbuf_2_3/X clk_QB
+ sky130_fd_sc_hs__clkbuf_2_3/a_43_192# sky130_fd_sc_hs__clkbuf_2
Xsky130_fd_sc_hs__dfxtp_2_1 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__mux4_4_1/A0 sky130_fd_sc_hs__clkbuf_1_1/X
+ din_2_dummy sky130_fd_sc_hs__dfxtp_2_1/a_431_508# sky130_fd_sc_hs__dfxtp_2_1/a_1125_508#
+ sky130_fd_sc_hs__dfxtp_2_1/a_206_368# sky130_fd_sc_hs__dfxtp_2_1/a_27_74# sky130_fd_sc_hs__dfxtp_2_1/a_708_101#
+ sky130_fd_sc_hs__dfxtp_2_1/a_1019_424# sky130_fd_sc_hs__dfxtp_2_1/a_1172_124# sky130_fd_sc_hs__dfxtp_2_1/a_644_504#
+ sky130_fd_sc_hs__dfxtp_2_1/a_1217_314# sky130_fd_sc_hs__dfxtp_2_1/a_538_429# sky130_fd_sc_hs__dfxtp_2_1/a_695_459#
+ sky130_fd_sc_hs__dfxtp_2
Xsky130_fd_sc_hs__mux4_4_0 DVSS DVDD DVDD DVSS clk_IB sky130_fd_sc_hs__mux4_4_1/A0
+ D1DQB_dummy sky130_fd_sc_hs__mux4_4_1/A2 D1DIB_dummy clk_QB mux_out_dummy sky130_fd_sc_hs__mux4_4_1/a_1278_121#
+ sky130_fd_sc_hs__mux4_4_1/a_1465_377# sky130_fd_sc_hs__mux4_4_1/a_2489_347# sky130_fd_sc_hs__mux4_4_1/a_114_126#
+ sky130_fd_sc_hs__mux4_4_1/a_509_392# sky130_fd_sc_hs__mux4_4_1/a_296_392# sky130_fd_sc_hs__mux4_4_1/a_2199_74#
+ sky130_fd_sc_hs__mux4_4_1/a_116_392# sky130_fd_sc_hs__mux4_4_1/a_1285_377# sky130_fd_sc_hs__mux4_4_1/a_299_126#
+ sky130_fd_sc_hs__mux4_4_1/a_758_306# sky130_fd_sc_hs__mux4_4_1/a_1191_121# sky130_fd_sc_hs__mux4_4_1/a_1450_121#
+ sky130_fd_sc_hs__mux4_4
Xsky130_fd_sc_hs__dfxtp_2_10 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__dfxtp_2_7/D sky130_fd_sc_hs__clkbuf_1_5/X
+ din[0] sky130_fd_sc_hs__dfxtp_2_11/a_431_508# sky130_fd_sc_hs__dfxtp_2_11/a_1125_508#
+ sky130_fd_sc_hs__dfxtp_2_11/a_206_368# sky130_fd_sc_hs__dfxtp_2_11/a_27_74# sky130_fd_sc_hs__dfxtp_2_11/a_708_101#
+ sky130_fd_sc_hs__dfxtp_2_11/a_1019_424# sky130_fd_sc_hs__dfxtp_2_11/a_1172_124#
+ sky130_fd_sc_hs__dfxtp_2_11/a_644_504# sky130_fd_sc_hs__dfxtp_2_11/a_1217_314# sky130_fd_sc_hs__dfxtp_2_11/a_538_429#
+ sky130_fd_sc_hs__dfxtp_2_11/a_695_459# sky130_fd_sc_hs__dfxtp_2
Xsky130_fd_sc_hs__dfxtp_2_2 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__mux4_4_1/A2 sky130_fd_sc_hs__clkbuf_2_3/X
+ din_3_dummy sky130_fd_sc_hs__dfxtp_2_3/a_431_508# sky130_fd_sc_hs__dfxtp_2_3/a_1125_508#
+ sky130_fd_sc_hs__dfxtp_2_3/a_206_368# sky130_fd_sc_hs__dfxtp_2_3/a_27_74# sky130_fd_sc_hs__dfxtp_2_3/a_708_101#
+ sky130_fd_sc_hs__dfxtp_2_3/a_1019_424# sky130_fd_sc_hs__dfxtp_2_3/a_1172_124# sky130_fd_sc_hs__dfxtp_2_3/a_644_504#
+ sky130_fd_sc_hs__dfxtp_2_3/a_1217_314# sky130_fd_sc_hs__dfxtp_2_3/a_538_429# sky130_fd_sc_hs__dfxtp_2_3/a_695_459#
+ sky130_fd_sc_hs__dfxtp_2
Xsky130_fd_sc_hs__mux4_4_1 DVSS DVDD DVDD DVSS clk_IB sky130_fd_sc_hs__mux4_4_1/A0
+ D1DQB_dummy sky130_fd_sc_hs__mux4_4_1/A2 D1DIB_dummy clk_QB mux_out_dummy sky130_fd_sc_hs__mux4_4_1/a_1278_121#
+ sky130_fd_sc_hs__mux4_4_1/a_1465_377# sky130_fd_sc_hs__mux4_4_1/a_2489_347# sky130_fd_sc_hs__mux4_4_1/a_114_126#
+ sky130_fd_sc_hs__mux4_4_1/a_509_392# sky130_fd_sc_hs__mux4_4_1/a_296_392# sky130_fd_sc_hs__mux4_4_1/a_2199_74#
+ sky130_fd_sc_hs__mux4_4_1/a_116_392# sky130_fd_sc_hs__mux4_4_1/a_1285_377# sky130_fd_sc_hs__mux4_4_1/a_299_126#
+ sky130_fd_sc_hs__mux4_4_1/a_758_306# sky130_fd_sc_hs__mux4_4_1/a_1191_121# sky130_fd_sc_hs__mux4_4_1/a_1450_121#
+ sky130_fd_sc_hs__mux4_4
Xsky130_fd_sc_hs__dfxtp_2_11 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__dfxtp_2_7/D sky130_fd_sc_hs__clkbuf_1_5/X
+ din[0] sky130_fd_sc_hs__dfxtp_2_11/a_431_508# sky130_fd_sc_hs__dfxtp_2_11/a_1125_508#
+ sky130_fd_sc_hs__dfxtp_2_11/a_206_368# sky130_fd_sc_hs__dfxtp_2_11/a_27_74# sky130_fd_sc_hs__dfxtp_2_11/a_708_101#
+ sky130_fd_sc_hs__dfxtp_2_11/a_1019_424# sky130_fd_sc_hs__dfxtp_2_11/a_1172_124#
+ sky130_fd_sc_hs__dfxtp_2_11/a_644_504# sky130_fd_sc_hs__dfxtp_2_11/a_1217_314# sky130_fd_sc_hs__dfxtp_2_11/a_538_429#
+ sky130_fd_sc_hs__dfxtp_2_11/a_695_459# sky130_fd_sc_hs__dfxtp_2
Xsky130_fd_sc_hs__dfxtp_2_3 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__mux4_4_1/A2 sky130_fd_sc_hs__clkbuf_2_3/X
+ din_3_dummy sky130_fd_sc_hs__dfxtp_2_3/a_431_508# sky130_fd_sc_hs__dfxtp_2_3/a_1125_508#
+ sky130_fd_sc_hs__dfxtp_2_3/a_206_368# sky130_fd_sc_hs__dfxtp_2_3/a_27_74# sky130_fd_sc_hs__dfxtp_2_3/a_708_101#
+ sky130_fd_sc_hs__dfxtp_2_3/a_1019_424# sky130_fd_sc_hs__dfxtp_2_3/a_1172_124# sky130_fd_sc_hs__dfxtp_2_3/a_644_504#
+ sky130_fd_sc_hs__dfxtp_2_3/a_1217_314# sky130_fd_sc_hs__dfxtp_2_3/a_538_429# sky130_fd_sc_hs__dfxtp_2_3/a_695_459#
+ sky130_fd_sc_hs__dfxtp_2
Xsky130_fd_sc_hs__dfxtp_2_4 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__mux4_1_1/A1 sky130_fd_sc_hs__clkbuf_2_3/X
+ sky130_fd_sc_hs__dfxtp_2_9/Q sky130_fd_sc_hs__dfxtp_2_5/a_431_508# sky130_fd_sc_hs__dfxtp_2_5/a_1125_508#
+ sky130_fd_sc_hs__dfxtp_2_5/a_206_368# sky130_fd_sc_hs__dfxtp_2_5/a_27_74# sky130_fd_sc_hs__dfxtp_2_5/a_708_101#
+ sky130_fd_sc_hs__dfxtp_2_5/a_1019_424# sky130_fd_sc_hs__dfxtp_2_5/a_1172_124# sky130_fd_sc_hs__dfxtp_2_5/a_644_504#
+ sky130_fd_sc_hs__dfxtp_2_5/a_1217_314# sky130_fd_sc_hs__dfxtp_2_5/a_538_429# sky130_fd_sc_hs__dfxtp_2_5/a_695_459#
+ sky130_fd_sc_hs__dfxtp_2
Xsky130_fd_sc_hs__dfxtp_2_5 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__mux4_1_1/A1 sky130_fd_sc_hs__clkbuf_2_3/X
+ sky130_fd_sc_hs__dfxtp_2_9/Q sky130_fd_sc_hs__dfxtp_2_5/a_431_508# sky130_fd_sc_hs__dfxtp_2_5/a_1125_508#
+ sky130_fd_sc_hs__dfxtp_2_5/a_206_368# sky130_fd_sc_hs__dfxtp_2_5/a_27_74# sky130_fd_sc_hs__dfxtp_2_5/a_708_101#
+ sky130_fd_sc_hs__dfxtp_2_5/a_1019_424# sky130_fd_sc_hs__dfxtp_2_5/a_1172_124# sky130_fd_sc_hs__dfxtp_2_5/a_644_504#
+ sky130_fd_sc_hs__dfxtp_2_5/a_1217_314# sky130_fd_sc_hs__dfxtp_2_5/a_538_429# sky130_fd_sc_hs__dfxtp_2_5/a_695_459#
+ sky130_fd_sc_hs__dfxtp_2
Xsky130_fd_sc_hs__dfxtp_2_6 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__mux4_1_1/A3 sky130_fd_sc_hs__clkbuf_1_1/X
+ sky130_fd_sc_hs__dfxtp_2_7/D sky130_fd_sc_hs__dfxtp_2_7/a_431_508# sky130_fd_sc_hs__dfxtp_2_7/a_1125_508#
+ sky130_fd_sc_hs__dfxtp_2_7/a_206_368# sky130_fd_sc_hs__dfxtp_2_7/a_27_74# sky130_fd_sc_hs__dfxtp_2_7/a_708_101#
+ sky130_fd_sc_hs__dfxtp_2_7/a_1019_424# sky130_fd_sc_hs__dfxtp_2_7/a_1172_124# sky130_fd_sc_hs__dfxtp_2_7/a_644_504#
+ sky130_fd_sc_hs__dfxtp_2_7/a_1217_314# sky130_fd_sc_hs__dfxtp_2_7/a_538_429# sky130_fd_sc_hs__dfxtp_2_7/a_695_459#
+ sky130_fd_sc_hs__dfxtp_2
Xsky130_fd_sc_hs__dfxtp_2_7 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__mux4_1_1/A3 sky130_fd_sc_hs__clkbuf_1_1/X
+ sky130_fd_sc_hs__dfxtp_2_7/D sky130_fd_sc_hs__dfxtp_2_7/a_431_508# sky130_fd_sc_hs__dfxtp_2_7/a_1125_508#
+ sky130_fd_sc_hs__dfxtp_2_7/a_206_368# sky130_fd_sc_hs__dfxtp_2_7/a_27_74# sky130_fd_sc_hs__dfxtp_2_7/a_708_101#
+ sky130_fd_sc_hs__dfxtp_2_7/a_1019_424# sky130_fd_sc_hs__dfxtp_2_7/a_1172_124# sky130_fd_sc_hs__dfxtp_2_7/a_644_504#
+ sky130_fd_sc_hs__dfxtp_2_7/a_1217_314# sky130_fd_sc_hs__dfxtp_2_7/a_538_429# sky130_fd_sc_hs__dfxtp_2_7/a_695_459#
+ sky130_fd_sc_hs__dfxtp_2
Xsky130_fd_sc_hs__dfxtp_2_8 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__dfxtp_2_9/Q sky130_fd_sc_hs__clkbuf_1_3/X
+ din[1] sky130_fd_sc_hs__dfxtp_2_9/a_431_508# sky130_fd_sc_hs__dfxtp_2_9/a_1125_508#
+ sky130_fd_sc_hs__dfxtp_2_9/a_206_368# sky130_fd_sc_hs__dfxtp_2_9/a_27_74# sky130_fd_sc_hs__dfxtp_2_9/a_708_101#
+ sky130_fd_sc_hs__dfxtp_2_9/a_1019_424# sky130_fd_sc_hs__dfxtp_2_9/a_1172_124# sky130_fd_sc_hs__dfxtp_2_9/a_644_504#
+ sky130_fd_sc_hs__dfxtp_2_9/a_1217_314# sky130_fd_sc_hs__dfxtp_2_9/a_538_429# sky130_fd_sc_hs__dfxtp_2_9/a_695_459#
+ sky130_fd_sc_hs__dfxtp_2
Xsky130_fd_sc_hs__dfxtp_2_9 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__dfxtp_2_9/Q sky130_fd_sc_hs__clkbuf_1_3/X
+ din[1] sky130_fd_sc_hs__dfxtp_2_9/a_431_508# sky130_fd_sc_hs__dfxtp_2_9/a_1125_508#
+ sky130_fd_sc_hs__dfxtp_2_9/a_206_368# sky130_fd_sc_hs__dfxtp_2_9/a_27_74# sky130_fd_sc_hs__dfxtp_2_9/a_708_101#
+ sky130_fd_sc_hs__dfxtp_2_9/a_1019_424# sky130_fd_sc_hs__dfxtp_2_9/a_1172_124# sky130_fd_sc_hs__dfxtp_2_9/a_644_504#
+ sky130_fd_sc_hs__dfxtp_2_9/a_1217_314# sky130_fd_sc_hs__dfxtp_2_9/a_538_429# sky130_fd_sc_hs__dfxtp_2_9/a_695_459#
+ sky130_fd_sc_hs__dfxtp_2
Xsky130_fd_sc_hs__clkbuf_1_0 DVSS DVDD DVDD DVSS clk_IB sky130_fd_sc_hs__clkbuf_1_1/X
+ sky130_fd_sc_hs__clkbuf_1_1/a_27_74# sky130_fd_sc_hs__clkbuf_1
Xsky130_fd_sc_hs__clkbuf_1_1 DVSS DVDD DVDD DVSS clk_IB sky130_fd_sc_hs__clkbuf_1_1/X
+ sky130_fd_sc_hs__clkbuf_1_1/a_27_74# sky130_fd_sc_hs__clkbuf_1
Xsky130_fd_sc_hs__clkbuf_1_2 DVSS DVDD DVDD DVSS clk_Q sky130_fd_sc_hs__clkbuf_1_3/X
+ sky130_fd_sc_hs__clkbuf_1_3/a_27_74# sky130_fd_sc_hs__clkbuf_1
Xsky130_fd_sc_hs__clkbuf_1_3 DVSS DVDD DVDD DVSS clk_Q sky130_fd_sc_hs__clkbuf_1_3/X
+ sky130_fd_sc_hs__clkbuf_1_3/a_27_74# sky130_fd_sc_hs__clkbuf_1
Xsky130_fd_sc_hs__clkbuf_1_4 DVSS DVDD DVDD DVSS clk_I sky130_fd_sc_hs__clkbuf_1_5/X
+ sky130_fd_sc_hs__clkbuf_1_5/a_27_74# sky130_fd_sc_hs__clkbuf_1
Xsky130_fd_sc_hs__clkbuf_1_5 DVSS DVDD DVDD DVSS clk_I sky130_fd_sc_hs__clkbuf_1_5/X
+ sky130_fd_sc_hs__clkbuf_1_5/a_27_74# sky130_fd_sc_hs__clkbuf_1
Xsky130_fd_sc_hs__mux4_1_0 DVSS DVDD DVDD DVSS clk_Q sky130_fd_sc_hs__mux4_1_1/A3
+ sky130_fd_sc_hs__mux4_1_1/A2 sky130_fd_sc_hs__mux4_1_1/A1 sky130_fd_sc_hs__mux4_1_1/A0
+ clk_I sky130_fd_sc_hs__mux4_1_1/X sky130_fd_sc_hs__mux4_1_1/a_450_74# sky130_fd_sc_hs__mux4_1_1/a_1396_99#
+ sky130_fd_sc_hs__mux4_1_1/a_768_74# sky130_fd_sc_hs__mux4_1_1/a_1338_125# sky130_fd_sc_hs__mux4_1_1/a_763_341#
+ sky130_fd_sc_hs__mux4_1_1/a_846_74# sky130_fd_sc_hs__mux4_1_1/a_27_74# sky130_fd_sc_hs__mux4_1_1/a_979_74#
+ sky130_fd_sc_hs__mux4_1_1/a_264_74# sky130_fd_sc_hs__mux4_1_1/a_342_74# sky130_fd_sc_hs__mux4_1_1/a_255_341#
+ sky130_fd_sc_hs__mux4_1_1/a_537_341# sky130_fd_sc_hs__mux4_1_1/a_1065_387# sky130_fd_sc_hs__mux4_1
Xsky130_fd_sc_hs__mux4_1_1 DVSS DVDD DVDD DVSS clk_Q sky130_fd_sc_hs__mux4_1_1/A3
+ sky130_fd_sc_hs__mux4_1_1/A2 sky130_fd_sc_hs__mux4_1_1/A1 sky130_fd_sc_hs__mux4_1_1/A0
+ clk_I sky130_fd_sc_hs__mux4_1_1/X sky130_fd_sc_hs__mux4_1_1/a_450_74# sky130_fd_sc_hs__mux4_1_1/a_1396_99#
+ sky130_fd_sc_hs__mux4_1_1/a_768_74# sky130_fd_sc_hs__mux4_1_1/a_1338_125# sky130_fd_sc_hs__mux4_1_1/a_763_341#
+ sky130_fd_sc_hs__mux4_1_1/a_846_74# sky130_fd_sc_hs__mux4_1_1/a_27_74# sky130_fd_sc_hs__mux4_1_1/a_979_74#
+ sky130_fd_sc_hs__mux4_1_1/a_264_74# sky130_fd_sc_hs__mux4_1_1/a_342_74# sky130_fd_sc_hs__mux4_1_1/a_255_341#
+ sky130_fd_sc_hs__mux4_1_1/a_537_341# sky130_fd_sc_hs__mux4_1_1/a_1065_387# sky130_fd_sc_hs__mux4_1
Xsky130_fd_sc_hs__clkinv_4_0 DVSS DVDD DVDD DVSS data sky130_fd_sc_hs__mux4_1_1/X
+ sky130_fd_sc_hs__clkinv_4
Xsky130_fd_sc_hs__clkinv_4_1 DVSS DVDD DVDD DVSS data sky130_fd_sc_hs__mux4_1_1/X
+ sky130_fd_sc_hs__clkinv_4
Xsky130_fd_sc_hs__dfxtp_4_0 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__mux4_1_1/A2 sky130_fd_sc_hs__dfxtp_4_1/D
+ sky130_fd_sc_hs__clkbuf_1_3/X sky130_fd_sc_hs__dfxtp_4_1/a_1226_296# sky130_fd_sc_hs__dfxtp_4_1/a_735_102#
+ sky130_fd_sc_hs__dfxtp_4_1/a_1141_508# sky130_fd_sc_hs__dfxtp_4_1/a_206_368# sky130_fd_sc_hs__dfxtp_4_1/a_437_503#
+ sky130_fd_sc_hs__dfxtp_4_1/a_27_74# sky130_fd_sc_hs__dfxtp_4_1/a_651_503# sky130_fd_sc_hs__dfxtp_4_1/a_696_458#
+ sky130_fd_sc_hs__dfxtp_4_1/a_544_485# sky130_fd_sc_hs__dfxtp_4_1/a_1178_124# sky130_fd_sc_hs__dfxtp_4_1/a_1034_424#
+ sky130_fd_sc_hs__dfxtp_4
Xsky130_fd_sc_hs__clkbuf_2_0 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__dfxtp_4_1/D din[3]
+ sky130_fd_sc_hs__clkbuf_2_1/a_43_192# sky130_fd_sc_hs__clkbuf_2
Xsky130_fd_sc_hs__dfxtp_4_1 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__mux4_1_1/A2 sky130_fd_sc_hs__dfxtp_4_1/D
+ sky130_fd_sc_hs__clkbuf_1_3/X sky130_fd_sc_hs__dfxtp_4_1/a_1226_296# sky130_fd_sc_hs__dfxtp_4_1/a_735_102#
+ sky130_fd_sc_hs__dfxtp_4_1/a_1141_508# sky130_fd_sc_hs__dfxtp_4_1/a_206_368# sky130_fd_sc_hs__dfxtp_4_1/a_437_503#
+ sky130_fd_sc_hs__dfxtp_4_1/a_27_74# sky130_fd_sc_hs__dfxtp_4_1/a_651_503# sky130_fd_sc_hs__dfxtp_4_1/a_696_458#
+ sky130_fd_sc_hs__dfxtp_4_1/a_544_485# sky130_fd_sc_hs__dfxtp_4_1/a_1178_124# sky130_fd_sc_hs__dfxtp_4_1/a_1034_424#
+ sky130_fd_sc_hs__dfxtp_4
Xsky130_fd_sc_hs__clkbuf_2_1 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__dfxtp_4_1/D din[3]
+ sky130_fd_sc_hs__clkbuf_2_1/a_43_192# sky130_fd_sc_hs__clkbuf_2
Xsky130_fd_sc_hs__dfxtp_4_2 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__mux4_1_1/A0 din[2]
+ sky130_fd_sc_hs__clkbuf_1_5/X sky130_fd_sc_hs__dfxtp_4_3/a_1226_296# sky130_fd_sc_hs__dfxtp_4_3/a_735_102#
+ sky130_fd_sc_hs__dfxtp_4_3/a_1141_508# sky130_fd_sc_hs__dfxtp_4_3/a_206_368# sky130_fd_sc_hs__dfxtp_4_3/a_437_503#
+ sky130_fd_sc_hs__dfxtp_4_3/a_27_74# sky130_fd_sc_hs__dfxtp_4_3/a_651_503# sky130_fd_sc_hs__dfxtp_4_3/a_696_458#
+ sky130_fd_sc_hs__dfxtp_4_3/a_544_485# sky130_fd_sc_hs__dfxtp_4_3/a_1178_124# sky130_fd_sc_hs__dfxtp_4_3/a_1034_424#
+ sky130_fd_sc_hs__dfxtp_4
Xsky130_fd_sc_hs__clkbuf_2_2 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__clkbuf_2_3/X clk_QB
+ sky130_fd_sc_hs__clkbuf_2_3/a_43_192# sky130_fd_sc_hs__clkbuf_2
Xsky130_fd_sc_hs__dfxtp_2_0 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__mux4_4_1/A0 sky130_fd_sc_hs__clkbuf_1_1/X
+ din_2_dummy sky130_fd_sc_hs__dfxtp_2_1/a_431_508# sky130_fd_sc_hs__dfxtp_2_1/a_1125_508#
+ sky130_fd_sc_hs__dfxtp_2_1/a_206_368# sky130_fd_sc_hs__dfxtp_2_1/a_27_74# sky130_fd_sc_hs__dfxtp_2_1/a_708_101#
+ sky130_fd_sc_hs__dfxtp_2_1/a_1019_424# sky130_fd_sc_hs__dfxtp_2_1/a_1172_124# sky130_fd_sc_hs__dfxtp_2_1/a_644_504#
+ sky130_fd_sc_hs__dfxtp_2_1/a_1217_314# sky130_fd_sc_hs__dfxtp_2_1/a_538_429# sky130_fd_sc_hs__dfxtp_2_1/a_695_459#
+ sky130_fd_sc_hs__dfxtp_2
Xsky130_fd_sc_hs__dfxtp_4_3 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__mux4_1_1/A0 din[2]
+ sky130_fd_sc_hs__clkbuf_1_5/X sky130_fd_sc_hs__dfxtp_4_3/a_1226_296# sky130_fd_sc_hs__dfxtp_4_3/a_735_102#
+ sky130_fd_sc_hs__dfxtp_4_3/a_1141_508# sky130_fd_sc_hs__dfxtp_4_3/a_206_368# sky130_fd_sc_hs__dfxtp_4_3/a_437_503#
+ sky130_fd_sc_hs__dfxtp_4_3/a_27_74# sky130_fd_sc_hs__dfxtp_4_3/a_651_503# sky130_fd_sc_hs__dfxtp_4_3/a_696_458#
+ sky130_fd_sc_hs__dfxtp_4_3/a_544_485# sky130_fd_sc_hs__dfxtp_4_3/a_1178_124# sky130_fd_sc_hs__dfxtp_4_3/a_1034_424#
+ sky130_fd_sc_hs__dfxtp_4
.ends

.subckt sky130_fd_sc_hs__buf_1 VNB VPB VPWR VGND A X a_27_164#
X0 X a_27_164# VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X1 X a_27_164# VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X2 VPWR A a_27_164# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X3 VGND A a_27_164# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=550000u l=150000u
.ends

.subckt sky130_fd_sc_hs__einvp_4 VNB VPB VPWR VGND TE Z A a_27_74# a_27_368# a_473_323#
X0 VPWR TE a_473_323# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X1 Z A a_27_368# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X2 Z A a_27_368# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X3 a_27_74# A Z VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X4 a_27_74# TE VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X5 Z A a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X6 Z A a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X7 a_27_368# A Z VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X8 VPWR a_473_323# a_27_368# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X9 a_27_368# a_473_323# VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X10 VGND TE a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X11 a_27_368# a_473_323# VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X12 VPWR a_473_323# a_27_368# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X13 a_27_74# A Z VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X14 a_27_74# TE VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X15 VGND TE a_473_323# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X16 VGND TE a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X17 a_27_368# A Z VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
.ends

.subckt sky130_fd_sc_hs__dlygate4sd3_1 VNB VPB VGND VPWR A X a_405_138# a_28_74# a_289_74#
X0 X a_405_138# VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X1 VGND A a_28_74# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 VPWR a_289_74# a_405_138# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X3 VGND a_289_74# a_405_138# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=420000u l=180000u
X4 X a_405_138# VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X5 a_289_74# a_28_74# VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X6 a_289_74# a_28_74# VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=420000u l=180000u
X7 VPWR A a_28_74# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
.ends

.subckt sky130_fd_sc_hs__inv_16 VNB VPB VPWR VGND Y A
X0 VPWR A Y VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X1 Y A VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X2 Y A VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X3 VGND A Y VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X4 VGND A Y VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X5 Y A VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X6 VPWR A Y VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X7 VPWR A Y VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X8 VGND A Y VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X9 Y A VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X10 Y A VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X11 VGND A Y VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X12 Y A VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X13 VPWR A Y VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X14 Y A VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X15 VPWR A Y VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X16 VGND A Y VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X17 Y A VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X18 VPWR A Y VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X19 Y A VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X20 VPWR A Y VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X21 VGND A Y VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X22 Y A VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X23 VGND A Y VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X24 Y A VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X25 VGND A Y VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X26 Y A VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X27 VPWR A Y VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X28 Y A VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X29 Y A VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X30 Y A VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X31 Y A VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
.ends

.subckt sky130_fd_sc_hs__einvp_1 VNB VPB VPWR VGND TE Z A a_44_549# a_318_74# a_310_392#
X0 a_310_392# a_44_549# VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 VGND TE a_44_549# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 VPWR TE a_44_549# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3 a_318_74# TE VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X4 Z A a_318_74# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X5 Z A a_310_392# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_sc_hs__nand2_8 VNB VPB VPWR VGND B A Y a_27_74#
X0 Y A VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X1 Y A a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X2 VPWR A Y VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X3 a_27_74# B VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X4 Y A VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X5 VPWR B Y VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X6 Y A a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X7 VGND B a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X8 VGND B a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X9 a_27_74# B VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X10 a_27_74# A Y VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X11 Y A a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X12 Y B VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X13 a_27_74# B VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X14 a_27_74# B VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X15 a_27_74# A Y VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X16 a_27_74# A Y VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X17 VPWR A Y VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X18 VPWR B Y VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X19 a_27_74# A Y VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X20 Y B VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X21 VGND B a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X22 VGND B a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X23 Y A a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
.ends

.subckt sky130_fd_sc_hs__and4_2 VNB VPB VPWR VGND D C B A X a_335_74# a_143_74# a_221_74#
+ a_56_74#
X0 a_221_74# B a_143_74# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X1 VGND a_56_74# X VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X2 VPWR a_56_74# X VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X3 a_56_74# A VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 X a_56_74# VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X5 VPWR D a_56_74# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 a_56_74# C VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 a_143_74# A a_56_74# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X8 VGND D a_335_74# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X9 a_335_74# C a_221_74# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X10 VPWR B a_56_74# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 X a_56_74# VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
.ends

.subckt sky130_fd_sc_hs__inv_1 VNB VPB VPWR VGND Y A
X0 Y A VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X1 Y A VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
.ends

.subckt sky130_fd_sc_hs__nand3_4 VNB VPB VPWR VGND C B A Y a_456_82# a_27_82#
X0 VGND C a_456_82# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X1 a_27_82# A Y VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X2 Y A a_27_82# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X3 VGND C a_456_82# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X4 a_27_82# B a_456_82# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X5 a_27_82# B a_456_82# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X6 VPWR B Y VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X7 a_456_82# C VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X8 a_27_82# A Y VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X9 Y B VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X10 a_456_82# B a_27_82# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X11 VPWR C Y VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X12 a_456_82# B a_27_82# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X13 Y C VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X14 a_456_82# C VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X15 VPWR A Y VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X16 Y A a_27_82# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X17 Y A VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
.ends

.subckt sky130_fd_sc_hs__inv_8 VNB VPB VPWR VGND A Y
X0 Y A VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X1 VPWR A Y VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X2 Y A VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X3 Y A VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X4 VPWR A Y VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X5 Y A VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X6 VGND A Y VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X7 VGND A Y VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X8 VPWR A Y VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X9 VGND A Y VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X10 Y A VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X11 Y A VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X12 VPWR A Y VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X13 Y A VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X14 VGND A Y VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X15 Y A VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
.ends

.subckt sky130_fd_sc_hs__dlygate4sd2_1 VNB VPB VGND VPWR A X a_405_138# a_28_74# a_288_74#
X0 X a_405_138# VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X1 VPWR a_288_74# a_405_138# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=250000u
X2 VGND A a_28_74# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3 VGND a_288_74# a_405_138# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=420000u l=180000u
X4 X a_405_138# VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X5 a_288_74# a_28_74# VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=250000u
X6 VPWR A a_28_74# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7 a_288_74# a_28_74# VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=420000u l=180000u
.ends

.subckt sky130_fd_sc_hs__bufbuf_8 VNB VPB VPWR VGND A X a_334_368# a_27_112# a_221_368#
X0 VGND a_334_368# X VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X1 X a_334_368# VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X2 a_221_368# a_27_112# VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X3 VPWR a_334_368# X VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X4 a_221_368# a_27_112# VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X5 X a_334_368# VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X6 VGND a_221_368# a_334_368# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X7 VPWR a_334_368# X VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X8 VPWR a_334_368# X VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X9 X a_334_368# VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X10 X a_334_368# VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X11 VPWR a_334_368# X VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X12 VGND a_334_368# X VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X13 X a_334_368# VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X14 X a_334_368# VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X15 X a_334_368# VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X16 VGND a_334_368# X VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X17 VGND a_221_368# a_334_368# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X18 X a_334_368# VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X19 VPWR a_221_368# a_334_368# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X20 VGND A a_27_112# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=550000u l=150000u
X21 a_334_368# a_221_368# VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X22 VGND a_334_368# X VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X23 VPWR a_221_368# a_334_368# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X24 a_334_368# a_221_368# VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X25 VPWR A a_27_112# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
.ends

.subckt sky130_fd_sc_hs__buf_4 VNB VPB VPWR VGND A X a_86_260#
X0 a_86_260# A VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X1 VPWR a_86_260# X VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X2 X a_86_260# VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X3 VPWR a_86_260# X VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X4 VGND a_86_260# X VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X5 X a_86_260# VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X6 X a_86_260# VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X7 X a_86_260# VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X8 VGND a_86_260# X VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X9 VPWR A a_86_260# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X10 a_86_260# A VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
.ends

.subckt osc_core glob_en delay_con_lsb[4] delay_con_lsb[3] delay_con_lsb[2] delay_con_lsb[1]
+ delay_con_lsb[0] delay_con_msb[7] delay_con_msb[6] delay_con_msb[5] delay_con_msb[4]
+ delay_con_msb[3] delay_con_msb[2] delay_con_msb[1] delay_con_msb[0] con_perb_1[3]
+ con_perb_1[2] con_perb_1[1] con_perb_1[0] con_perb_2[3] con_perb_2[2] con_perb_2[1]
+ con_perb_2[0] con_perb_3[3] con_perb_3[2] con_perb_3[1] con_perb_3[0] con_perb_4[3]
+ con_perb_4[2] con_perb_4[1] con_perb_4[0] con_perb_5[3] con_perb_5[2] con_perb_5[1]
+ con_perb_5[0] ref_clk pi1_l[3] pi1_l[2] pi1_l[1] pi1_l[0] pi1_r[3] pi1_r[2] pi1_r[1]
+ pi1_r[0] pi2_l[3] pi2_l[2] pi2_l[1] pi2_l[0] pi2_r[3] pi2_r[2] pi2_r[1] pi2_r[0]
+ pi3_l[3] pi3_l[2] pi3_l[1] pi3_l[0] pi3_r[3] pi3_r[2] pi3_r[1] pi3_r[0] pi4_l[3]
+ pi4_l[2] pi4_l[1] pi4_l[0] pi4_r[3] pi4_r[2] pi4_r[1] pi4_r[0] pi5_l[3] pi5_l[2]
+ pi5_l[1] pi5_l[0] pi5_r[3] pi5_r[2] pi5_r[1] pi5_r[0] osc_000 osc_036 osc_072 osc_108
+ osc_144 inj_en inj_out osc_hold p1 p2 p3 p4 p5 DVSS DVDD sky130_fd_sc_hs__einvp_2_5/a_36_74#
+ sky130_fd_sc_hs__dlygate4sd3_1_75/X sky130_fd_sc_hs__nand2_2_93/Y sky130_fd_sc_hs__dlygate4sd3_1_1/X
+ sky130_fd_sc_hs__dlygate4sd3_1_11/a_28_74# sky130_fd_sc_hs__inv_4_5/Y sky130_fd_sc_hs__dlygate4sd3_1_27/a_289_74#
+ sky130_fd_sc_hs__nand2_8_9/B sky130_fd_sc_hs__dlygate4sd3_1_7/a_405_138# sky130_fd_sc_hs__nand2_4_40/a_27_74#
+ sky130_fd_sc_hs__dfrtp_4_3/a_890_138# sky130_fd_sc_hs__nand2_1_9/B sky130_fd_sc_hs__nand2_4_137/a_27_74#
+ sky130_fd_sc_hs__dlygate4sd3_1_56/A sky130_fd_sc_hs__inv_4_17/Y sky130_fd_sc_hs__nand2_2_55/Y
+ sky130_fd_sc_hs__nand2_8_31/a_27_74# sky130_fd_sc_hs__nand2_4_53/a_27_74# sky130_fd_sc_hs__nand2_4_123/Y
+ sky130_fd_sc_hs__einvp_1_1/a_44_549# sky130_fd_sc_hs__nand2_1_5/a_117_74# sky130_fd_sc_hs__inv_4_3/Y
+ sky130_fd_sc_hs__nand2_2_69/a_27_74# sky130_fd_sc_hs__einvp_2_11/a_263_323# sky130_fd_sc_hs__einvp_8_3/a_27_368#
+ sky130_fd_sc_hs__nand2_2_84/B sky130_fd_sc_hs__a21oi_1_9/a_29_368# sky130_fd_sc_hs__nand2_4_51/Y
+ sky130_fd_sc_hs__dlygate4sd3_1_68/X sky130_fd_sc_hs__einvp_4_9/a_473_323# sky130_fd_sc_hs__nand2_2_109/a_27_74#
+ sky130_fd_sc_hs__inv_16_3/Y sky130_fd_sc_hs__dlygate4sd3_1_31/X sky130_fd_sc_hs__dlygate4sd3_1_5/A
+ sky130_fd_sc_hs__nand2_2_45/B sky130_fd_sc_hs__nand2_2_3/a_27_74# sky130_fd_sc_hs__einvp_8_14/a_802_323#
+ sky130_fd_sc_hs__einvp_2_19/a_36_74# sky130_fd_sc_hs__nand2_4_15/Y sky130_fd_sc_hs__nand2_4_153/Y
+ sky130_fd_sc_hs__nand2_4_107/a_27_74# sky130_fd_sc_hs__and4_2_3/X sky130_fd_sc_hs__and2_2_1/a_118_74#
+ sky130_fd_sc_hs__nand2_4_93/a_27_74# sky130_fd_sc_hs__einvp_1_5/a_44_549# sky130_fd_sc_hs__nand2_1_9/a_117_74#
+ sky130_fd_sc_hs__and4_2_3/a_335_74# sky130_fd_sc_hs__a21oi_1_49/Y sky130_fd_sc_hs__einvp_1_5/a_310_392#
+ sky130_fd_sc_hs__einvp_8_5/a_27_368# sky130_fd_sc_hs__inv_16_9/Y sky130_fd_sc_hs__nand2_4_45/Y
+ sky130_fd_sc_hs__a21oi_1_43/a_29_368# sky130_fd_sc_hs__nand2_2_77/Y sky130_fd_sc_hs__clkbuf_2_3/A
+ sky130_fd_sc_hs__nand2_4_9/a_27_74# sky130_fd_sc_hs__nand2_8_25/a_27_74# sky130_fd_sc_hs__inv_16_1/Y
+ sky130_fd_sc_hs__einvp_4_17/a_473_323# sky130_fd_sc_hs__nand2_2_53/a_27_74# sky130_fd_sc_hs__inv_16_13/Y
+ sky130_fd_sc_hs__nand2_4_47/a_27_74# sky130_fd_sc_hs__dlygate4sd3_1_78/a_289_74#
+ sky130_fd_sc_hs__inv_8_3/A sky130_fd_sc_hs__dlygate4sd3_1_14/a_289_74# sky130_fd_sc_hs__inv_8_9/A
+ sky130_fd_sc_hs__nand2_4_75/Y sky130_fd_sc_hs__nand2_4_61/a_27_74# sky130_fd_sc_hs__nand2_4_110/Y
+ sky130_fd_sc_hs__inv_4_9/Y sky130_fd_sc_hs__einvp_1_9/a_44_549# sky130_fd_sc_hs__inv_4_7/Y
+ sky130_fd_sc_hs__einvp_8_8/a_27_368# sky130_fd_sc_hs__inv_4_23/Y sky130_fd_sc_hs__dlygate4sd3_1_78/a_405_138#
+ sky130_fd_sc_hs__dlygate4sd3_1_45/a_28_74# sky130_fd_sc_hs__nand2_2_77/a_27_74#
+ sky130_fd_sc_hs__nand2_2_23/Y sky130_fd_sc_hs__einvp_8_9/a_27_368# sky130_fd_sc_hs__clkbuf_4_3/X
+ sky130_fd_sc_hs__nand2_4_40/Y sky130_fd_sc_hs__a21oi_1_13/a_29_368# sky130_fd_sc_hs__nand2_1_3/B
+ sky130_fd_sc_hs__nand2_8_1/a_27_74# sky130_fd_sc_hs__dlygate4sd3_1_25/X sky130_fd_sc_hs__dlygate4sd3_1_71/X
+ sky130_fd_sc_hs__nand2_2_21/a_27_74# sky130_fd_sc_hs__inv_4_1/Y sky130_fd_sc_hs__nand2_4_87/a_27_74#
+ sky130_fd_sc_hs__nand2_4_139/Y sky130_fd_sc_hs__nand2_4_115/a_27_74# sky130_fd_sc_hs__dlygate4sd2_1_1/a_28_74#
+ sky130_fd_sc_hs__dlygate4sd3_1_17/a_289_74# sky130_fd_sc_hs__dlygate4sd3_1_5/a_405_138#
+ sky130_fd_sc_hs__dlygate4sd3_1_79/A sky130_fd_sc_hs__clkbuf_2_14/a_43_192# sky130_fd_sc_hs__dlygate4sd3_1_62/a_289_74#
+ sky130_fd_sc_hs__dlygate4sd3_1_35/X sky130_fd_sc_hs__nand2_2_53/Y sky130_fd_sc_hs__nand2_4_31/a_27_74#
+ sky130_fd_sc_hs__nand2_8_19/a_27_74# sky130_fd_sc_hs__einvp_8_14/a_27_368# sky130_fd_sc_hs__inv_4_25/Y
+ sky130_fd_sc_hs__inv_8_1/A sky130_fd_sc_hs__inv_4_15/Y sky130_fd_sc_hs__dlygate4sd3_1_15/a_28_74#
+ sky130_fd_sc_hs__nand2_2_47/a_27_74# sky130_fd_sc_hs__and2_2_3/X sky130_fd_sc_hs__nand2_2_15/Y
+ sky130_fd_sc_hs__dlygate4sd3_1_3/a_289_74# sky130_fd_sc_hs__dlygate4sd3_1_63/A sky130_fd_sc_hs__a21oi_1_17/a_29_368#
+ sky130_fd_sc_hs__nand2_8_33/a_27_74# sky130_fd_sc_hs__einvp_8_9/a_802_323# sky130_fd_sc_hs__inv_16_5/Y
+ sky130_fd_sc_hs__dlygate4sd3_1_65/X sky130_fd_sc_hs__nand2_2_85/Y sky130_fd_sc_hs__nand2_2_61/a_27_74#
+ sky130_fd_sc_hs__einvp_2_1/a_263_323# sky130_fd_sc_hs__nand2_4_155/a_27_74# sky130_fd_sc_hs__dlygate4sd3_1_57/X
+ sky130_fd_sc_hs__dlygate4sd3_1_21/a_405_138# sky130_fd_sc_hs__dlygate4sd3_1_59/a_405_138#
+ sky130_fd_sc_hs__a21oi_1_47/a_117_74# sky130_fd_sc_hs__nand2_4_13/Y sky130_fd_sc_hs__nand2_4_151/Y
+ sky130_fd_sc_hs__dlygate4sd3_1_39/a_28_74# sky130_fd_sc_hs__nand2_2_61/B sky130_fd_sc_hs__inv_4_11/Y
+ sky130_fd_sc_hs__nand2_2_102/a_27_74# sky130_fd_sc_hs__einvp_2_13/a_27_368# sky130_fd_sc_hs__einvp_8_15/a_802_323#
+ sky130_fd_sc_hs__dlygate4sd3_1_65/a_289_74# sky130_fd_sc_hs__nand2_4_71/a_27_74#
+ sky130_fd_sc_hs__einvp_8_19/a_27_368# sky130_fd_sc_hs__dlygate4sd3_1_53/a_28_74#
+ sky130_fd_sc_hs__nand2_2_88/a_27_74# sky130_fd_sc_hs__nand2_2_15/a_27_74# sky130_fd_sc_hs__nand2_2_5/a_27_74#
+ sky130_fd_sc_hs__and4_2_3/C sky130_fd_sc_hs__a21oi_1_45/Y sky130_fd_sc_hs__nand2_4_110/a_27_74#
+ sky130_fd_sc_hs__inv_16_7/Y sky130_fd_sc_hs__einvp_4_5/a_27_368# sky130_fd_sc_hs__nand2_2_99/B
+ sky130_fd_sc_hs__dlygate4sd3_1_49/a_405_138# sky130_fd_sc_hs__a21oi_1_33/a_29_368#
+ sky130_fd_sc_hs__clkbuf_2_1/A sky130_fd_sc_hs__nand2_2_5/B sky130_fd_sc_hs__nand2_2_31/a_27_74#
+ sky130_fd_sc_hs__nand2_4_25/a_27_74# sky130_fd_sc_hs__inv_4_36/Y sky130_fd_sc_hs__nand2_2_9/B
+ sky130_fd_sc_hs__inv_4_39/Y sky130_fd_sc_hs__nand2_2_9/Y sky130_fd_sc_hs__dlygate4sd3_1_78/a_28_74#
+ sky130_fd_sc_hs__dfrtp_4_3/a_313_74# sky130_fd_sc_hs__nand2_2_39/Y sky130_fd_sc_hs__and4_2_1/a_143_74#
+ sky130_fd_sc_hs__inv_8_7/A sky130_fd_sc_hs__nand2_8_27/a_27_74# sky130_fd_sc_hs__nand2_4_73/Y
+ sky130_fd_sc_hs__buf_4_1/a_86_260# sky130_fd_sc_hs__inv_4_33/Y sky130_fd_sc_hs__dfrtp_4_3/a_494_366#
+ sky130_fd_sc_hs__dlygate4sd3_1_23/a_28_74# sky130_fd_sc_hs__clkbuf_4_3/a_83_270#
+ sky130_fd_sc_hs__einvp_1_19/a_310_392# sky130_fd_sc_hs__dlygate4sd3_1_49/X sky130_fd_sc_hs__dlygate4sd3_1_39/a_405_138#
+ sky130_fd_sc_hs__clkbuf_2_9/a_43_192# sky130_fd_sc_hs__nand2_8_43/a_27_74# sky130_fd_sc_hs__nand2_4_35/Y
+ sky130_fd_sc_hs__einvp_4_9/a_27_368# sky130_fd_sc_hs__nand2_2_69/Y sky130_fd_sc_hs__a21oi_1_35/a_29_368#
+ sky130_fd_sc_hs__nand2_1_1/B sky130_fd_sc_hs__nand2_2_71/a_27_74# sky130_fd_sc_hs__inv_4_29/Y
+ sky130_fd_sc_hs__nand2_4_65/a_27_74# sky130_fd_sc_hs__nand2_2_43/B sky130_fd_sc_hs__dfrtp_4_1/a_1647_81#
+ sky130_fd_sc_hs__nand2_4_137/Y sky130_fd_sc_hs__dlygate4sd3_1_47/a_28_74# sky130_fd_sc_hs__and4_2_5/a_143_74#
+ sky130_fd_sc_hs__a21oi_1_32/a_117_74# sky130_fd_sc_hs__einvp_2_5/a_27_368# sky130_fd_sc_hs__dlygate4sd3_1_45/A
+ sky130_fd_sc_hs__nand2_2_97/B sky130_fd_sc_hs__inv_8_5/A sky130_fd_sc_hs__nand2_2_51/Y
+ sky130_fd_sc_hs__dfrtp_4_1/a_890_138# sky130_fd_sc_hs__dlygate4sd3_1_29/a_405_138#
+ sky130_fd_sc_hs__dlygate4sd3_1_69/a_405_138# sky130_fd_sc_hs__nand2_2_97/a_27_74#
+ sky130_fd_sc_hs__nand2_2_25/a_27_74# sky130_fd_sc_hs__nand2_2_99/Y sky130_fd_sc_hs__nand2_4_19/a_27_74#
+ sky130_fd_sc_hs__nand2_4_117/a_27_74# sky130_fd_sc_hs__inv_16_9/A sky130_fd_sc_hs__nand2_4_29/Y
+ sky130_fd_sc_hs__einvp_8_19/a_27_74# sky130_fd_sc_hs__nand2_2_85/B sky130_fd_sc_hs__einvp_2_19/a_263_323#
+ sky130_fd_sc_hs__dfrtp_4_3/D sky130_fd_sc_hs__nand2_2_83/Y sky130_fd_sc_hs__dlygate4sd3_1_17/a_28_74#
+ sky130_fd_sc_hs__einvp_4_7/a_473_323# sky130_fd_sc_hs__nand2_4_11/Y sky130_fd_sc_hs__dlygate4sd3_1_20/a_405_138#
+ sky130_fd_sc_hs__a21oi_1_37/a_117_74# sky130_fd_sc_hs__einvp_2_9/a_27_368# sky130_fd_sc_hs__nand2_8_37/a_27_74#
+ sky130_fd_sc_hs__dlygate4sd3_1_56/a_289_74# sky130_fd_sc_hs__inv_4_31/Y sky130_fd_sc_hs__inv_1_9/Y
+ sky130_fd_sc_hs__nand2_2_65/a_27_74# sky130_fd_sc_hs__inv_16_31/A sky130_fd_sc_hs__einvp_4_7/a_27_74#
+ sky130_fd_sc_hs__dlygate4sd3_1_9/A sky130_fd_sc_hs__and2_2_1/B sky130_fd_sc_hs__nand2_4_159/Y
+ sky130_fd_sc_hs__einvp_1_3/a_318_74# sky130_fd_sc_hs__nand2_2_71/B sky130_fd_sc_hs__inv_4_19/Y
+ sky130_fd_sc_hs__einvp_2_15/a_36_74# sky130_fd_sc_hs__nand2_2_108/Y sky130_fd_sc_hs__buf_4_1/X
+ sky130_fd_sc_hs__nand2_2_73/Y sky130_fd_sc_hs__einvp_1_3/a_310_392# sky130_fd_sc_hs__nand2_4_89/Y
+ sky130_fd_sc_hs__dlygate4sd3_1_47/a_405_138# sky130_fd_sc_hs__nand2_2_19/a_27_74#
+ sky130_fd_sc_hs__nand2_2_9/a_27_74# sky130_fd_sc_hs__nand2_2_57/B sky130_fd_sc_hs__einvp_4_15/a_473_323#
+ sky130_fd_sc_hs__nand2_2_37/Y sky130_fd_sc_hs__dlygate4sd3_1_59/a_289_74# sky130_fd_sc_hs__einvp_1_11/a_44_549#
+ sky130_fd_sc_hs__dlygate4sd3_1_71/a_28_74# sky130_fd_sc_hs__dlygate4sd3_1_25/a_289_74#
+ sky130_fd_sc_hs__clkbuf_2_9/A sky130_fd_sc_hs__nand2_4_99/a_27_74# sky130_fd_sc_hs__nand2_4_27/a_27_74#
+ sky130_fd_sc_hs__nand2_4_71/Y sky130_fd_sc_hs__dlygate4sd2_1_1/X sky130_fd_sc_hs__nand2_4_106/Y
+ sky130_fd_sc_hs__nand2_4_127/a_27_74# sky130_fd_sc_hs__a21oi_1_1/a_117_74# sky130_fd_sc_hs__and4_2_5/D
+ sky130_fd_sc_hs__nand2_4_5/a_27_74# sky130_fd_sc_hs__einvp_1_7/a_318_74# sky130_fd_sc_hs__einvp_8_9/a_27_74#
+ sky130_fd_sc_hs__conb_1_1/LO sky130_fd_sc_hs__nand2_2_67/Y sky130_fd_sc_hs__einvp_4_11/a_27_368#
+ sky130_fd_sc_hs__inv_4_37/Y sky130_fd_sc_hs__dlygate4sd3_1_25/a_28_74# sky130_fd_sc_hs__einvp_8_2/a_27_368#
+ sky130_fd_sc_hs__nand3_4_3/a_27_82# sky130_fd_sc_hs__dfrtp_4_3/a_2010_409# sky130_fd_sc_hs__einvp_1_15/a_44_549#
+ sky130_fd_sc_hs__dlygate4sd3_1_41/a_28_74# sky130_fd_sc_hs__nand2_2_73/a_27_74#
+ sky130_fd_sc_hs__a21oi_1_23/a_117_74# sky130_fd_sc_hs__dlygate4sd3_1_75/a_289_74#
+ sky130_fd_sc_hs__dlygate4sd3_1_3/a_405_138# sky130_fd_sc_hs__dlygate4sd3_1_78/X
+ sky130_fd_sc_hs__dlygate4sd3_1_41/a_289_74# sky130_fd_sc_hs__a21oi_1_5/a_117_74#
+ sky130_fd_sc_hs__dlygate4sd3_1_68/a_405_138# sky130_fd_sc_hs__dlygate4sd3_1_59/X
+ sky130_fd_sc_hs__nand2_2_13/Y sky130_fd_sc_hs__nand2_4_83/a_27_74# sky130_fd_sc_hs__inv_4_21/Y
+ sky130_fd_sc_hs__nand2_2_59/Y sky130_fd_sc_hs__einvp_4_15/a_27_368# sky130_fd_sc_hs__einvp_4_19/a_27_74#
+ sky130_fd_sc_hs__nand2_8_7/a_27_74# sky130_fd_sc_hs__a21oi_1_29/a_29_368# sky130_fd_sc_hs__dlygate4sd3_1_62/X
+ sky130_fd_sc_hs__nand2_2_99/a_27_74# sky130_fd_sc_hs__einvp_8_7/a_802_323# sky130_fd_sc_hs__a21oi_1_42/a_29_368#
+ sky130_fd_sc_hs__dlygate4sd3_1_1/a_28_74# sky130_fd_sc_hs__nand2_8_15/a_27_74# sky130_fd_sc_hs__dfrtp_4_1/a_37_78#
+ sky130_fd_sc_hs__einvp_2_9/a_263_323# sky130_fd_sc_hs__einvp_1_19/a_44_549# sky130_fd_sc_hs__nand2_2_88/B
+ sky130_fd_sc_hs__nand2_2_43/Y sky130_fd_sc_hs__nand3_4_3/a_456_82# sky130_fd_sc_hs__and4_2_5/a_56_74#
+ sky130_fd_sc_hs__nand2_4_57/Y sky130_fd_sc_hs__nand2_4_39/a_27_74# sky130_fd_sc_hs__inv_1_7/Y
+ sky130_fd_sc_hs__nand2_4_135/a_27_74# sky130_fd_sc_hs__dlygate4sd3_1_45/a_289_74#
+ sky130_fd_sc_hs__a21oi_1_9/a_117_74# sky130_fd_sc_hs__dlygate4sd3_1_21/a_28_74#
+ sky130_fd_sc_hs__dlygate4sd3_1_7/A sky130_fd_sc_hs__and2_2_1/A sky130_fd_sc_hs__dfrtp_4_1/a_2010_409#
+ sky130_fd_sc_hs__einvp_4_1/a_27_74# sky130_fd_sc_hs__nand2_4_51/a_27_74# sky130_fd_sc_hs__clkbuf_4_1/A
+ sky130_fd_sc_hs__nand2_4_151/a_27_74# sky130_fd_sc_hs__einvp_4_19/a_27_368# sky130_fd_sc_hs__dlygate4sd3_1_35/a_28_74#
+ sky130_fd_sc_hs__dlygate4sd3_1_53/X sky130_fd_sc_hs__nand2_4_87/Y sky130_fd_sc_hs__dlygate4sd3_1_7/X
+ sky130_fd_sc_hs__a21oi_1_45/a_29_368# sky130_fd_sc_hs__nand2_1_5/B sky130_fd_sc_hs__nand2_2_108/a_27_74#
+ sky130_fd_sc_hs__nand2_2_79/B sky130_fd_sc_hs__dlygate4sd3_1_1/A sky130_fd_sc_hs__nand2_2_35/Y
+ sky130_fd_sc_hs__nand2_2_85/a_27_74# sky130_fd_sc_hs__nand2_2_13/a_27_74# sky130_fd_sc_hs__einvp_4_13/a_473_323#
+ sky130_fd_sc_hs__nand2_4_77/a_27_74# sky130_fd_sc_hs__nand2_2_1/a_27_74# sky130_fd_sc_hs__nand2_4_106/a_27_74#
+ sky130_fd_sc_hs__dlygate4sd3_1_49/a_289_74# sky130_fd_sc_hs__nand2_4_102/Y sky130_fd_sc_hs__a21oi_1_43/a_117_74#
+ sky130_fd_sc_hs__bufbuf_8_1/X sky130_fd_sc_hs__nand2_4_21/a_27_74# sky130_fd_sc_hs__dfrtp_4_1/a_494_366#
+ sky130_fd_sc_hs__einvp_8_15/a_27_368# sky130_fd_sc_hs__einvp_1_17/a_310_392# sky130_fd_sc_hs__and2_2_3/a_31_74#
+ sky130_fd_sc_hs__dlygate4sd3_1_37/a_405_138# sky130_fd_sc_hs__nand2_2_65/Y sky130_fd_sc_hs__nand2_2_37/a_27_74#
+ sky130_fd_sc_hs__and4_2_1/a_221_74# sky130_fd_sc_hs__a21oi_1_49/a_29_368# sky130_fd_sc_hs__clkbuf_2_1/a_43_192#
+ sky130_fd_sc_hs__einvp_4_1/a_27_368# sky130_fd_sc_hs__dlygate4sd3_1_75/A sky130_fd_sc_hs__nand2_4_145/a_27_74#
+ sky130_fd_sc_hs__nand2_4_61/Y sky130_fd_sc_hs__dlygate4sd3_1_21/a_289_74# sky130_fd_sc_hs__dlygate4sd3_1_29/a_28_74#
+ sky130_fd_sc_hs__a21oi_1_13/a_117_74# sky130_fd_sc_hs__nand2_2_96/Y sky130_fd_sc_hs__dlygate4sd3_1_31/a_289_74#
+ sky130_fd_sc_hs__dlygate4sd3_1_27/a_405_138# sky130_fd_sc_hs__nand2_4_60/a_27_74#
+ sky130_fd_sc_hs__dlygate4sd3_1_37/A sky130_fd_sc_hs__nand2_8_49/a_27_74# sky130_fd_sc_hs__nand2_4_25/Y
+ sky130_fd_sc_hs__and4_2_5/a_221_74# sky130_fd_sc_hs__dlygate4sd3_1_7/a_289_74# sky130_fd_sc_hs__clkbuf_2_5/a_43_192#
+ sky130_fd_sc_hs__nand2_2_93/a_27_74# sky130_fd_sc_hs__nand2_4_85/a_27_74# sky130_fd_sc_hs__nand2_4_15/a_27_74#
+ sky130_fd_sc_hs__dlygate4sd3_1_68/A sky130_fd_sc_hs__einvp_4_5/a_473_323# sky130_fd_sc_hs__nand2_4_55/Y
+ sky130_fd_sc_hs__dlygate4sd3_1_17/a_405_138# sky130_fd_sc_hs__dlygate4sd3_1_57/a_405_138#
+ sky130_fd_sc_hs__inv_1_9/A sky130_fd_sc_hs__a21oi_1_17/a_117_74# sky130_fd_sc_hs__nand2_2_89/Y
+ sky130_fd_sc_hs__einvp_2_17/a_27_368# sky130_fd_sc_hs__dlygate4sd3_1_51/X sky130_fd_sc_hs__dlygate4sd3_1_69/a_289_74#
+ sky130_fd_sc_hs__einvp_8_8/a_802_323# sky130_fd_sc_hs__and4_2_3/A sky130_fd_sc_hs__einvp_8_14/a_27_74#
+ sky130_fd_sc_hs__dfrtp_4_3/a_699_463# sky130_fd_sc_hs__dlygate4sd3_1_35/a_289_74#
+ sky130_fd_sc_hs__dlygate4sd3_1_3/a_28_74# sky130_fd_sc_hs__einvp_2_1/a_27_368# sky130_fd_sc_hs__and4_2_5/C
+ sky130_fd_sc_hs__nand2_8_17/a_27_74# sky130_fd_sc_hs__dlygate4sd3_1_14/a_28_74#
+ sky130_fd_sc_hs__conb_1_1/a_21_290# sky130_fd_sc_hs__nand2_4_139/a_27_74# sky130_fd_sc_hs__inv_1_1/Y
+ sky130_fd_sc_hs__clkbuf_2_8/a_43_192# sky130_fd_sc_hs__einvp_1_1/a_310_392# sky130_fd_sc_hs__nand2_2_3/Y
+ sky130_fd_sc_hs__nand2_4_55/a_27_74# sky130_fd_sc_hs__nand2_2_33/Y sky130_fd_sc_hs__and4_2_3/a_143_74#
+ sky130_fd_sc_hs__and4_2_3/B sky130_fd_sc_hs__dlygate4sd3_1_39/a_289_74# sky130_fd_sc_hs__a21oi_1_33/a_117_74#
+ sky130_fd_sc_hs__buf_4_1/A sky130_fd_sc_hs__clkbuf_4_5/a_83_270# sky130_fd_sc_hs__nand2_2_63/Y
+ sky130_fd_sc_hs__clkbuf_4_3/A sky130_fd_sc_hs__a21oi_1_39/a_29_368# sky130_fd_sc_hs__nand2_4_131/Y
+ sky130_fd_sc_hs__nand2_4_95/a_27_74# sky130_fd_sc_hs__nand2_4_123/a_27_74# sky130_fd_sc_hs__clkbuf_4_5/X
+ sky130_fd_sc_hs__nand2_4_1/a_27_74# sky130_fd_sc_hs__clkbuf_1_1/A sky130_fd_sc_hs__einvp_1_13/a_318_74#
+ sky130_fd_sc_hs__einvp_8_5/a_27_74# sky130_fd_sc_hs__a21oi_1_35/a_117_74# sky130_fd_sc_hs__nand2_1_9/Y
+ sky130_fd_sc_hs__dlygate4sd3_1_53/a_289_74# sky130_fd_sc_hs__dlygate4sd3_1_25/a_405_138#
+ sky130_fd_sc_hs__nand2_2_55/a_27_74# sky130_fd_sc_hs__nand2_4_23/Y sky130_fd_sc_hs__dlygate4sd3_1_65/a_405_138#
+ sky130_fd_sc_hs__nand2_4_49/a_27_74# sky130_fd_sc_hs__nand2_4_147/a_27_74# sky130_fd_sc_hs__nand2_8_41/a_27_74#
+ sky130_fd_sc_hs__dlygate4sd3_1_3/A sky130_fd_sc_hs__and2_2_3/A sky130_fd_sc_hs__nand2_2_7/B
+ sky130_fd_sc_hs__nand2_2_19/Y sky130_fd_sc_hs__einvp_2_17/a_263_323# sky130_fd_sc_hs__einvp_8_5/a_802_323#
+ sky130_fd_sc_hs__a21oi_1_21/a_29_368# sky130_fd_sc_hs__nand2_2_79/a_27_74# sky130_fd_sc_hs__nand2_4_53/Y
+ sky130_fd_sc_hs__clkbuf_2_8/A sky130_fd_sc_hs__and4_2_3/D sky130_fd_sc_hs__a21oi_1_3/a_29_368#
+ sky130_fd_sc_hs__einvp_1_17/a_318_74# sky130_fd_sc_hs__dlygate4sd2_1_1/A sky130_fd_sc_hs__dlygate4sd3_1_56/a_405_138#
+ sky130_fd_sc_hs__clkbuf_1_1/a_27_74# sky130_fd_sc_hs__einvp_4_15/a_27_74# sky130_fd_sc_hs__nand2_8_3/a_27_74#
+ sky130_fd_sc_hs__dlygate4sd3_1_63/a_28_74# sky130_fd_sc_hs__nand2_2_96/a_27_74#
+ sky130_fd_sc_hs__nand2_4_89/a_27_74# sky130_fd_sc_hs__inv_4_13/Y sky130_fd_sc_hs__nand2_2_49/Y
+ sky130_fd_sc_hs__einvp_2_1/a_36_74# sky130_fd_sc_hs__nand2_8_11/a_27_74# sky130_fd_sc_hs__nand2_2_102/Y
+ sky130_fd_sc_hs__and2_2_3/B sky130_fd_sc_hs__dfrtp_4_3/a_124_78# sky130_fd_sc_hs__nand2_4_83/Y
+ sky130_fd_sc_hs__and4_2_1/a_56_74# sky130_fd_sc_hs__nand2_4_33/a_27_74# sky130_fd_sc_hs__dlygate4sd3_1_7/a_28_74#
+ sky130_fd_sc_hs__nand2_1_3/a_117_74# sky130_fd_sc_hs__a21oi_1_25/a_29_368# sky130_fd_sc_hs__nand2_2_31/Y
+ sky130_fd_sc_hs__dlygate4sd3_1_45/a_405_138# sky130_fd_sc_hs__nand2_2_49/a_27_74#
+ sky130_fd_sc_hs__a21oi_1_7/a_29_368# sky130_fd_sc_hs__nand2_2_78/Y sky130_fd_sc_hs__dlygate4sd2_1_1/a_288_74#
+ sky130_fd_sc_hs__dlygate4sd3_1_31/a_28_74# sky130_fd_sc_hs__dlygate4sd3_1_29/a_289_74#
+ sky130_fd_sc_hs__clkbuf_2_7/X sky130_fd_sc_hs__dlygate4sd3_1_74/a_289_74# sky130_fd_sc_hs__nand2_4_157/a_27_74#
+ sky130_fd_sc_hs__dlygate4sd3_1_43/X sky130_fd_sc_hs__nand2_4_111/Y sky130_fd_sc_hs__einvp_1_15/a_310_392#
+ sky130_fd_sc_hs__nand2_4_73/a_27_74# sky130_fd_sc_hs__dlygate4sd3_1_35/a_405_138#
+ sky130_fd_sc_hs__dlygate4sd3_1_75/a_405_138# sky130_fd_sc_hs__einvp_1_3/a_44_549#
+ sky130_fd_sc_hs__einvp_4_13/a_27_368# sky130_fd_sc_hs__nand2_1_7/a_117_74# sky130_fd_sc_hs__a21oi_1_28/a_29_368#
+ sky130_fd_sc_hs__dlygate4sd3_1_57/a_28_74# sky130_fd_sc_hs__nand2_4_9/Y sky130_fd_sc_hs__nand2_2_7/a_27_74#
+ sky130_fd_sc_hs__dfrtp_4_3/a_1827_81# sky130_fd_sc_hs__nand2_2_92/Y sky130_fd_sc_hs__nand2_1_7/Y
+ sky130_fd_sc_hs__nand2_2_33/a_27_74# sky130_fd_sc_hs__dlygate4sd3_1_33/A sky130_fd_sc_hs__nand2_2_65/B
+ sky130_fd_sc_hs__nand2_4_21/Y sky130_fd_sc_hs__dlygate4sd3_1_1/a_405_138# sky130_fd_sc_hs__dlygate4sd3_1_11/a_289_74#
+ sky130_fd_sc_hs__nand2_4_69/Y sky130_fd_sc_hs__and2_2_3/a_118_74# sky130_fd_sc_hs__and4_2_1/X
+ sky130_fd_sc_hs__nand2_4_41/a_27_74# sky130_fd_sc_hs__einvp_1_7/a_44_549# sky130_fd_sc_hs__nand2_4_141/a_27_74#
+ sky130_fd_sc_hs__nand2_4_121/Y sky130_fd_sc_hs__nand2_2_17/Y sky130_fd_sc_hs__einvp_8_7/a_27_368#
+ sky130_fd_sc_hs__einvp_2_15/a_263_323# sky130_fd_sc_hs__a21oi_1_11/a_29_368# sky130_fd_sc_hs__nand2_8_45/a_27_74#
+ sky130_fd_sc_hs__einvp_2_7/a_263_323# sky130_fd_sc_hs__nand2_4_99/Y sky130_fd_sc_hs__nand2_4_67/a_27_74#
+ sky130_fd_sc_hs__a21oi_1_29/a_117_74# sky130_fd_sc_hs__dlygate4sd3_1_3/X sky130_fd_sc_hs__dlygate4sd3_1_53/a_405_138#
+ sky130_fd_sc_hs__dlygate4sd3_1_47/a_289_74# sky130_fd_sc_hs__nand2_2_73/B sky130_fd_sc_hs__dfrtp_4_1/a_699_463#
+ sky130_fd_sc_hs__a21oi_1_42/a_117_74# sky130_fd_sc_hs__nand2_2_47/Y sky130_fd_sc_hs__nand2_4_11/a_27_74#
+ sky130_fd_sc_hs__nand2_4_81/Y sky130_fd_sc_hs__nand2_4_115/Y sky130_fd_sc_hs__dlygate4sd3_1_65/a_28_74#
+ sky130_fd_sc_hs__nand2_2_27/a_27_74# sky130_fd_sc_hs__einvp_8_8/a_27_74# sky130_fd_sc_hs__nand2_4_119/a_27_74#
+ sky130_fd_sc_hs__nand2_4_43/Y sky130_fd_sc_hs__einvp_2_3/a_36_74# sky130_fd_sc_hs__a21oi_1_15/a_29_368#
+ sky130_fd_sc_hs__nand2_8_13/a_27_74# sky130_fd_sc_hs__and4_2_3/a_56_74# sky130_fd_sc_hs__nand2_2_43/a_27_74#
+ sky130_fd_sc_hs__dlygate4sd3_1_20/A sky130_fd_sc_hs__nand2_4_35/a_27_74# sky130_fd_sc_hs__nand2_2_37/B
+ sky130_fd_sc_hs__einvp_4_11/a_473_323# sky130_fd_sc_hs__dlygate4sd3_1_9/X sky130_fd_sc_hs__and4_2_5/B
+ sky130_fd_sc_hs__nand2_4_145/Y sky130_fd_sc_hs__dlygate4sd3_1_20/a_289_74# sky130_fd_sc_hs__a21oi_1_45/a_117_74#
+ sky130_fd_sc_hs__dlygate4sd3_1_20/a_28_74# sky130_fd_sc_hs__clkbuf_2_17/a_43_192#
+ sky130_fd_sc_hs__nand3_4_3/C sky130_fd_sc_hs__dfrtp_4_3/a_789_463# sky130_fd_sc_hs__einvp_8_17/a_27_368#
+ sky130_fd_sc_hs__nand2_8_39/a_27_74# sky130_fd_sc_hs__bufbuf_8_1/a_221_368# sky130_fd_sc_hs__and4_2_3/a_221_74#
+ sky130_fd_sc_hs__nand2_2_67/a_27_74# sky130_fd_sc_hs__einvp_4_9/a_27_74# sky130_fd_sc_hs__dlygate4sd3_1_74/a_405_138#
+ sky130_fd_sc_hs__nand2_2_21/Y sky130_fd_sc_hs__nand2_4_159/a_27_74# sky130_fd_sc_hs__dlygate4sd3_1_5/a_289_74#
+ sky130_fd_sc_hs__nand2_4_39/Y sky130_fd_sc_hs__nand2_4_7/Y sky130_fd_sc_hs__a21oi_1_19/a_29_368#
+ sky130_fd_sc_hs__nand2_2_105/a_27_74# sky130_fd_sc_hs__nand2_2_12/a_27_74# sky130_fd_sc_hs__nand2_2_84/a_27_74#
+ sky130_fd_sc_hs__nand2_1_5/Y sky130_fd_sc_hs__nand2_4_103/a_27_74# sky130_fd_sc_hs__a21oi_1_49/a_117_74#
+ sky130_fd_sc_hs__dlygate4sd3_1_59/a_28_74# sky130_fd_sc_hs__einvp_2_15/a_27_368#
+ sky130_fd_sc_hs__dfrtp_4_1/a_313_74# sky130_fd_sc_hs__dlygate4sd3_1_68/a_289_74#
+ sky130_fd_sc_hs__dlygate4sd3_1_79/X sky130_fd_sc_hs__inv_1_7/A sky130_fd_sc_hs__nand2_4_91/a_27_74#
+ sky130_fd_sc_hs__nand2_4_67/Y sky130_fd_sc_hs__inv_4_27/Y sky130_fd_sc_hs__dlygate4sd3_1_75/a_28_74#
+ sky130_fd_sc_hs__clkbuf_4_1/a_83_270# sky130_fd_sc_hs__einvp_8_3/a_27_74# sky130_fd_sc_hs__nand2_4_129/a_27_74#
+ sky130_fd_sc_hs__nand2_8_23/a_27_74# sky130_fd_sc_hs__nand2_4_7/a_27_74# sky130_fd_sc_hs__einvp_4_7/a_27_368#
+ sky130_fd_sc_hs__nand2_2_51/a_27_74# sky130_fd_sc_hs__dfrtp_4_3/a_834_355# sky130_fd_sc_hs__nand2_4_45/a_27_74#
+ sky130_fd_sc_hs__nand2_2_84/Y sky130_fd_sc_hs__nand2_4_97/Y sky130_fd_sc_hs__einvp_2_5/a_263_323#
+ sky130_fd_sc_hs__einvp_4_3/a_473_323# sky130_fd_sc_hs__dlygate4sd3_1_15/a_405_138#
+ sky130_fd_sc_hs__dfrtp_4_3/a_1627_493# sky130_fd_sc_hs__einvp_2_19/a_27_368# sky130_fd_sc_hs__einvp_8_19/a_802_323#
+ sky130_fd_sc_hs__nand2_2_45/Y sky130_fd_sc_hs__einvp_2_3/a_27_368# sky130_fd_sc_hs__dfrtp_4_3/a_812_138#
+ sky130_fd_sc_hs__dlygate4sd3_1_43/a_28_74# sky130_fd_sc_hs__nand2_4_113/Y sky130_fd_sc_hs__dlygate4sd3_1_53/A
+ sky130_fd_sc_hs__einvp_4_11/a_27_74# sky130_fd_sc_hs__nand2_4_41/Y sky130_fd_sc_hs__nand2_2_92/a_27_74#
+ sky130_fd_sc_hs__nand2_2_109/Y sky130_fd_sc_hs__einvp_1_9/a_310_392# sky130_fd_sc_hs__dlygate4sd3_1_43/a_405_138#
+ sky130_fd_sc_hs__nand2_4_113/a_27_74# sky130_fd_sc_hs__clkbuf_2_1/X sky130_fd_sc_hs__nand2_8_9/a_27_74#
+ sky130_fd_sc_hs__nand2_2_35/B sky130_fd_sc_hs__dlygate4sd3_1_69/a_28_74# sky130_fd_sc_hs__nand2_2_7/Y
+ sky130_fd_sc_hs__nand2_4_143/Y sky130_fd_sc_hs__einvp_8_15/a_27_74# sky130_fd_sc_hs__einvp_2_7/a_36_74#
+ sky130_fd_sc_hs__dfrtp_4_3/a_37_78# sky130_fd_sc_hs__nand2_4_107/Y sky130_fd_sc_hs__nand2_2_45/a_27_74#
+ sky130_fd_sc_hs__einvp_1_13/a_310_392# sky130_fd_sc_hs__dfrtp_4_1/a_1627_493# sky130_fd_sc_hs__einvp_1_1/a_318_74#
+ sky130_fd_sc_hs__dlygate4sd3_1_33/a_405_138# sky130_fd_sc_hs__nand2_4_5/Y sky130_fd_sc_hs__dlygate4sd3_1_71/a_405_138#
+ sky130_fd_sc_hs__einvp_4_3/a_27_74# sky130_fd_sc_hs__nand2_4_153/a_27_74# sky130_fd_sc_hs__dlygate4sd3_1_37/a_28_74#
+ sky130_fd_sc_hs__nand2_1_3/Y sky130_fd_sc_hs__nand2_4_135/Y sky130_fd_sc_hs__dfrtp_4_1/a_1827_81#
+ sky130_fd_sc_hs__a21oi_1_39/a_117_74# sky130_fd_sc_hs__einvp_2_11/a_36_74# sky130_fd_sc_hs__inv_1_5/A
+ sky130_fd_sc_hs__dlygate4sd3_1_51/a_28_74# sky130_fd_sc_hs__nand2_4_65/Y sky130_fd_sc_hs__nand2_4_79/a_27_74#
+ sky130_fd_sc_hs__dlygate4sd3_1_23/a_405_138# sky130_fd_sc_hs__dlygate4sd3_1_63/a_405_138#
+ sky130_fd_sc_hs__einvp_1_5/a_318_74# sky130_fd_sc_hs__nand2_4_27/Y sky130_fd_sc_hs__nand2_4_23/a_27_74#
+ sky130_fd_sc_hs__nand2_4_121/a_27_74# sky130_fd_sc_hs__einvp_2_13/a_263_323# sky130_fd_sc_hs__nand2_4_129/Y
+ sky130_fd_sc_hs__nand2_2_39/a_27_74# sky130_fd_sc_hs__nand2_4_95/Y sky130_fd_sc_hs__clkbuf_2_17/A
+ sky130_fd_sc_hs__dlygate4sd3_1_14/a_405_138# sky130_fd_sc_hs__dlygate4sd3_1_51/a_405_138#
+ sky130_fd_sc_hs__einvp_1_13/a_44_549# sky130_fd_sc_hs__a21oi_1_21/a_117_74# sky130_fd_sc_hs__dlygate4sd3_1_71/a_289_74#
+ sky130_fd_sc_hs__a21oi_1_3/a_117_74# sky130_fd_sc_hs__einvp_1_9/a_318_74# sky130_fd_sc_hs__conb_1_1/a_165_290#
+ sky130_fd_sc_hs__nand2_4_63/a_27_74# sky130_fd_sc_hs__nand2_2_105/Y sky130_fd_sc_hs__and4_2_1/a_335_74#
+ sky130_fd_sc_hs__nand2_2_78/a_27_74# sky130_fd_sc_hs__nand2_2_5/Y sky130_fd_sc_hs__nand2_4_141/Y
+ sky130_fd_sc_hs__dfrtp_4_3/a_1678_395# sky130_fd_sc_hs__einvp_1_17/a_44_549# sky130_fd_sc_hs__einvp_4_13/a_27_74#
+ sky130_fd_sc_hs__dlygate4sd3_1_62/a_28_74# sky130_fd_sc_hs__nand2_2_23/a_27_74#
+ sky130_fd_sc_hs__nand3_4_1/a_456_82# sky130_fd_sc_hs__a21oi_1_25/a_117_74# sky130_fd_sc_hs__nand2_4_17/a_27_74#
+ sky130_fd_sc_hs__nand2_4_103/Y sky130_fd_sc_hs__dlygate4sd3_1_43/a_289_74# sky130_fd_sc_hs__dfrtp_4_1/a_789_463#
+ sky130_fd_sc_hs__a21oi_1_7/a_117_74# sky130_fd_sc_hs__einvp_8_17/a_27_74# sky130_fd_sc_hs__dlygate4sd3_1_5/a_28_74#
+ sky130_fd_sc_hs__nand2_4_3/Y sky130_fd_sc_hs__nand2_4_33/Y sky130_fd_sc_hs__einvp_2_9/a_36_74#
+ sky130_fd_sc_hs__einvp_4_17/a_27_368# sky130_fd_sc_hs__nand2_4_131/a_27_74# sky130_fd_sc_hs__and4_2_5/a_335_74#
+ sky130_fd_sc_hs__nand2_1_1/Y sky130_fd_sc_hs__clkbuf_4_5/A sky130_fd_sc_hs__nand2_4_133/Y
+ sky130_fd_sc_hs__nand2_8_35/a_27_74# sky130_fd_sc_hs__nand2_2_29/Y sky130_fd_sc_hs__dlygate4sd2_1_1/a_405_138#
+ sky130_fd_sc_hs__nand2_2_63/a_27_74# sky130_fd_sc_hs__a21oi_1_28/a_117_74# sky130_fd_sc_hs__einvp_4_5/a_27_74#
+ sky130_fd_sc_hs__nand2_4_57/a_27_74# sky130_fd_sc_hs__dlygate4sd3_1_79/a_289_74#
+ sky130_fd_sc_hs__nand2_4_63/Y sky130_fd_sc_hs__dlygate4sd3_1_9/a_405_138# sky130_fd_sc_hs__dlygate4sd3_1_15/a_289_74#
+ sky130_fd_sc_hs__nand2_2_97/Y sky130_fd_sc_hs__nand2_2_103/a_27_74# sky130_fd_sc_hs__dlygate4sd3_1_62/a_405_138#
+ sky130_fd_sc_hs__nand2_2_12/Y sky130_fd_sc_hs__einvp_2_13/a_36_74# sky130_fd_sc_hs__dfrtp_4_1/a_1678_395#
+ sky130_fd_sc_hs__dlygate4sd3_1_56/a_28_74# sky130_fd_sc_hs__bufbuf_8_1/a_334_368#
+ sky130_fd_sc_hs__nand2_2_17/a_27_74# sky130_fd_sc_hs__nand2_2_89/a_27_74# sky130_fd_sc_hs__nand2_4_111/a_27_74#
+ sky130_fd_sc_hs__a21oi_1_47/a_29_368# sky130_fd_sc_hs__nand2_4_127/Y sky130_fd_sc_hs__dlygate4sd3_1_1/a_289_74#
+ sky130_fd_sc_hs__nand2_4_93/Y sky130_fd_sc_hs__einvp_8_3/a_802_323# sky130_fd_sc_hs__dfrtp_4_1/a_834_355#
+ sky130_fd_sc_hs__einvp_2_3/a_263_323# sky130_fd_sc_hs__einvp_4_1/a_473_323# sky130_fd_sc_hs__nand2_4_97/a_27_74#
+ sky130_fd_sc_hs__nand2_2_42/Y sky130_fd_sc_hs__nand2_4_125/a_27_74# sky130_fd_sc_hs__nand2_4_3/a_27_74#
+ sky130_fd_sc_hs__dlygate4sd3_1_79/a_28_74# sky130_fd_sc_hs__einvp_8_17/a_802_323#
+ sky130_fd_sc_hs__a21oi_1_11/a_117_74# sky130_fd_sc_hs__and4_2_5/A sky130_fd_sc_hs__einvp_2_11/a_27_368#
+ sky130_fd_sc_hs__clkbuf_2_15/a_43_192# sky130_fd_sc_hs__dlygate4sd3_1_63/a_289_74#
+ sky130_fd_sc_hs__dfrtp_4_1/a_812_138# sky130_fd_sc_hs__einvp_8_7/a_27_74# sky130_fd_sc_hs__nand2_4_157/Y
+ sky130_fd_sc_hs__nand2_4_19/Y sky130_fd_sc_hs__nand2_8_29/a_27_74# sky130_fd_sc_hs__nand2_2_57/a_27_74#
+ sky130_fd_sc_hs__nand3_4_1/a_27_82# sky130_fd_sc_hs__nand2_2_71/Y sky130_fd_sc_hs__nand2_4_149/a_27_74#
+ sky130_fd_sc_hs__nand2_4_119/Y sky130_fd_sc_hs__nand2_4_85/Y sky130_fd_sc_hs__clkbuf_2_3/a_43_192#
+ sky130_fd_sc_hs__einvp_1_7/a_310_392# sky130_fd_sc_hs__einvp_4_3/a_27_368# sky130_fd_sc_hs__dlygate4sd3_1_41/a_405_138#
+ sky130_fd_sc_hs__dfrtp_4_3/a_1350_392# sky130_fd_sc_hs__nand2_4_49/Y sky130_fd_sc_hs__einvp_4_19/a_473_323#
+ sky130_fd_sc_hs__dlygate4sd3_1_49/a_28_74# sky130_fd_sc_hs__a21oi_1_15/a_117_74#
+ sky130_fd_sc_hs__dlygate4sd3_1_33/a_289_74# sky130_fd_sc_hs__nand2_4_81/a_27_74#
+ sky130_fd_sc_hs__nand2_4_149/Y sky130_fd_sc_hs__einvp_4_17/a_27_74# sky130_fd_sc_hs__nand2_8_5/a_27_74#
+ sky130_fd_sc_hs__nand2_4_1/Y sky130_fd_sc_hs__nand2_4_31/Y sky130_fd_sc_hs__einvp_1_11/a_310_392#
+ sky130_fd_sc_hs__dlygate4sd3_1_31/a_405_138# sky130_fd_sc_hs__nand2_4_79/Y sky130_fd_sc_hs__dlygate4sd3_1_9/a_289_74#
+ sky130_fd_sc_hs__clkbuf_2_7/a_43_192# sky130_fd_sc_hs__a21oi_1_32/a_29_368# sky130_fd_sc_hs__nand2_2_42/a_27_74#
+ sky130_fd_sc_hs__dlygate4sd3_1_9/a_28_74# sky130_fd_sc_hs__nand2_2_27/Y sky130_fd_sc_hs__nand2_4_133/a_27_74#
+ sky130_fd_sc_hs__nand2_1_7/B sky130_fd_sc_hs__nand2_4_60/Y sky130_fd_sc_hs__a21oi_1_19/a_117_74#
+ sky130_fd_sc_hs__dlygate4sd3_1_37/a_289_74# sky130_fd_sc_hs__dfrtp_4_1/a_1350_392#
+ sky130_fd_sc_hs__dlygate4sd3_1_33/a_28_74# sky130_fd_sc_hs__nand2_2_57/Y sky130_fd_sc_hs__nand2_4_125/Y
+ sky130_fd_sc_hs__nand2_4_91/Y sky130_fd_sc_hs__a21oi_1_37/a_29_368# sky130_fd_sc_hs__nand2_2_83/a_27_74#
+ sky130_fd_sc_hs__nand2_4_75/a_27_74# sky130_fd_sc_hs__einvp_8_2/a_802_323# sky130_fd_sc_hs__einvp_2_17/a_36_74#
+ sky130_fd_sc_hs__nand2_4_102/a_27_74# sky130_fd_sc_hs__dlygate4sd3_1_11/a_405_138#
+ sky130_fd_sc_hs__einvp_1_11/a_318_74# sky130_fd_sc_hs__nand2_2_88/Y sky130_fd_sc_hs__einvp_2_7/a_27_368#
+ sky130_fd_sc_hs__and2_2_1/a_31_74# sky130_fd_sc_hs__dlygate4sd3_1_51/a_289_74# sky130_fd_sc_hs__nand2_4_17/Y
+ sky130_fd_sc_hs__dlygate4sd3_1_74/a_28_74# sky130_fd_sc_hs__nand2_4_155/Y sky130_fd_sc_hs__nand2_2_35/a_27_74#
+ sky130_fd_sc_hs__nand2_4_29/a_27_74# sky130_fd_sc_hs__einvp_8_2/a_27_74# sky130_fd_sc_hs__nand2_2_103/Y
+ sky130_fd_sc_hs__nand2_8_21/a_27_74# sky130_fd_sc_hs__nand2_4_117/Y sky130_fd_sc_hs__nand2_2_1/Y
+ sky130_fd_sc_hs__nand2_4_43/a_27_74# sky130_fd_sc_hs__nand2_4_143/a_27_74# sky130_fd_sc_hs__dlygate4sd3_1_27/a_28_74#
+ sky130_fd_sc_hs__nand2_4_47/Y sky130_fd_sc_hs__nand2_2_59/a_27_74# sky130_fd_sc_hs__einvp_1_15/a_318_74#
+ sky130_fd_sc_hs__a21oi_1_1/a_29_368# sky130_fd_sc_hs__nand2_2_79/Y sky130_fd_sc_hs__nand2_8_47/a_27_74#
+ sky130_fd_sc_hs__dlygate4sd3_1_57/a_289_74# sky130_fd_sc_hs__bufbuf_8_1/a_27_112#
+ sky130_fd_sc_hs__nand2_4_147/Y sky130_fd_sc_hs__dlygate4sd3_1_23/a_289_74# sky130_fd_sc_hs__nand2_4_69/a_27_74#
+ sky130_fd_sc_hs__nand2_2_61/Y sky130_fd_sc_hs__nand2_4_77/Y sky130_fd_sc_hs__dfrtp_4_1/a_124_78#
+ sky130_fd_sc_hs__dlygate4sd3_1_79/a_405_138# sky130_fd_sc_hs__nand2_4_13/a_27_74#
+ sky130_fd_sc_hs__nand2_2_25/Y sky130_fd_sc_hs__nand2_1_1/a_117_74# sky130_fd_sc_hs__dlygate4sd3_1_68/a_28_74#
+ sky130_fd_sc_hs__a21oi_1_23/a_29_368# sky130_fd_sc_hs__nand2_2_29/a_27_74# sky130_fd_sc_hs__einvp_1_19/a_318_74#
+ sky130_fd_sc_hs__a21oi_1_5/a_29_368# sky130_fd_sc_hs__dfrtp_4_3/a_1647_81#
Xsky130_fd_sc_hs__nand2_4_13 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_4_13/Y delay_con_msb[2]
+ osc_144 sky130_fd_sc_hs__nand2_4_13/a_27_74# sky130_fd_sc_hs__nand2_4
Xsky130_fd_sc_hs__nand2_4_24 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_4_25/Y delay_con_msb[1]
+ osc_000 sky130_fd_sc_hs__nand2_4_25/a_27_74# sky130_fd_sc_hs__nand2_4
Xsky130_fd_sc_hs__nand2_4_35 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_4_35/Y delay_con_msb[2]
+ osc_144 sky130_fd_sc_hs__nand2_4_35/a_27_74# sky130_fd_sc_hs__nand2_4
Xsky130_fd_sc_hs__nand2_4_46 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_4_47/Y delay_con_msb[0]
+ osc_144 sky130_fd_sc_hs__nand2_4_47/a_27_74# sky130_fd_sc_hs__nand2_4
Xsky130_fd_sc_hs__nand2_4_57 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_4_57/Y delay_con_msb[0]
+ osc_000 sky130_fd_sc_hs__nand2_4_57/a_27_74# sky130_fd_sc_hs__nand2_4
Xsky130_fd_sc_hs__nand2_4_68 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_4_69/Y delay_con_msb[0]
+ osc_144 sky130_fd_sc_hs__nand2_4_69/a_27_74# sky130_fd_sc_hs__nand2_4
Xsky130_fd_sc_hs__nand2_4_79 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_4_79/Y delay_con_msb[1]
+ osc_108 sky130_fd_sc_hs__nand2_4_79/a_27_74# sky130_fd_sc_hs__nand2_4
Xsky130_fd_sc_hs__einvp_4_3 DVSS DVDD DVDD DVSS pi3_r[2] sky130_fd_sc_hs__inv_8_1/A
+ sky130_fd_sc_hs__inv_4_5/Y sky130_fd_sc_hs__einvp_4_3/a_27_74# sky130_fd_sc_hs__einvp_4_3/a_27_368#
+ sky130_fd_sc_hs__einvp_4_3/a_473_323# sky130_fd_sc_hs__einvp_4
Xsky130_fd_sc_hs__and2_2_0 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__and2_2_1/A sky130_fd_sc_hs__and2_2_1/B
+ inj_out sky130_fd_sc_hs__and2_2_1/a_31_74# sky130_fd_sc_hs__and2_2_1/a_118_74# sky130_fd_sc_hs__and2_2
Xsky130_fd_sc_hs__inv_4_8 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_9/Y osc_000 sky130_fd_sc_hs__inv_4
Xsky130_fd_sc_hs__einvp_2_0 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_8_1/A sky130_fd_sc_hs__inv_4_3/Y
+ pi3_l[1] sky130_fd_sc_hs__einvp_2_1/a_263_323# sky130_fd_sc_hs__einvp_2_1/a_36_74#
+ sky130_fd_sc_hs__einvp_2_1/a_27_368# sky130_fd_sc_hs__einvp_2
Xsky130_fd_sc_hs__clkbuf_2_14 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__clkbuf_2_8/A sky130_fd_sc_hs__clkbuf_4_5/X
+ sky130_fd_sc_hs__clkbuf_2_14/a_43_192# sky130_fd_sc_hs__clkbuf_2
Xsky130_fd_sc_hs__clkbuf_2_3 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__clkbuf_4_3/A sky130_fd_sc_hs__clkbuf_2_3/A
+ sky130_fd_sc_hs__clkbuf_2_3/a_43_192# sky130_fd_sc_hs__clkbuf_2
Xsky130_fd_sc_hs__einvp_4_18 DVSS DVDD DVDD DVSS pi5_r[2] sky130_fd_sc_hs__inv_8_9/A
+ sky130_fd_sc_hs__inv_4_21/Y sky130_fd_sc_hs__einvp_4_19/a_27_74# sky130_fd_sc_hs__einvp_4_19/a_27_368#
+ sky130_fd_sc_hs__einvp_4_19/a_473_323# sky130_fd_sc_hs__einvp_4
Xsky130_fd_sc_hs__dlygate4sd3_1_15 DVSS DVDD DVSS DVDD sky130_fd_sc_hs__dlygate4sd3_1_7/X
+ sky130_fd_sc_hs__dlygate4sd3_1_20/A sky130_fd_sc_hs__dlygate4sd3_1_15/a_405_138#
+ sky130_fd_sc_hs__dlygate4sd3_1_15/a_28_74# sky130_fd_sc_hs__dlygate4sd3_1_15/a_289_74#
+ sky130_fd_sc_hs__dlygate4sd3_1
Xsky130_fd_sc_hs__dlygate4sd3_1_37 DVSS DVDD DVSS DVDD sky130_fd_sc_hs__dlygate4sd3_1_37/A
+ sky130_fd_sc_hs__dlygate4sd3_1_56/A sky130_fd_sc_hs__dlygate4sd3_1_37/a_405_138#
+ sky130_fd_sc_hs__dlygate4sd3_1_37/a_28_74# sky130_fd_sc_hs__dlygate4sd3_1_37/a_289_74#
+ sky130_fd_sc_hs__dlygate4sd3_1
Xsky130_fd_sc_hs__dlygate4sd3_1_48 DVSS DVDD DVSS DVDD sky130_fd_sc_hs__dlygate4sd3_1_51/X
+ sky130_fd_sc_hs__dlygate4sd3_1_49/X sky130_fd_sc_hs__dlygate4sd3_1_49/a_405_138#
+ sky130_fd_sc_hs__dlygate4sd3_1_49/a_28_74# sky130_fd_sc_hs__dlygate4sd3_1_49/a_289_74#
+ sky130_fd_sc_hs__dlygate4sd3_1
Xsky130_fd_sc_hs__dlygate4sd3_1_59 DVSS DVDD DVSS DVDD sky130_fd_sc_hs__dlygate4sd3_1_65/X
+ sky130_fd_sc_hs__dlygate4sd3_1_59/X sky130_fd_sc_hs__dlygate4sd3_1_59/a_405_138#
+ sky130_fd_sc_hs__dlygate4sd3_1_59/a_28_74# sky130_fd_sc_hs__dlygate4sd3_1_59/a_289_74#
+ sky130_fd_sc_hs__dlygate4sd3_1
Xsky130_fd_sc_hs__dlygate4sd3_1_26 DVSS DVDD DVSS DVDD sky130_fd_sc_hs__dlygate4sd3_1_31/X
+ sky130_fd_sc_hs__dlygate4sd3_1_33/A sky130_fd_sc_hs__dlygate4sd3_1_27/a_405_138#
+ sky130_fd_sc_hs__dlygate4sd3_1_27/a_28_74# sky130_fd_sc_hs__dlygate4sd3_1_27/a_289_74#
+ sky130_fd_sc_hs__dlygate4sd3_1
Xsky130_fd_sc_hs__nand2_4_9 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_4_9/Y delay_con_msb[2]
+ osc_144 sky130_fd_sc_hs__nand2_4_9/a_27_74# sky130_fd_sc_hs__nand2_4
Xsky130_fd_sc_hs__nand2_2_90 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_2_92/Y sky130_fd_sc_hs__nand2_2_97/B
+ osc_036 sky130_fd_sc_hs__nand2_2_92/a_27_74# sky130_fd_sc_hs__nand2_2
Xsky130_fd_sc_hs__nand2_2_108 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_2_108/Y sky130_fd_sc_hs__a21oi_1_49/Y
+ osc_036 sky130_fd_sc_hs__nand2_2_108/a_27_74# sky130_fd_sc_hs__nand2_2
Xsky130_fd_sc_hs__inv_16_15 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__and4_2_5/A sky130_fd_sc_hs__inv_16_7/Y
+ sky130_fd_sc_hs__inv_16
Xsky130_fd_sc_hs__inv_16_26 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_16_31/A sky130_fd_sc_hs__inv_4_27/Y
+ sky130_fd_sc_hs__inv_16
Xsky130_fd_sc_hs__nand2_2_6 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_2_7/Y sky130_fd_sc_hs__nand2_2_7/B
+ osc_144 sky130_fd_sc_hs__nand2_2_7/a_27_74# sky130_fd_sc_hs__nand2_2
Xsky130_fd_sc_hs__einvp_1_19 DVSS DVDD DVDD DVSS pi5_r[0] sky130_fd_sc_hs__inv_8_9/A
+ sky130_fd_sc_hs__inv_4_21/Y sky130_fd_sc_hs__einvp_1_19/a_44_549# sky130_fd_sc_hs__einvp_1_19/a_318_74#
+ sky130_fd_sc_hs__einvp_1_19/a_310_392# sky130_fd_sc_hs__einvp_1
Xsky130_fd_sc_hs__nand2_4_14 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_4_15/Y delay_con_msb[1]
+ osc_000 sky130_fd_sc_hs__nand2_4_15/a_27_74# sky130_fd_sc_hs__nand2_4
Xsky130_fd_sc_hs__nand2_4_25 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_4_25/Y delay_con_msb[1]
+ osc_000 sky130_fd_sc_hs__nand2_4_25/a_27_74# sky130_fd_sc_hs__nand2_4
Xsky130_fd_sc_hs__nand2_4_36 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_4_39/Y delay_con_msb[2]
+ osc_000 sky130_fd_sc_hs__nand2_4_39/a_27_74# sky130_fd_sc_hs__nand2_4
Xsky130_fd_sc_hs__nand2_4_47 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_4_47/Y delay_con_msb[0]
+ osc_144 sky130_fd_sc_hs__nand2_4_47/a_27_74# sky130_fd_sc_hs__nand2_4
Xsky130_fd_sc_hs__nand2_4_58 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_4_60/Y delay_con_msb[3]
+ osc_108 sky130_fd_sc_hs__nand2_4_60/a_27_74# sky130_fd_sc_hs__nand2_4
Xsky130_fd_sc_hs__nand2_4_69 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_4_69/Y delay_con_msb[0]
+ osc_144 sky130_fd_sc_hs__nand2_4_69/a_27_74# sky130_fd_sc_hs__nand2_4
Xsky130_fd_sc_hs__einvp_4_4 DVSS DVDD DVDD DVSS pi2_l[2] sky130_fd_sc_hs__inv_8_3/A
+ sky130_fd_sc_hs__inv_4_7/Y sky130_fd_sc_hs__einvp_4_5/a_27_74# sky130_fd_sc_hs__einvp_4_5/a_27_368#
+ sky130_fd_sc_hs__einvp_4_5/a_473_323# sky130_fd_sc_hs__einvp_4
Xsky130_fd_sc_hs__and2_2_1 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__and2_2_1/A sky130_fd_sc_hs__and2_2_1/B
+ inj_out sky130_fd_sc_hs__and2_2_1/a_31_74# sky130_fd_sc_hs__and2_2_1/a_118_74# sky130_fd_sc_hs__and2_2
Xsky130_fd_sc_hs__inv_4_9 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_9/Y osc_000 sky130_fd_sc_hs__inv_4
Xsky130_fd_sc_hs__einvp_2_1 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_8_1/A sky130_fd_sc_hs__inv_4_3/Y
+ pi3_l[1] sky130_fd_sc_hs__einvp_2_1/a_263_323# sky130_fd_sc_hs__einvp_2_1/a_36_74#
+ sky130_fd_sc_hs__einvp_2_1/a_27_368# sky130_fd_sc_hs__einvp_2
Xsky130_fd_sc_hs__clkbuf_2_4 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__clkbuf_2_9/A sky130_fd_sc_hs__clkbuf_2_7/X
+ sky130_fd_sc_hs__clkbuf_2_5/a_43_192# sky130_fd_sc_hs__clkbuf_2
Xsky130_fd_sc_hs__clkbuf_2_15 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__clkbuf_2_17/A sky130_fd_sc_hs__buf_4_1/X
+ sky130_fd_sc_hs__clkbuf_2_15/a_43_192# sky130_fd_sc_hs__clkbuf_2
Xsky130_fd_sc_hs__einvp_4_19 DVSS DVDD DVDD DVSS pi5_r[2] sky130_fd_sc_hs__inv_8_9/A
+ sky130_fd_sc_hs__inv_4_21/Y sky130_fd_sc_hs__einvp_4_19/a_27_74# sky130_fd_sc_hs__einvp_4_19/a_27_368#
+ sky130_fd_sc_hs__einvp_4_19/a_473_323# sky130_fd_sc_hs__einvp_4
Xsky130_fd_sc_hs__dlygate4sd3_1_16 DVSS DVDD DVSS DVDD sky130_fd_sc_hs__clkbuf_2_1/X
+ sky130_fd_sc_hs__dlygate4sd3_1_1/A sky130_fd_sc_hs__dlygate4sd3_1_17/a_405_138#
+ sky130_fd_sc_hs__dlygate4sd3_1_17/a_28_74# sky130_fd_sc_hs__dlygate4sd3_1_17/a_289_74#
+ sky130_fd_sc_hs__dlygate4sd3_1
Xsky130_fd_sc_hs__dlygate4sd3_1_38 DVSS DVDD DVSS DVDD sky130_fd_sc_hs__dlygate4sd3_1_59/X
+ sky130_fd_sc_hs__dlygate4sd3_1_53/A sky130_fd_sc_hs__dlygate4sd3_1_39/a_405_138#
+ sky130_fd_sc_hs__dlygate4sd3_1_39/a_28_74# sky130_fd_sc_hs__dlygate4sd3_1_39/a_289_74#
+ sky130_fd_sc_hs__dlygate4sd3_1
Xsky130_fd_sc_hs__dlygate4sd3_1_49 DVSS DVDD DVSS DVDD sky130_fd_sc_hs__dlygate4sd3_1_51/X
+ sky130_fd_sc_hs__dlygate4sd3_1_49/X sky130_fd_sc_hs__dlygate4sd3_1_49/a_405_138#
+ sky130_fd_sc_hs__dlygate4sd3_1_49/a_28_74# sky130_fd_sc_hs__dlygate4sd3_1_49/a_289_74#
+ sky130_fd_sc_hs__dlygate4sd3_1
Xsky130_fd_sc_hs__dlygate4sd3_1_27 DVSS DVDD DVSS DVDD sky130_fd_sc_hs__dlygate4sd3_1_31/X
+ sky130_fd_sc_hs__dlygate4sd3_1_33/A sky130_fd_sc_hs__dlygate4sd3_1_27/a_405_138#
+ sky130_fd_sc_hs__dlygate4sd3_1_27/a_28_74# sky130_fd_sc_hs__dlygate4sd3_1_27/a_289_74#
+ sky130_fd_sc_hs__dlygate4sd3_1
Xsky130_fd_sc_hs__nand2_2_80 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_2_83/Y sky130_fd_sc_hs__nand2_2_84/B
+ osc_072 sky130_fd_sc_hs__nand2_2_83/a_27_74# sky130_fd_sc_hs__nand2_2
Xsky130_fd_sc_hs__nand2_2_91 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_2_93/Y sky130_fd_sc_hs__nand2_2_97/B
+ osc_036 sky130_fd_sc_hs__nand2_2_93/a_27_74# sky130_fd_sc_hs__nand2_2
Xsky130_fd_sc_hs__nand2_4_150 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_4_151/Y delay_con_msb[0]
+ osc_036 sky130_fd_sc_hs__nand2_4_151/a_27_74# sky130_fd_sc_hs__nand2_4
Xsky130_fd_sc_hs__nand2_2_109 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_2_109/Y sky130_fd_sc_hs__a21oi_1_49/Y
+ osc_036 sky130_fd_sc_hs__nand2_2_109/a_27_74# sky130_fd_sc_hs__nand2_2
Xsky130_fd_sc_hs__inv_16_16 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__and4_2_3/B sky130_fd_sc_hs__inv_16_31/A
+ sky130_fd_sc_hs__inv_16
Xsky130_fd_sc_hs__inv_16_27 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_16_9/A sky130_fd_sc_hs__inv_4_25/Y
+ sky130_fd_sc_hs__inv_16
Xsky130_fd_sc_hs__nand2_2_7 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_2_7/Y sky130_fd_sc_hs__nand2_2_7/B
+ osc_144 sky130_fd_sc_hs__nand2_2_7/a_27_74# sky130_fd_sc_hs__nand2_2
Xsky130_fd_sc_hs__conb_1_0 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__conb_1_1/LO sky130_fd_sc_hs__dfrtp_4_3/D
+ sky130_fd_sc_hs__conb_1_1/a_165_290# sky130_fd_sc_hs__conb_1_1/a_21_290# sky130_fd_sc_hs__conb_1
Xsky130_fd_sc_hs__nand2_4_15 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_4_15/Y delay_con_msb[1]
+ osc_000 sky130_fd_sc_hs__nand2_4_15/a_27_74# sky130_fd_sc_hs__nand2_4
Xsky130_fd_sc_hs__nand2_4_26 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_4_27/Y delay_con_msb[1]
+ osc_144 sky130_fd_sc_hs__nand2_4_27/a_27_74# sky130_fd_sc_hs__nand2_4
Xsky130_fd_sc_hs__nand2_4_37 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_4_40/Y delay_con_msb[2]
+ osc_000 sky130_fd_sc_hs__nand2_4_40/a_27_74# sky130_fd_sc_hs__nand2_4
Xsky130_fd_sc_hs__nand2_4_48 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_4_49/Y delay_con_msb[0]
+ osc_000 sky130_fd_sc_hs__nand2_4_49/a_27_74# sky130_fd_sc_hs__nand2_4
Xsky130_fd_sc_hs__nand2_4_59 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_4_61/Y delay_con_msb[3]
+ osc_108 sky130_fd_sc_hs__nand2_4_61/a_27_74# sky130_fd_sc_hs__nand2_4
Xsky130_fd_sc_hs__einvp_4_5 DVSS DVDD DVDD DVSS pi2_l[2] sky130_fd_sc_hs__inv_8_3/A
+ sky130_fd_sc_hs__inv_4_7/Y sky130_fd_sc_hs__einvp_4_5/a_27_74# sky130_fd_sc_hs__einvp_4_5/a_27_368#
+ sky130_fd_sc_hs__einvp_4_5/a_473_323# sky130_fd_sc_hs__einvp_4
Xsky130_fd_sc_hs__and2_2_2 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__and2_2_3/A sky130_fd_sc_hs__and2_2_3/B
+ sky130_fd_sc_hs__and2_2_3/X sky130_fd_sc_hs__and2_2_3/a_31_74# sky130_fd_sc_hs__and2_2_3/a_118_74#
+ sky130_fd_sc_hs__and2_2
Xsky130_fd_sc_hs__einvp_2_2 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_8_1/A sky130_fd_sc_hs__inv_4_5/Y
+ pi3_r[1] sky130_fd_sc_hs__einvp_2_3/a_263_323# sky130_fd_sc_hs__einvp_2_3/a_36_74#
+ sky130_fd_sc_hs__einvp_2_3/a_27_368# sky130_fd_sc_hs__einvp_2
Xsky130_fd_sc_hs__clkbuf_2_5 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__clkbuf_2_9/A sky130_fd_sc_hs__clkbuf_2_7/X
+ sky130_fd_sc_hs__clkbuf_2_5/a_43_192# sky130_fd_sc_hs__clkbuf_2
Xsky130_fd_sc_hs__clkbuf_2_16 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__clkbuf_2_3/A sky130_fd_sc_hs__clkbuf_2_17/A
+ sky130_fd_sc_hs__clkbuf_2_17/a_43_192# sky130_fd_sc_hs__clkbuf_2
Xsky130_fd_sc_hs__dlygate4sd3_1_17 DVSS DVDD DVSS DVDD sky130_fd_sc_hs__clkbuf_2_1/X
+ sky130_fd_sc_hs__dlygate4sd3_1_1/A sky130_fd_sc_hs__dlygate4sd3_1_17/a_405_138#
+ sky130_fd_sc_hs__dlygate4sd3_1_17/a_28_74# sky130_fd_sc_hs__dlygate4sd3_1_17/a_289_74#
+ sky130_fd_sc_hs__dlygate4sd3_1
Xsky130_fd_sc_hs__dlygate4sd3_1_39 DVSS DVDD DVSS DVDD sky130_fd_sc_hs__dlygate4sd3_1_59/X
+ sky130_fd_sc_hs__dlygate4sd3_1_53/A sky130_fd_sc_hs__dlygate4sd3_1_39/a_405_138#
+ sky130_fd_sc_hs__dlygate4sd3_1_39/a_28_74# sky130_fd_sc_hs__dlygate4sd3_1_39/a_289_74#
+ sky130_fd_sc_hs__dlygate4sd3_1
Xsky130_fd_sc_hs__dlygate4sd3_1_28 DVSS DVDD DVSS DVDD sky130_fd_sc_hs__dlygate4sd3_1_35/X
+ sky130_fd_sc_hs__dlygate4sd3_1_37/A sky130_fd_sc_hs__dlygate4sd3_1_29/a_405_138#
+ sky130_fd_sc_hs__dlygate4sd3_1_29/a_28_74# sky130_fd_sc_hs__dlygate4sd3_1_29/a_289_74#
+ sky130_fd_sc_hs__dlygate4sd3_1
Xsky130_fd_sc_hs__nand2_2_70 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_2_71/Y sky130_fd_sc_hs__nand2_2_71/B
+ osc_144 sky130_fd_sc_hs__nand2_2_71/a_27_74# sky130_fd_sc_hs__nand2_2
Xsky130_fd_sc_hs__nand2_2_81 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_2_84/Y sky130_fd_sc_hs__nand2_2_84/B
+ osc_072 sky130_fd_sc_hs__nand2_2_84/a_27_74# sky130_fd_sc_hs__nand2_2
Xsky130_fd_sc_hs__nand2_2_92 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_2_92/Y sky130_fd_sc_hs__nand2_2_97/B
+ osc_036 sky130_fd_sc_hs__nand2_2_92/a_27_74# sky130_fd_sc_hs__nand2_2
Xsky130_fd_sc_hs__nand2_4_140 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_4_141/Y delay_con_msb[3]
+ osc_036 sky130_fd_sc_hs__nand2_4_141/a_27_74# sky130_fd_sc_hs__nand2_4
Xsky130_fd_sc_hs__nand2_4_151 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_4_151/Y delay_con_msb[0]
+ osc_036 sky130_fd_sc_hs__nand2_4_151/a_27_74# sky130_fd_sc_hs__nand2_4
Xsky130_fd_sc_hs__inv_16_17 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__and4_2_3/B sky130_fd_sc_hs__inv_16_31/A
+ sky130_fd_sc_hs__inv_16
Xsky130_fd_sc_hs__inv_16_28 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__and4_2_3/C sky130_fd_sc_hs__inv_16_31/A
+ sky130_fd_sc_hs__inv_16
Xsky130_fd_sc_hs__nand2_2_8 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_2_9/Y sky130_fd_sc_hs__nand2_2_9/B
+ osc_000 sky130_fd_sc_hs__nand2_2_9/a_27_74# sky130_fd_sc_hs__nand2_2
Xsky130_fd_sc_hs__conb_1_1 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__conb_1_1/LO sky130_fd_sc_hs__dfrtp_4_3/D
+ sky130_fd_sc_hs__conb_1_1/a_165_290# sky130_fd_sc_hs__conb_1_1/a_21_290# sky130_fd_sc_hs__conb_1
Xsky130_fd_sc_hs__nand2_4_16 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_4_17/Y delay_con_msb[1]
+ osc_144 sky130_fd_sc_hs__nand2_4_17/a_27_74# sky130_fd_sc_hs__nand2_4
Xsky130_fd_sc_hs__nand2_4_27 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_4_27/Y delay_con_msb[1]
+ osc_144 sky130_fd_sc_hs__nand2_4_27/a_27_74# sky130_fd_sc_hs__nand2_4
Xsky130_fd_sc_hs__nand2_4_38 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_4_41/Y delay_con_msb[3]
+ osc_000 sky130_fd_sc_hs__nand2_4_41/a_27_74# sky130_fd_sc_hs__nand2_4
Xsky130_fd_sc_hs__nand2_4_49 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_4_49/Y delay_con_msb[0]
+ osc_000 sky130_fd_sc_hs__nand2_4_49/a_27_74# sky130_fd_sc_hs__nand2_4
Xsky130_fd_sc_hs__einvp_4_6 DVSS DVDD DVDD DVSS pi2_r[2] sky130_fd_sc_hs__inv_8_3/A
+ sky130_fd_sc_hs__inv_4_9/Y sky130_fd_sc_hs__einvp_4_7/a_27_74# sky130_fd_sc_hs__einvp_4_7/a_27_368#
+ sky130_fd_sc_hs__einvp_4_7/a_473_323# sky130_fd_sc_hs__einvp_4
Xsky130_fd_sc_hs__and2_2_3 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__and2_2_3/A sky130_fd_sc_hs__and2_2_3/B
+ sky130_fd_sc_hs__and2_2_3/X sky130_fd_sc_hs__and2_2_3/a_31_74# sky130_fd_sc_hs__and2_2_3/a_118_74#
+ sky130_fd_sc_hs__and2_2
Xsky130_fd_sc_hs__einvp_2_3 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_8_1/A sky130_fd_sc_hs__inv_4_5/Y
+ pi3_r[1] sky130_fd_sc_hs__einvp_2_3/a_263_323# sky130_fd_sc_hs__einvp_2_3/a_36_74#
+ sky130_fd_sc_hs__einvp_2_3/a_27_368# sky130_fd_sc_hs__einvp_2
Xsky130_fd_sc_hs__clkbuf_2_6 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__clkbuf_2_7/X glob_en
+ sky130_fd_sc_hs__clkbuf_2_7/a_43_192# sky130_fd_sc_hs__clkbuf_2
Xsky130_fd_sc_hs__clkbuf_2_17 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__clkbuf_2_3/A sky130_fd_sc_hs__clkbuf_2_17/A
+ sky130_fd_sc_hs__clkbuf_2_17/a_43_192# sky130_fd_sc_hs__clkbuf_2
Xsky130_fd_sc_hs__dlygate4sd3_1_18 DVSS DVDD DVSS DVDD sky130_fd_sc_hs__dlygate4sd3_1_20/A
+ sky130_fd_sc_hs__dlygate4sd3_1_9/A sky130_fd_sc_hs__dlygate4sd3_1_20/a_405_138#
+ sky130_fd_sc_hs__dlygate4sd3_1_20/a_28_74# sky130_fd_sc_hs__dlygate4sd3_1_20/a_289_74#
+ sky130_fd_sc_hs__dlygate4sd3_1
Xsky130_fd_sc_hs__dlygate4sd3_1_29 DVSS DVDD DVSS DVDD sky130_fd_sc_hs__dlygate4sd3_1_35/X
+ sky130_fd_sc_hs__dlygate4sd3_1_37/A sky130_fd_sc_hs__dlygate4sd3_1_29/a_405_138#
+ sky130_fd_sc_hs__dlygate4sd3_1_29/a_28_74# sky130_fd_sc_hs__dlygate4sd3_1_29/a_289_74#
+ sky130_fd_sc_hs__dlygate4sd3_1
Xsky130_fd_sc_hs__nand2_2_60 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_2_61/Y sky130_fd_sc_hs__nand2_2_61/B
+ osc_108 sky130_fd_sc_hs__nand2_2_61/a_27_74# sky130_fd_sc_hs__nand2_2
Xsky130_fd_sc_hs__nand2_2_71 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_2_71/Y sky130_fd_sc_hs__nand2_2_71/B
+ osc_144 sky130_fd_sc_hs__nand2_2_71/a_27_74# sky130_fd_sc_hs__nand2_2
Xsky130_fd_sc_hs__nand2_2_82 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_2_85/Y sky130_fd_sc_hs__nand2_2_85/B
+ osc_072 sky130_fd_sc_hs__nand2_2_85/a_27_74# sky130_fd_sc_hs__nand2_2
Xsky130_fd_sc_hs__nand2_4_130 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_4_131/Y delay_con_msb[3]
+ osc_072 sky130_fd_sc_hs__nand2_4_131/a_27_74# sky130_fd_sc_hs__nand2_4
Xsky130_fd_sc_hs__nand2_4_141 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_4_141/Y delay_con_msb[3]
+ osc_036 sky130_fd_sc_hs__nand2_4_141/a_27_74# sky130_fd_sc_hs__nand2_4
Xsky130_fd_sc_hs__nand2_2_93 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_2_93/Y sky130_fd_sc_hs__nand2_2_97/B
+ osc_036 sky130_fd_sc_hs__nand2_2_93/a_27_74# sky130_fd_sc_hs__nand2_2
Xsky130_fd_sc_hs__nand2_4_152 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_4_153/Y delay_con_msb[1]
+ osc_036 sky130_fd_sc_hs__nand2_4_153/a_27_74# sky130_fd_sc_hs__nand2_4
Xsky130_fd_sc_hs__inv_16_18 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__and4_2_5/D sky130_fd_sc_hs__inv_16_7/Y
+ sky130_fd_sc_hs__inv_16
Xsky130_fd_sc_hs__inv_16_29 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__and4_2_3/D sky130_fd_sc_hs__inv_16_31/A
+ sky130_fd_sc_hs__inv_16
Xsky130_fd_sc_hs__nand2_2_9 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_2_9/Y sky130_fd_sc_hs__nand2_2_9/B
+ osc_000 sky130_fd_sc_hs__nand2_2_9/a_27_74# sky130_fd_sc_hs__nand2_2
Xsky130_fd_sc_hs__nand2_4_17 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_4_17/Y delay_con_msb[1]
+ osc_144 sky130_fd_sc_hs__nand2_4_17/a_27_74# sky130_fd_sc_hs__nand2_4
Xsky130_fd_sc_hs__nand2_4_28 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_4_29/Y delay_con_msb[2]
+ osc_000 sky130_fd_sc_hs__nand2_4_29/a_27_74# sky130_fd_sc_hs__nand2_4
Xsky130_fd_sc_hs__nand2_4_39 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_4_39/Y delay_con_msb[2]
+ osc_000 sky130_fd_sc_hs__nand2_4_39/a_27_74# sky130_fd_sc_hs__nand2_4
Xsky130_fd_sc_hs__einvp_4_7 DVSS DVDD DVDD DVSS pi2_r[2] sky130_fd_sc_hs__inv_8_3/A
+ sky130_fd_sc_hs__inv_4_9/Y sky130_fd_sc_hs__einvp_4_7/a_27_74# sky130_fd_sc_hs__einvp_4_7/a_27_368#
+ sky130_fd_sc_hs__einvp_4_7/a_473_323# sky130_fd_sc_hs__einvp_4
Xsky130_fd_sc_hs__einvp_2_10 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_8_5/A sky130_fd_sc_hs__inv_4_13/Y
+ pi4_r[1] sky130_fd_sc_hs__einvp_2_11/a_263_323# sky130_fd_sc_hs__einvp_2_11/a_36_74#
+ sky130_fd_sc_hs__einvp_2_11/a_27_368# sky130_fd_sc_hs__einvp_2
Xsky130_fd_sc_hs__dfrtp_4_0 DVSS DVDD sky130_fd_sc_hs__and4_2_3/X DVDD DVSS sky130_fd_sc_hs__dfrtp_4_3/D
+ sky130_fd_sc_hs__inv_4_1/Y sky130_fd_sc_hs__and2_2_3/B sky130_fd_sc_hs__dfrtp_4_1/a_37_78#
+ sky130_fd_sc_hs__dfrtp_4_1/a_494_366# sky130_fd_sc_hs__dfrtp_4_1/a_699_463# sky130_fd_sc_hs__dfrtp_4_1/a_313_74#
+ sky130_fd_sc_hs__dfrtp_4_1/a_1627_493# sky130_fd_sc_hs__dfrtp_4_1/a_1678_395# sky130_fd_sc_hs__dfrtp_4_1/a_1827_81#
+ sky130_fd_sc_hs__dfrtp_4_1/a_789_463# sky130_fd_sc_hs__dfrtp_4_1/a_1350_392# sky130_fd_sc_hs__dfrtp_4_1/a_834_355#
+ sky130_fd_sc_hs__dfrtp_4_1/a_812_138# sky130_fd_sc_hs__dfrtp_4_1/a_124_78# sky130_fd_sc_hs__dfrtp_4_1/a_1647_81#
+ sky130_fd_sc_hs__dfrtp_4_1/a_2010_409# sky130_fd_sc_hs__dfrtp_4_1/a_890_138# sky130_fd_sc_hs__dfrtp_4
Xsky130_fd_sc_hs__einvp_2_4 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_8_3/A sky130_fd_sc_hs__inv_4_7/Y
+ pi2_l[1] sky130_fd_sc_hs__einvp_2_5/a_263_323# sky130_fd_sc_hs__einvp_2_5/a_36_74#
+ sky130_fd_sc_hs__einvp_2_5/a_27_368# sky130_fd_sc_hs__einvp_2
Xsky130_fd_sc_hs__clkbuf_2_7 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__clkbuf_2_7/X glob_en
+ sky130_fd_sc_hs__clkbuf_2_7/a_43_192# sky130_fd_sc_hs__clkbuf_2
Xsky130_fd_sc_hs__dlygate4sd3_1_19 DVSS DVDD DVSS DVDD sky130_fd_sc_hs__dlygate4sd3_1_1/X
+ sky130_fd_sc_hs__dlygate4sd3_1_3/A sky130_fd_sc_hs__dlygate4sd3_1_21/a_405_138#
+ sky130_fd_sc_hs__dlygate4sd3_1_21/a_28_74# sky130_fd_sc_hs__dlygate4sd3_1_21/a_289_74#
+ sky130_fd_sc_hs__dlygate4sd3_1
Xsky130_fd_sc_hs__nand2_2_50 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_2_51/Y sky130_fd_sc_hs__nand2_2_65/B
+ osc_144 sky130_fd_sc_hs__nand2_2_51/a_27_74# sky130_fd_sc_hs__nand2_2
Xsky130_fd_sc_hs__nand2_2_61 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_2_61/Y sky130_fd_sc_hs__nand2_2_61/B
+ osc_108 sky130_fd_sc_hs__nand2_2_61/a_27_74# sky130_fd_sc_hs__nand2_2
Xsky130_fd_sc_hs__nand2_2_72 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_2_73/Y sky130_fd_sc_hs__nand2_2_73/B
+ osc_108 sky130_fd_sc_hs__nand2_2_73/a_27_74# sky130_fd_sc_hs__nand2_2
Xsky130_fd_sc_hs__nand2_4_120 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_4_121/Y delay_con_msb[3]
+ osc_072 sky130_fd_sc_hs__nand2_4_121/a_27_74# sky130_fd_sc_hs__nand2_4
Xsky130_fd_sc_hs__nand2_2_83 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_2_83/Y sky130_fd_sc_hs__nand2_2_84/B
+ osc_072 sky130_fd_sc_hs__nand2_2_83/a_27_74# sky130_fd_sc_hs__nand2_2
Xsky130_fd_sc_hs__nand2_4_131 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_4_131/Y delay_con_msb[3]
+ osc_072 sky130_fd_sc_hs__nand2_4_131/a_27_74# sky130_fd_sc_hs__nand2_4
Xsky130_fd_sc_hs__nand2_4_142 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_4_143/Y delay_con_msb[1]
+ osc_036 sky130_fd_sc_hs__nand2_4_143/a_27_74# sky130_fd_sc_hs__nand2_4
Xsky130_fd_sc_hs__nand2_2_94 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_2_96/Y sky130_fd_sc_hs__nand2_2_99/B
+ osc_036 sky130_fd_sc_hs__nand2_2_96/a_27_74# sky130_fd_sc_hs__nand2_2
Xsky130_fd_sc_hs__nand2_4_153 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_4_153/Y delay_con_msb[1]
+ osc_036 sky130_fd_sc_hs__nand2_4_153/a_27_74# sky130_fd_sc_hs__nand2_4
Xsky130_fd_sc_hs__inv_16_19 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__and4_2_5/D sky130_fd_sc_hs__inv_16_7/Y
+ sky130_fd_sc_hs__inv_16
Xsky130_fd_sc_hs__nand2_4_18 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_4_19/Y delay_con_msb[2]
+ osc_144 sky130_fd_sc_hs__nand2_4_19/a_27_74# sky130_fd_sc_hs__nand2_4
Xsky130_fd_sc_hs__nand2_4_29 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_4_29/Y delay_con_msb[2]
+ osc_000 sky130_fd_sc_hs__nand2_4_29/a_27_74# sky130_fd_sc_hs__nand2_4
Xsky130_fd_sc_hs__einvp_4_8 DVSS DVDD DVDD DVSS pi4_l[2] sky130_fd_sc_hs__inv_8_5/A
+ sky130_fd_sc_hs__inv_4_11/Y sky130_fd_sc_hs__einvp_4_9/a_27_74# sky130_fd_sc_hs__einvp_4_9/a_27_368#
+ sky130_fd_sc_hs__einvp_4_9/a_473_323# sky130_fd_sc_hs__einvp_4
Xsky130_fd_sc_hs__einvp_2_11 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_8_5/A sky130_fd_sc_hs__inv_4_13/Y
+ pi4_r[1] sky130_fd_sc_hs__einvp_2_11/a_263_323# sky130_fd_sc_hs__einvp_2_11/a_36_74#
+ sky130_fd_sc_hs__einvp_2_11/a_27_368# sky130_fd_sc_hs__einvp_2
Xsky130_fd_sc_hs__dfrtp_4_1 DVSS DVDD sky130_fd_sc_hs__and4_2_3/X DVDD DVSS sky130_fd_sc_hs__dfrtp_4_3/D
+ sky130_fd_sc_hs__inv_4_1/Y sky130_fd_sc_hs__and2_2_3/B sky130_fd_sc_hs__dfrtp_4_1/a_37_78#
+ sky130_fd_sc_hs__dfrtp_4_1/a_494_366# sky130_fd_sc_hs__dfrtp_4_1/a_699_463# sky130_fd_sc_hs__dfrtp_4_1/a_313_74#
+ sky130_fd_sc_hs__dfrtp_4_1/a_1627_493# sky130_fd_sc_hs__dfrtp_4_1/a_1678_395# sky130_fd_sc_hs__dfrtp_4_1/a_1827_81#
+ sky130_fd_sc_hs__dfrtp_4_1/a_789_463# sky130_fd_sc_hs__dfrtp_4_1/a_1350_392# sky130_fd_sc_hs__dfrtp_4_1/a_834_355#
+ sky130_fd_sc_hs__dfrtp_4_1/a_812_138# sky130_fd_sc_hs__dfrtp_4_1/a_124_78# sky130_fd_sc_hs__dfrtp_4_1/a_1647_81#
+ sky130_fd_sc_hs__dfrtp_4_1/a_2010_409# sky130_fd_sc_hs__dfrtp_4_1/a_890_138# sky130_fd_sc_hs__dfrtp_4
Xsky130_fd_sc_hs__einvp_2_5 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_8_3/A sky130_fd_sc_hs__inv_4_7/Y
+ pi2_l[1] sky130_fd_sc_hs__einvp_2_5/a_263_323# sky130_fd_sc_hs__einvp_2_5/a_36_74#
+ sky130_fd_sc_hs__einvp_2_5/a_27_368# sky130_fd_sc_hs__einvp_2
Xsky130_fd_sc_hs__clkbuf_2_8 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__buf_4_1/A sky130_fd_sc_hs__clkbuf_2_8/A
+ sky130_fd_sc_hs__clkbuf_2_8/a_43_192# sky130_fd_sc_hs__clkbuf_2
Xsky130_fd_sc_hs__einvp_8_10 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_8_5/A pi4_l[3]
+ sky130_fd_sc_hs__inv_4_11/Y sky130_fd_sc_hs__einvp_8_8/a_802_323# sky130_fd_sc_hs__einvp_8_8/a_27_74#
+ sky130_fd_sc_hs__einvp_8_8/a_27_368# sky130_fd_sc_hs__einvp_8
Xsky130_fd_sc_hs__nand2_2_40 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_2_42/Y sky130_fd_sc_hs__nand2_2_61/B
+ osc_108 sky130_fd_sc_hs__nand2_2_42/a_27_74# sky130_fd_sc_hs__nand2_2
Xsky130_fd_sc_hs__nand2_2_51 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_2_51/Y sky130_fd_sc_hs__nand2_2_65/B
+ osc_144 sky130_fd_sc_hs__nand2_2_51/a_27_74# sky130_fd_sc_hs__nand2_2
Xsky130_fd_sc_hs__nand2_2_62 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_2_63/Y sky130_fd_sc_hs__nand2_2_73/B
+ osc_108 sky130_fd_sc_hs__nand2_2_63/a_27_74# sky130_fd_sc_hs__nand2_2
Xsky130_fd_sc_hs__nand2_2_73 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_2_73/Y sky130_fd_sc_hs__nand2_2_73/B
+ osc_108 sky130_fd_sc_hs__nand2_2_73/a_27_74# sky130_fd_sc_hs__nand2_2
Xsky130_fd_sc_hs__nand2_4_110 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_4_110/Y delay_con_msb[1]
+ osc_072 sky130_fd_sc_hs__nand2_4_110/a_27_74# sky130_fd_sc_hs__nand2_4
Xsky130_fd_sc_hs__nand2_4_121 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_4_121/Y delay_con_msb[3]
+ osc_072 sky130_fd_sc_hs__nand2_4_121/a_27_74# sky130_fd_sc_hs__nand2_4
Xsky130_fd_sc_hs__nand2_2_84 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_2_84/Y sky130_fd_sc_hs__nand2_2_84/B
+ osc_072 sky130_fd_sc_hs__nand2_2_84/a_27_74# sky130_fd_sc_hs__nand2_2
Xsky130_fd_sc_hs__nand2_4_132 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_4_133/Y delay_con_msb[0]
+ osc_036 sky130_fd_sc_hs__nand2_4_133/a_27_74# sky130_fd_sc_hs__nand2_4
Xsky130_fd_sc_hs__nand2_4_143 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_4_143/Y delay_con_msb[1]
+ osc_036 sky130_fd_sc_hs__nand2_4_143/a_27_74# sky130_fd_sc_hs__nand2_4
Xsky130_fd_sc_hs__nand2_2_95 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_2_97/Y sky130_fd_sc_hs__nand2_2_97/B
+ osc_036 sky130_fd_sc_hs__nand2_2_97/a_27_74# sky130_fd_sc_hs__nand2_2
Xsky130_fd_sc_hs__nand2_4_154 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_4_155/Y delay_con_msb[3]
+ osc_036 sky130_fd_sc_hs__nand2_4_155/a_27_74# sky130_fd_sc_hs__nand2_4
Xsky130_fd_sc_hs__diode_2_0 sky130_fd_sc_hs__clkbuf_4_1/A DVSS DVDD DVDD DVSS sky130_fd_sc_hs__diode_2
Xsky130_fd_sc_hs__nand2_4_19 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_4_19/Y delay_con_msb[2]
+ osc_144 sky130_fd_sc_hs__nand2_4_19/a_27_74# sky130_fd_sc_hs__nand2_4
Xsky130_fd_sc_hs__einvp_4_9 DVSS DVDD DVDD DVSS pi4_l[2] sky130_fd_sc_hs__inv_8_5/A
+ sky130_fd_sc_hs__inv_4_11/Y sky130_fd_sc_hs__einvp_4_9/a_27_74# sky130_fd_sc_hs__einvp_4_9/a_27_368#
+ sky130_fd_sc_hs__einvp_4_9/a_473_323# sky130_fd_sc_hs__einvp_4
Xsky130_fd_sc_hs__einvp_2_12 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_8_7/A sky130_fd_sc_hs__inv_4_15/Y
+ pi1_l[1] sky130_fd_sc_hs__einvp_2_13/a_263_323# sky130_fd_sc_hs__einvp_2_13/a_36_74#
+ sky130_fd_sc_hs__einvp_2_13/a_27_368# sky130_fd_sc_hs__einvp_2
Xsky130_fd_sc_hs__dfrtp_4_2 DVSS DVDD sky130_fd_sc_hs__and4_2_3/X DVDD DVSS sky130_fd_sc_hs__dfrtp_4_3/D
+ sky130_fd_sc_hs__inv_4_1/Y sky130_fd_sc_hs__and2_2_3/A sky130_fd_sc_hs__dfrtp_4_3/a_37_78#
+ sky130_fd_sc_hs__dfrtp_4_3/a_494_366# sky130_fd_sc_hs__dfrtp_4_3/a_699_463# sky130_fd_sc_hs__dfrtp_4_3/a_313_74#
+ sky130_fd_sc_hs__dfrtp_4_3/a_1627_493# sky130_fd_sc_hs__dfrtp_4_3/a_1678_395# sky130_fd_sc_hs__dfrtp_4_3/a_1827_81#
+ sky130_fd_sc_hs__dfrtp_4_3/a_789_463# sky130_fd_sc_hs__dfrtp_4_3/a_1350_392# sky130_fd_sc_hs__dfrtp_4_3/a_834_355#
+ sky130_fd_sc_hs__dfrtp_4_3/a_812_138# sky130_fd_sc_hs__dfrtp_4_3/a_124_78# sky130_fd_sc_hs__dfrtp_4_3/a_1647_81#
+ sky130_fd_sc_hs__dfrtp_4_3/a_2010_409# sky130_fd_sc_hs__dfrtp_4_3/a_890_138# sky130_fd_sc_hs__dfrtp_4
Xsky130_fd_sc_hs__einvp_2_6 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_8_3/A sky130_fd_sc_hs__inv_4_9/Y
+ pi2_r[1] sky130_fd_sc_hs__einvp_2_7/a_263_323# sky130_fd_sc_hs__einvp_2_7/a_36_74#
+ sky130_fd_sc_hs__einvp_2_7/a_27_368# sky130_fd_sc_hs__einvp_2
Xsky130_fd_sc_hs__clkbuf_2_9 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__clkbuf_4_5/A sky130_fd_sc_hs__clkbuf_2_9/A
+ sky130_fd_sc_hs__clkbuf_2_9/a_43_192# sky130_fd_sc_hs__clkbuf_2
Xsky130_fd_sc_hs__einvp_8_11 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_8_5/A pi4_r[3]
+ sky130_fd_sc_hs__inv_4_13/Y sky130_fd_sc_hs__einvp_8_9/a_802_323# sky130_fd_sc_hs__einvp_8_9/a_27_74#
+ sky130_fd_sc_hs__einvp_8_9/a_27_368# sky130_fd_sc_hs__einvp_8
Xsky130_fd_sc_hs__nand2_2_30 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_2_31/Y sky130_fd_sc_hs__nand2_2_7/B
+ osc_144 sky130_fd_sc_hs__nand2_2_31/a_27_74# sky130_fd_sc_hs__nand2_2
Xsky130_fd_sc_hs__nand2_2_41 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_2_43/Y sky130_fd_sc_hs__nand2_2_43/B
+ osc_108 sky130_fd_sc_hs__nand2_2_43/a_27_74# sky130_fd_sc_hs__nand2_2
Xsky130_fd_sc_hs__nand2_2_52 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_2_53/Y sky130_fd_sc_hs__nand2_2_85/B
+ osc_072 sky130_fd_sc_hs__nand2_2_53/a_27_74# sky130_fd_sc_hs__nand2_2
Xsky130_fd_sc_hs__nand2_2_63 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_2_63/Y sky130_fd_sc_hs__nand2_2_73/B
+ osc_108 sky130_fd_sc_hs__nand2_2_63/a_27_74# sky130_fd_sc_hs__nand2_2
Xsky130_fd_sc_hs__nand2_4_100 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_4_102/Y delay_con_msb[0]
+ osc_072 sky130_fd_sc_hs__nand2_4_102/a_27_74# sky130_fd_sc_hs__nand2_4
Xsky130_fd_sc_hs__nand2_2_74 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_2_77/Y sky130_fd_sc_hs__nand2_2_79/B
+ osc_072 sky130_fd_sc_hs__nand2_2_77/a_27_74# sky130_fd_sc_hs__nand2_2
Xsky130_fd_sc_hs__nand2_2_85 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_2_85/Y sky130_fd_sc_hs__nand2_2_85/B
+ osc_072 sky130_fd_sc_hs__nand2_2_85/a_27_74# sky130_fd_sc_hs__nand2_2
Xsky130_fd_sc_hs__nand2_2_96 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_2_96/Y sky130_fd_sc_hs__nand2_2_99/B
+ osc_036 sky130_fd_sc_hs__nand2_2_96/a_27_74# sky130_fd_sc_hs__nand2_2
Xsky130_fd_sc_hs__nand2_4_111 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_4_111/Y delay_con_msb[1]
+ osc_072 sky130_fd_sc_hs__nand2_4_111/a_27_74# sky130_fd_sc_hs__nand2_4
Xsky130_fd_sc_hs__nand2_4_122 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_4_123/Y delay_con_msb[1]
+ osc_072 sky130_fd_sc_hs__nand2_4_123/a_27_74# sky130_fd_sc_hs__nand2_4
Xsky130_fd_sc_hs__nand2_4_133 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_4_133/Y delay_con_msb[0]
+ osc_036 sky130_fd_sc_hs__nand2_4_133/a_27_74# sky130_fd_sc_hs__nand2_4
Xsky130_fd_sc_hs__nand2_4_144 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_4_145/Y delay_con_msb[2]
+ osc_036 sky130_fd_sc_hs__nand2_4_145/a_27_74# sky130_fd_sc_hs__nand2_4
Xsky130_fd_sc_hs__nand2_4_155 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_4_155/Y delay_con_msb[3]
+ osc_036 sky130_fd_sc_hs__nand2_4_155/a_27_74# sky130_fd_sc_hs__nand2_4
Xsky130_fd_sc_hs__diode_2_1 sky130_fd_sc_hs__clkbuf_4_1/A DVSS DVDD DVDD DVSS sky130_fd_sc_hs__diode_2
Xsky130_fd_sc_hs__nand2_8_40 DVSS DVDD DVDD DVSS inj_out osc_072 osc_108 sky130_fd_sc_hs__nand2_8_41/a_27_74#
+ sky130_fd_sc_hs__nand2_8
Xsky130_fd_sc_hs__einvp_2_13 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_8_7/A sky130_fd_sc_hs__inv_4_15/Y
+ pi1_l[1] sky130_fd_sc_hs__einvp_2_13/a_263_323# sky130_fd_sc_hs__einvp_2_13/a_36_74#
+ sky130_fd_sc_hs__einvp_2_13/a_27_368# sky130_fd_sc_hs__einvp_2
Xsky130_fd_sc_hs__dfrtp_4_3 DVSS DVDD sky130_fd_sc_hs__and4_2_3/X DVDD DVSS sky130_fd_sc_hs__dfrtp_4_3/D
+ sky130_fd_sc_hs__inv_4_1/Y sky130_fd_sc_hs__and2_2_3/A sky130_fd_sc_hs__dfrtp_4_3/a_37_78#
+ sky130_fd_sc_hs__dfrtp_4_3/a_494_366# sky130_fd_sc_hs__dfrtp_4_3/a_699_463# sky130_fd_sc_hs__dfrtp_4_3/a_313_74#
+ sky130_fd_sc_hs__dfrtp_4_3/a_1627_493# sky130_fd_sc_hs__dfrtp_4_3/a_1678_395# sky130_fd_sc_hs__dfrtp_4_3/a_1827_81#
+ sky130_fd_sc_hs__dfrtp_4_3/a_789_463# sky130_fd_sc_hs__dfrtp_4_3/a_1350_392# sky130_fd_sc_hs__dfrtp_4_3/a_834_355#
+ sky130_fd_sc_hs__dfrtp_4_3/a_812_138# sky130_fd_sc_hs__dfrtp_4_3/a_124_78# sky130_fd_sc_hs__dfrtp_4_3/a_1647_81#
+ sky130_fd_sc_hs__dfrtp_4_3/a_2010_409# sky130_fd_sc_hs__dfrtp_4_3/a_890_138# sky130_fd_sc_hs__dfrtp_4
Xsky130_fd_sc_hs__inv_4_30 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_31/Y delay_con_lsb[4]
+ sky130_fd_sc_hs__inv_4
Xsky130_fd_sc_hs__einvp_2_7 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_8_3/A sky130_fd_sc_hs__inv_4_9/Y
+ pi2_r[1] sky130_fd_sc_hs__einvp_2_7/a_263_323# sky130_fd_sc_hs__einvp_2_7/a_36_74#
+ sky130_fd_sc_hs__einvp_2_7/a_27_368# sky130_fd_sc_hs__einvp_2
Xsky130_fd_sc_hs__einvp_8_12 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_8_7/A pi1_l[3]
+ sky130_fd_sc_hs__inv_4_15/Y sky130_fd_sc_hs__einvp_8_14/a_802_323# sky130_fd_sc_hs__einvp_8_14/a_27_74#
+ sky130_fd_sc_hs__einvp_8_14/a_27_368# sky130_fd_sc_hs__einvp_8
Xsky130_fd_sc_hs__nand2_2_20 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_2_21/Y sky130_fd_sc_hs__nand2_2_7/B
+ osc_144 sky130_fd_sc_hs__nand2_2_21/a_27_74# sky130_fd_sc_hs__nand2_2
Xsky130_fd_sc_hs__nand2_2_31 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_2_31/Y sky130_fd_sc_hs__nand2_2_7/B
+ osc_144 sky130_fd_sc_hs__nand2_2_31/a_27_74# sky130_fd_sc_hs__nand2_2
Xsky130_fd_sc_hs__nand2_2_42 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_2_42/Y sky130_fd_sc_hs__nand2_2_61/B
+ osc_108 sky130_fd_sc_hs__nand2_2_42/a_27_74# sky130_fd_sc_hs__nand2_2
Xsky130_fd_sc_hs__nand2_2_53 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_2_53/Y sky130_fd_sc_hs__nand2_2_85/B
+ osc_072 sky130_fd_sc_hs__nand2_2_53/a_27_74# sky130_fd_sc_hs__nand2_2
Xsky130_fd_sc_hs__nand2_2_64 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_2_65/Y sky130_fd_sc_hs__nand2_2_65/B
+ osc_144 sky130_fd_sc_hs__nand2_2_65/a_27_74# sky130_fd_sc_hs__nand2_2
Xsky130_fd_sc_hs__nand2_4_101 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_4_103/Y delay_con_msb[0]
+ osc_072 sky130_fd_sc_hs__nand2_4_103/a_27_74# sky130_fd_sc_hs__nand2_4
Xsky130_fd_sc_hs__nand2_4_112 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_4_113/Y delay_con_msb[2]
+ osc_072 sky130_fd_sc_hs__nand2_4_113/a_27_74# sky130_fd_sc_hs__nand2_4
Xsky130_fd_sc_hs__nand2_2_75 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_2_78/Y sky130_fd_sc_hs__nand2_2_79/B
+ osc_072 sky130_fd_sc_hs__nand2_2_78/a_27_74# sky130_fd_sc_hs__nand2_2
Xsky130_fd_sc_hs__nand2_4_123 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_4_123/Y delay_con_msb[1]
+ osc_072 sky130_fd_sc_hs__nand2_4_123/a_27_74# sky130_fd_sc_hs__nand2_4
Xsky130_fd_sc_hs__nand2_2_86 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_2_88/Y sky130_fd_sc_hs__nand2_2_88/B
+ osc_072 sky130_fd_sc_hs__nand2_2_88/a_27_74# sky130_fd_sc_hs__nand2_2
Xsky130_fd_sc_hs__nand2_4_134 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_4_135/Y delay_con_msb[2]
+ osc_036 sky130_fd_sc_hs__nand2_4_135/a_27_74# sky130_fd_sc_hs__nand2_4
Xsky130_fd_sc_hs__nand2_2_97 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_2_97/Y sky130_fd_sc_hs__nand2_2_97/B
+ osc_036 sky130_fd_sc_hs__nand2_2_97/a_27_74# sky130_fd_sc_hs__nand2_2
Xsky130_fd_sc_hs__nand2_4_145 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_4_145/Y delay_con_msb[2]
+ osc_036 sky130_fd_sc_hs__nand2_4_145/a_27_74# sky130_fd_sc_hs__nand2_4
Xsky130_fd_sc_hs__nand2_4_156 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_4_157/Y delay_con_msb[1]
+ osc_036 sky130_fd_sc_hs__nand2_4_157/a_27_74# sky130_fd_sc_hs__nand2_4
Xsky130_fd_sc_hs__nand2_8_30 DVSS DVDD DVDD DVSS inj_out osc_072 osc_108 sky130_fd_sc_hs__nand2_8_31/a_27_74#
+ sky130_fd_sc_hs__nand2_8
Xsky130_fd_sc_hs__nand2_8_41 DVSS DVDD DVDD DVSS inj_out osc_072 osc_108 sky130_fd_sc_hs__nand2_8_41/a_27_74#
+ sky130_fd_sc_hs__nand2_8
Xsky130_fd_sc_hs__einvp_2_14 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_8_7/A sky130_fd_sc_hs__inv_4_17/Y
+ pi1_r[1] sky130_fd_sc_hs__einvp_2_15/a_263_323# sky130_fd_sc_hs__einvp_2_15/a_36_74#
+ sky130_fd_sc_hs__einvp_2_15/a_27_368# sky130_fd_sc_hs__einvp_2
Xsky130_fd_sc_hs__inv_4_20 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_21/Y osc_000
+ sky130_fd_sc_hs__inv_4
Xsky130_fd_sc_hs__inv_4_31 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_31/Y delay_con_lsb[4]
+ sky130_fd_sc_hs__inv_4
Xsky130_fd_sc_hs__einvp_2_8 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_8_5/A sky130_fd_sc_hs__inv_4_11/Y
+ pi4_l[1] sky130_fd_sc_hs__einvp_2_9/a_263_323# sky130_fd_sc_hs__einvp_2_9/a_36_74#
+ sky130_fd_sc_hs__einvp_2_9/a_27_368# sky130_fd_sc_hs__einvp_2
Xsky130_fd_sc_hs__einvp_8_13 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_8_7/A pi1_r[3]
+ sky130_fd_sc_hs__inv_4_17/Y sky130_fd_sc_hs__einvp_8_15/a_802_323# sky130_fd_sc_hs__einvp_8_15/a_27_74#
+ sky130_fd_sc_hs__einvp_8_15/a_27_368# sky130_fd_sc_hs__einvp_8
Xsky130_fd_sc_hs__nand2_2_10 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_2_12/Y sky130_fd_sc_hs__nand2_2_9/B
+ osc_000 sky130_fd_sc_hs__nand2_2_12/a_27_74# sky130_fd_sc_hs__nand2_2
Xsky130_fd_sc_hs__nand2_2_21 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_2_21/Y sky130_fd_sc_hs__nand2_2_7/B
+ osc_144 sky130_fd_sc_hs__nand2_2_21/a_27_74# sky130_fd_sc_hs__nand2_2
Xsky130_fd_sc_hs__nand2_2_32 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_2_33/Y sky130_fd_sc_hs__nand2_2_35/B
+ osc_000 sky130_fd_sc_hs__nand2_2_33/a_27_74# sky130_fd_sc_hs__nand2_2
Xsky130_fd_sc_hs__nand2_2_43 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_2_43/Y sky130_fd_sc_hs__nand2_2_43/B
+ osc_108 sky130_fd_sc_hs__nand2_2_43/a_27_74# sky130_fd_sc_hs__nand2_2
Xsky130_fd_sc_hs__nand2_2_54 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_2_55/Y sky130_fd_sc_hs__nand2_2_85/B
+ osc_072 sky130_fd_sc_hs__nand2_2_55/a_27_74# sky130_fd_sc_hs__nand2_2
Xsky130_fd_sc_hs__nand2_2_65 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_2_65/Y sky130_fd_sc_hs__nand2_2_65/B
+ osc_144 sky130_fd_sc_hs__nand2_2_65/a_27_74# sky130_fd_sc_hs__nand2_2
Xsky130_fd_sc_hs__nand2_4_102 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_4_102/Y delay_con_msb[0]
+ osc_072 sky130_fd_sc_hs__nand2_4_102/a_27_74# sky130_fd_sc_hs__nand2_4
Xsky130_fd_sc_hs__nand2_4_113 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_4_113/Y delay_con_msb[2]
+ osc_072 sky130_fd_sc_hs__nand2_4_113/a_27_74# sky130_fd_sc_hs__nand2_4
Xsky130_fd_sc_hs__nand2_2_76 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_2_79/Y sky130_fd_sc_hs__nand2_2_79/B
+ osc_072 sky130_fd_sc_hs__nand2_2_79/a_27_74# sky130_fd_sc_hs__nand2_2
Xsky130_fd_sc_hs__nand2_4_124 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_4_125/Y delay_con_msb[1]
+ osc_036 sky130_fd_sc_hs__nand2_4_125/a_27_74# sky130_fd_sc_hs__nand2_4
Xsky130_fd_sc_hs__nand2_2_87 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_2_89/Y sky130_fd_sc_hs__nand2_2_97/B
+ osc_036 sky130_fd_sc_hs__nand2_2_89/a_27_74# sky130_fd_sc_hs__nand2_2
Xsky130_fd_sc_hs__nand2_4_135 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_4_135/Y delay_con_msb[2]
+ osc_036 sky130_fd_sc_hs__nand2_4_135/a_27_74# sky130_fd_sc_hs__nand2_4
Xsky130_fd_sc_hs__nand2_4_146 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_4_147/Y delay_con_msb[0]
+ osc_036 sky130_fd_sc_hs__nand2_4_147/a_27_74# sky130_fd_sc_hs__nand2_4
Xsky130_fd_sc_hs__nand2_2_98 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_2_99/Y sky130_fd_sc_hs__nand2_2_99/B
+ osc_036 sky130_fd_sc_hs__nand2_2_99/a_27_74# sky130_fd_sc_hs__nand2_2
Xsky130_fd_sc_hs__nand2_4_157 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_4_157/Y delay_con_msb[1]
+ osc_036 sky130_fd_sc_hs__nand2_4_157/a_27_74# sky130_fd_sc_hs__nand2_4
Xsky130_fd_sc_hs__a21oi_1_0 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_31/Y sky130_fd_sc_hs__nand2_2_7/B
+ con_perb_4[0] sky130_fd_sc_hs__inv_4_29/Y sky130_fd_sc_hs__a21oi_1_1/a_117_74# sky130_fd_sc_hs__a21oi_1_1/a_29_368#
+ sky130_fd_sc_hs__a21oi_1
Xsky130_fd_sc_hs__nand2_8_20 DVSS DVDD DVDD DVSS inj_out osc_072 osc_108 sky130_fd_sc_hs__nand2_8_21/a_27_74#
+ sky130_fd_sc_hs__nand2_8
Xsky130_fd_sc_hs__nand2_8_31 DVSS DVDD DVDD DVSS inj_out osc_072 osc_108 sky130_fd_sc_hs__nand2_8_31/a_27_74#
+ sky130_fd_sc_hs__nand2_8
Xsky130_fd_sc_hs__nand2_8_42 DVSS DVDD DVDD DVSS osc_hold osc_036 osc_072 sky130_fd_sc_hs__nand2_8_43/a_27_74#
+ sky130_fd_sc_hs__nand2_8
Xsky130_fd_sc_hs__einvp_2_15 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_8_7/A sky130_fd_sc_hs__inv_4_17/Y
+ pi1_r[1] sky130_fd_sc_hs__einvp_2_15/a_263_323# sky130_fd_sc_hs__einvp_2_15/a_36_74#
+ sky130_fd_sc_hs__einvp_2_15/a_27_368# sky130_fd_sc_hs__einvp_2
Xsky130_fd_sc_hs__inv_4_10 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_11/Y osc_108
+ sky130_fd_sc_hs__inv_4
Xsky130_fd_sc_hs__inv_4_21 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_21/Y osc_000
+ sky130_fd_sc_hs__inv_4
Xsky130_fd_sc_hs__inv_4_32 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_33/Y delay_con_lsb[0]
+ sky130_fd_sc_hs__inv_4
Xsky130_fd_sc_hs__einvp_2_9 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_8_5/A sky130_fd_sc_hs__inv_4_11/Y
+ pi4_l[1] sky130_fd_sc_hs__einvp_2_9/a_263_323# sky130_fd_sc_hs__einvp_2_9/a_36_74#
+ sky130_fd_sc_hs__einvp_2_9/a_27_368# sky130_fd_sc_hs__einvp_2
Xsky130_fd_sc_hs__einvp_8_14 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_8_7/A pi1_l[3]
+ sky130_fd_sc_hs__inv_4_15/Y sky130_fd_sc_hs__einvp_8_14/a_802_323# sky130_fd_sc_hs__einvp_8_14/a_27_74#
+ sky130_fd_sc_hs__einvp_8_14/a_27_368# sky130_fd_sc_hs__einvp_8
Xsky130_fd_sc_hs__nand2_2_11 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_2_13/Y sky130_fd_sc_hs__nand2_2_5/B
+ osc_000 sky130_fd_sc_hs__nand2_2_13/a_27_74# sky130_fd_sc_hs__nand2_2
Xsky130_fd_sc_hs__nand2_2_22 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_2_23/Y sky130_fd_sc_hs__nand2_2_57/B
+ osc_144 sky130_fd_sc_hs__nand2_2_23/a_27_74# sky130_fd_sc_hs__nand2_2
Xsky130_fd_sc_hs__nand2_2_33 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_2_33/Y sky130_fd_sc_hs__nand2_2_35/B
+ osc_000 sky130_fd_sc_hs__nand2_2_33/a_27_74# sky130_fd_sc_hs__nand2_2
Xsky130_fd_sc_hs__nand2_2_44 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_2_45/Y sky130_fd_sc_hs__nand2_2_45/B
+ osc_108 sky130_fd_sc_hs__nand2_2_45/a_27_74# sky130_fd_sc_hs__nand2_2
Xsky130_fd_sc_hs__nand2_2_55 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_2_55/Y sky130_fd_sc_hs__nand2_2_85/B
+ osc_072 sky130_fd_sc_hs__nand2_2_55/a_27_74# sky130_fd_sc_hs__nand2_2
Xsky130_fd_sc_hs__nand2_2_66 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_2_67/Y sky130_fd_sc_hs__nand2_2_79/B
+ osc_072 sky130_fd_sc_hs__nand2_2_67/a_27_74# sky130_fd_sc_hs__nand2_2
Xsky130_fd_sc_hs__nand2_4_103 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_4_103/Y delay_con_msb[0]
+ osc_072 sky130_fd_sc_hs__nand2_4_103/a_27_74# sky130_fd_sc_hs__nand2_4
Xsky130_fd_sc_hs__nand2_4_114 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_4_115/Y delay_con_msb[2]
+ osc_072 sky130_fd_sc_hs__nand2_4_115/a_27_74# sky130_fd_sc_hs__nand2_4
Xsky130_fd_sc_hs__nand2_2_77 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_2_77/Y sky130_fd_sc_hs__nand2_2_79/B
+ osc_072 sky130_fd_sc_hs__nand2_2_77/a_27_74# sky130_fd_sc_hs__nand2_2
Xsky130_fd_sc_hs__nand2_4_125 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_4_125/Y delay_con_msb[1]
+ osc_036 sky130_fd_sc_hs__nand2_4_125/a_27_74# sky130_fd_sc_hs__nand2_4
Xsky130_fd_sc_hs__nand2_2_88 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_2_88/Y sky130_fd_sc_hs__nand2_2_88/B
+ osc_072 sky130_fd_sc_hs__nand2_2_88/a_27_74# sky130_fd_sc_hs__nand2_2
Xsky130_fd_sc_hs__nand2_4_136 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_4_137/Y delay_con_msb[2]
+ osc_036 sky130_fd_sc_hs__nand2_4_137/a_27_74# sky130_fd_sc_hs__nand2_4
Xsky130_fd_sc_hs__nand2_4_147 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_4_147/Y delay_con_msb[0]
+ osc_036 sky130_fd_sc_hs__nand2_4_147/a_27_74# sky130_fd_sc_hs__nand2_4
Xsky130_fd_sc_hs__nand2_2_99 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_2_99/Y sky130_fd_sc_hs__nand2_2_99/B
+ osc_036 sky130_fd_sc_hs__nand2_2_99/a_27_74# sky130_fd_sc_hs__nand2_2
Xsky130_fd_sc_hs__nand2_4_158 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_4_159/Y delay_con_msb[3]
+ osc_036 sky130_fd_sc_hs__nand2_4_159/a_27_74# sky130_fd_sc_hs__nand2_4
Xsky130_fd_sc_hs__a21oi_1_1 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_31/Y sky130_fd_sc_hs__nand2_2_7/B
+ con_perb_4[0] sky130_fd_sc_hs__inv_4_29/Y sky130_fd_sc_hs__a21oi_1_1/a_117_74# sky130_fd_sc_hs__a21oi_1_1/a_29_368#
+ sky130_fd_sc_hs__a21oi_1
Xsky130_fd_sc_hs__inv_16_0 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_16_1/Y sky130_fd_sc_hs__inv_16_9/A
+ sky130_fd_sc_hs__inv_16
Xsky130_fd_sc_hs__nand2_8_10 DVSS DVDD DVDD DVSS inj_out osc_072 osc_108 sky130_fd_sc_hs__nand2_8_11/a_27_74#
+ sky130_fd_sc_hs__nand2_8
Xsky130_fd_sc_hs__nand2_8_21 DVSS DVDD DVDD DVSS inj_out osc_072 osc_108 sky130_fd_sc_hs__nand2_8_21/a_27_74#
+ sky130_fd_sc_hs__nand2_8
Xsky130_fd_sc_hs__nand2_8_32 DVSS DVDD DVDD DVSS osc_hold osc_036 osc_072 sky130_fd_sc_hs__nand2_8_33/a_27_74#
+ sky130_fd_sc_hs__nand2_8
Xsky130_fd_sc_hs__nand2_8_43 DVSS DVDD DVDD DVSS osc_hold osc_036 osc_072 sky130_fd_sc_hs__nand2_8_43/a_27_74#
+ sky130_fd_sc_hs__nand2_8
Xsky130_fd_sc_hs__einvp_2_16 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_8_9/A sky130_fd_sc_hs__inv_4_19/Y
+ pi5_l[1] sky130_fd_sc_hs__einvp_2_17/a_263_323# sky130_fd_sc_hs__einvp_2_17/a_36_74#
+ sky130_fd_sc_hs__einvp_2_17/a_27_368# sky130_fd_sc_hs__einvp_2
Xsky130_fd_sc_hs__inv_4_11 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_11/Y osc_108
+ sky130_fd_sc_hs__inv_4
Xsky130_fd_sc_hs__inv_4_22 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_23/Y sky130_fd_sc_hs__inv_1_1/Y
+ sky130_fd_sc_hs__inv_4
Xsky130_fd_sc_hs__inv_4_33 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_33/Y delay_con_lsb[0]
+ sky130_fd_sc_hs__inv_4
Xsky130_fd_sc_hs__einvp_8_15 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_8_7/A pi1_r[3]
+ sky130_fd_sc_hs__inv_4_17/Y sky130_fd_sc_hs__einvp_8_15/a_802_323# sky130_fd_sc_hs__einvp_8_15/a_27_74#
+ sky130_fd_sc_hs__einvp_8_15/a_27_368# sky130_fd_sc_hs__einvp_8
Xsky130_fd_sc_hs__nand2_2_12 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_2_12/Y sky130_fd_sc_hs__nand2_2_9/B
+ osc_000 sky130_fd_sc_hs__nand2_2_12/a_27_74# sky130_fd_sc_hs__nand2_2
Xsky130_fd_sc_hs__nand2_2_23 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_2_23/Y sky130_fd_sc_hs__nand2_2_57/B
+ osc_144 sky130_fd_sc_hs__nand2_2_23/a_27_74# sky130_fd_sc_hs__nand2_2
Xsky130_fd_sc_hs__nand2_2_34 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_2_35/Y sky130_fd_sc_hs__nand2_2_35/B
+ osc_000 sky130_fd_sc_hs__nand2_2_35/a_27_74# sky130_fd_sc_hs__nand2_2
Xsky130_fd_sc_hs__nand2_2_45 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_2_45/Y sky130_fd_sc_hs__nand2_2_45/B
+ osc_108 sky130_fd_sc_hs__nand2_2_45/a_27_74# sky130_fd_sc_hs__nand2_2
Xsky130_fd_sc_hs__nand2_2_56 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_2_57/Y sky130_fd_sc_hs__nand2_2_57/B
+ osc_144 sky130_fd_sc_hs__nand2_2_57/a_27_74# sky130_fd_sc_hs__nand2_2
Xsky130_fd_sc_hs__nand2_2_67 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_2_67/Y sky130_fd_sc_hs__nand2_2_79/B
+ osc_072 sky130_fd_sc_hs__nand2_2_67/a_27_74# sky130_fd_sc_hs__nand2_2
Xsky130_fd_sc_hs__nand2_2_78 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_2_78/Y sky130_fd_sc_hs__nand2_2_79/B
+ osc_072 sky130_fd_sc_hs__nand2_2_78/a_27_74# sky130_fd_sc_hs__nand2_2
Xsky130_fd_sc_hs__nand2_4_104 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_4_106/Y delay_con_msb[1]
+ osc_072 sky130_fd_sc_hs__nand2_4_106/a_27_74# sky130_fd_sc_hs__nand2_4
Xsky130_fd_sc_hs__nand2_4_115 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_4_115/Y delay_con_msb[2]
+ osc_072 sky130_fd_sc_hs__nand2_4_115/a_27_74# sky130_fd_sc_hs__nand2_4
Xsky130_fd_sc_hs__nand2_4_126 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_4_127/Y delay_con_msb[0]
+ osc_036 sky130_fd_sc_hs__nand2_4_127/a_27_74# sky130_fd_sc_hs__nand2_4
Xsky130_fd_sc_hs__nand2_2_89 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_2_89/Y sky130_fd_sc_hs__nand2_2_97/B
+ osc_036 sky130_fd_sc_hs__nand2_2_89/a_27_74# sky130_fd_sc_hs__nand2_2
Xsky130_fd_sc_hs__nand2_4_137 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_4_137/Y delay_con_msb[2]
+ osc_036 sky130_fd_sc_hs__nand2_4_137/a_27_74# sky130_fd_sc_hs__nand2_4
Xsky130_fd_sc_hs__nand2_4_148 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_4_149/Y delay_con_msb[2]
+ osc_036 sky130_fd_sc_hs__nand2_4_149/a_27_74# sky130_fd_sc_hs__nand2_4
Xsky130_fd_sc_hs__nand2_4_159 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_4_159/Y delay_con_msb[3]
+ osc_036 sky130_fd_sc_hs__nand2_4_159/a_27_74# sky130_fd_sc_hs__nand2_4
Xsky130_fd_sc_hs__a21oi_1_2 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_33/Y sky130_fd_sc_hs__nand2_1_1/B
+ con_perb_4[0] sky130_fd_sc_hs__inv_4_29/Y sky130_fd_sc_hs__a21oi_1_3/a_117_74# sky130_fd_sc_hs__a21oi_1_3/a_29_368#
+ sky130_fd_sc_hs__a21oi_1
Xsky130_fd_sc_hs__inv_16_1 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_16_1/Y sky130_fd_sc_hs__inv_16_9/A
+ sky130_fd_sc_hs__inv_16
Xsky130_fd_sc_hs__nand2_8_11 DVSS DVDD DVDD DVSS inj_out osc_072 osc_108 sky130_fd_sc_hs__nand2_8_11/a_27_74#
+ sky130_fd_sc_hs__nand2_8
Xsky130_fd_sc_hs__nand2_8_22 DVSS DVDD DVDD DVSS osc_hold osc_036 osc_072 sky130_fd_sc_hs__nand2_8_23/a_27_74#
+ sky130_fd_sc_hs__nand2_8
Xsky130_fd_sc_hs__nand2_8_33 DVSS DVDD DVDD DVSS osc_hold osc_036 osc_072 sky130_fd_sc_hs__nand2_8_33/a_27_74#
+ sky130_fd_sc_hs__nand2_8
Xsky130_fd_sc_hs__nand2_8_44 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_8_9/B osc_108
+ osc_144 sky130_fd_sc_hs__nand2_8_45/a_27_74# sky130_fd_sc_hs__nand2_8
Xsky130_fd_sc_hs__einvp_2_17 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_8_9/A sky130_fd_sc_hs__inv_4_19/Y
+ pi5_l[1] sky130_fd_sc_hs__einvp_2_17/a_263_323# sky130_fd_sc_hs__einvp_2_17/a_36_74#
+ sky130_fd_sc_hs__einvp_2_17/a_27_368# sky130_fd_sc_hs__einvp_2
Xsky130_fd_sc_hs__inv_4_12 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_13/Y osc_144
+ sky130_fd_sc_hs__inv_4
Xsky130_fd_sc_hs__inv_4_23 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_23/Y sky130_fd_sc_hs__inv_1_1/Y
+ sky130_fd_sc_hs__inv_4
Xsky130_fd_sc_hs__inv_4_34 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_36/Y delay_con_lsb[1]
+ sky130_fd_sc_hs__inv_4
Xsky130_fd_sc_hs__einvp_8_16 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_8_9/A pi5_l[3]
+ sky130_fd_sc_hs__inv_4_19/Y sky130_fd_sc_hs__einvp_8_17/a_802_323# sky130_fd_sc_hs__einvp_8_17/a_27_74#
+ sky130_fd_sc_hs__einvp_8_17/a_27_368# sky130_fd_sc_hs__einvp_8
Xsky130_fd_sc_hs__nand2_2_13 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_2_13/Y sky130_fd_sc_hs__nand2_2_5/B
+ osc_000 sky130_fd_sc_hs__nand2_2_13/a_27_74# sky130_fd_sc_hs__nand2_2
Xsky130_fd_sc_hs__nand2_2_24 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_2_25/Y sky130_fd_sc_hs__nand2_2_9/B
+ osc_000 sky130_fd_sc_hs__nand2_2_25/a_27_74# sky130_fd_sc_hs__nand2_2
Xsky130_fd_sc_hs__nand2_2_35 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_2_35/Y sky130_fd_sc_hs__nand2_2_35/B
+ osc_000 sky130_fd_sc_hs__nand2_2_35/a_27_74# sky130_fd_sc_hs__nand2_2
Xsky130_fd_sc_hs__nand2_2_46 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_2_47/Y sky130_fd_sc_hs__nand2_2_65/B
+ osc_144 sky130_fd_sc_hs__nand2_2_47/a_27_74# sky130_fd_sc_hs__nand2_2
Xsky130_fd_sc_hs__nand2_2_57 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_2_57/Y sky130_fd_sc_hs__nand2_2_57/B
+ osc_144 sky130_fd_sc_hs__nand2_2_57/a_27_74# sky130_fd_sc_hs__nand2_2
Xsky130_fd_sc_hs__nand2_2_68 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_2_69/Y sky130_fd_sc_hs__nand2_2_85/B
+ osc_072 sky130_fd_sc_hs__nand2_2_69/a_27_74# sky130_fd_sc_hs__nand2_2
Xsky130_fd_sc_hs__nand2_4_105 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_4_107/Y delay_con_msb[1]
+ osc_108 sky130_fd_sc_hs__nand2_4_107/a_27_74# sky130_fd_sc_hs__nand2_4
Xsky130_fd_sc_hs__nand2_4_116 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_4_117/Y delay_con_msb[2]
+ osc_072 sky130_fd_sc_hs__nand2_4_117/a_27_74# sky130_fd_sc_hs__nand2_4
Xsky130_fd_sc_hs__nand2_2_79 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_2_79/Y sky130_fd_sc_hs__nand2_2_79/B
+ osc_072 sky130_fd_sc_hs__nand2_2_79/a_27_74# sky130_fd_sc_hs__nand2_2
Xsky130_fd_sc_hs__nand2_4_127 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_4_127/Y delay_con_msb[0]
+ osc_036 sky130_fd_sc_hs__nand2_4_127/a_27_74# sky130_fd_sc_hs__nand2_4
Xsky130_fd_sc_hs__nand2_4_138 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_4_139/Y delay_con_msb[3]
+ osc_036 sky130_fd_sc_hs__nand2_4_139/a_27_74# sky130_fd_sc_hs__nand2_4
Xsky130_fd_sc_hs__nand2_4_149 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_4_149/Y delay_con_msb[2]
+ osc_036 sky130_fd_sc_hs__nand2_4_149/a_27_74# sky130_fd_sc_hs__nand2_4
Xsky130_fd_sc_hs__a21oi_1_3 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_33/Y sky130_fd_sc_hs__nand2_1_1/B
+ con_perb_4[0] sky130_fd_sc_hs__inv_4_29/Y sky130_fd_sc_hs__a21oi_1_3/a_117_74# sky130_fd_sc_hs__a21oi_1_3/a_29_368#
+ sky130_fd_sc_hs__a21oi_1
Xsky130_fd_sc_hs__inv_16_2 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_16_3/Y sky130_fd_sc_hs__inv_16_9/A
+ sky130_fd_sc_hs__inv_16
Xsky130_fd_sc_hs__nand2_8_12 DVSS DVDD DVDD DVSS osc_hold osc_036 osc_072 sky130_fd_sc_hs__nand2_8_13/a_27_74#
+ sky130_fd_sc_hs__nand2_8
Xsky130_fd_sc_hs__nand2_8_23 DVSS DVDD DVDD DVSS osc_hold osc_036 osc_072 sky130_fd_sc_hs__nand2_8_23/a_27_74#
+ sky130_fd_sc_hs__nand2_8
Xsky130_fd_sc_hs__nand2_8_34 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_8_9/B osc_108
+ osc_144 sky130_fd_sc_hs__nand2_8_35/a_27_74# sky130_fd_sc_hs__nand2_8
Xsky130_fd_sc_hs__nand2_8_45 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_8_9/B osc_108
+ osc_144 sky130_fd_sc_hs__nand2_8_45/a_27_74# sky130_fd_sc_hs__nand2_8
Xsky130_fd_sc_hs__einvp_2_18 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_8_9/A sky130_fd_sc_hs__inv_4_21/Y
+ pi5_r[1] sky130_fd_sc_hs__einvp_2_19/a_263_323# sky130_fd_sc_hs__einvp_2_19/a_36_74#
+ sky130_fd_sc_hs__einvp_2_19/a_27_368# sky130_fd_sc_hs__einvp_2
Xsky130_fd_sc_hs__inv_4_13 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_13/Y osc_144
+ sky130_fd_sc_hs__inv_4
Xsky130_fd_sc_hs__inv_4_24 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_25/Y sky130_fd_sc_hs__inv_1_7/Y
+ sky130_fd_sc_hs__inv_4
Xsky130_fd_sc_hs__inv_4_35 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_37/Y delay_con_lsb[2]
+ sky130_fd_sc_hs__inv_4
Xsky130_fd_sc_hs__einvp_8_17 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_8_9/A pi5_l[3]
+ sky130_fd_sc_hs__inv_4_19/Y sky130_fd_sc_hs__einvp_8_17/a_802_323# sky130_fd_sc_hs__einvp_8_17/a_27_74#
+ sky130_fd_sc_hs__einvp_8_17/a_27_368# sky130_fd_sc_hs__einvp_8
Xsky130_fd_sc_hs__nand2_2_14 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_2_15/Y sky130_fd_sc_hs__nand2_2_7/B
+ osc_144 sky130_fd_sc_hs__nand2_2_15/a_27_74# sky130_fd_sc_hs__nand2_2
Xsky130_fd_sc_hs__nand2_2_25 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_2_25/Y sky130_fd_sc_hs__nand2_2_9/B
+ osc_000 sky130_fd_sc_hs__nand2_2_25/a_27_74# sky130_fd_sc_hs__nand2_2
Xsky130_fd_sc_hs__nand2_2_36 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_2_37/Y sky130_fd_sc_hs__nand2_2_37/B
+ osc_000 sky130_fd_sc_hs__nand2_2_37/a_27_74# sky130_fd_sc_hs__nand2_2
Xsky130_fd_sc_hs__nand2_2_47 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_2_47/Y sky130_fd_sc_hs__nand2_2_65/B
+ osc_144 sky130_fd_sc_hs__nand2_2_47/a_27_74# sky130_fd_sc_hs__nand2_2
Xsky130_fd_sc_hs__nand2_2_58 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_2_59/Y sky130_fd_sc_hs__nand2_2_61/B
+ osc_108 sky130_fd_sc_hs__nand2_2_59/a_27_74# sky130_fd_sc_hs__nand2_2
Xsky130_fd_sc_hs__nand2_2_69 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_2_69/Y sky130_fd_sc_hs__nand2_2_85/B
+ osc_072 sky130_fd_sc_hs__nand2_2_69/a_27_74# sky130_fd_sc_hs__nand2_2
Xsky130_fd_sc_hs__nand2_4_106 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_4_106/Y delay_con_msb[1]
+ osc_072 sky130_fd_sc_hs__nand2_4_106/a_27_74# sky130_fd_sc_hs__nand2_4
Xsky130_fd_sc_hs__nand2_4_117 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_4_117/Y delay_con_msb[2]
+ osc_072 sky130_fd_sc_hs__nand2_4_117/a_27_74# sky130_fd_sc_hs__nand2_4
Xsky130_fd_sc_hs__nand2_4_128 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_4_129/Y delay_con_msb[3]
+ osc_072 sky130_fd_sc_hs__nand2_4_129/a_27_74# sky130_fd_sc_hs__nand2_4
Xsky130_fd_sc_hs__nand2_4_139 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_4_139/Y delay_con_msb[3]
+ osc_036 sky130_fd_sc_hs__nand2_4_139/a_27_74# sky130_fd_sc_hs__nand2_4
Xsky130_fd_sc_hs__a21oi_1_4 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_31/Y sky130_fd_sc_hs__nand2_2_5/B
+ con_perb_5[0] sky130_fd_sc_hs__inv_4_29/Y sky130_fd_sc_hs__a21oi_1_5/a_117_74# sky130_fd_sc_hs__a21oi_1_5/a_29_368#
+ sky130_fd_sc_hs__a21oi_1
Xsky130_fd_sc_hs__inv_16_3 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_16_3/Y sky130_fd_sc_hs__inv_16_9/A
+ sky130_fd_sc_hs__inv_16
Xsky130_fd_sc_hs__nand2_8_13 DVSS DVDD DVDD DVSS osc_hold osc_036 osc_072 sky130_fd_sc_hs__nand2_8_13/a_27_74#
+ sky130_fd_sc_hs__nand2_8
Xsky130_fd_sc_hs__nand2_8_24 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_8_9/B osc_108
+ osc_144 sky130_fd_sc_hs__nand2_8_25/a_27_74# sky130_fd_sc_hs__nand2_8
Xsky130_fd_sc_hs__nand2_8_35 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_8_9/B osc_108
+ osc_144 sky130_fd_sc_hs__nand2_8_35/a_27_74# sky130_fd_sc_hs__nand2_8
Xsky130_fd_sc_hs__nand2_8_46 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_8_9/B osc_000
+ osc_036 sky130_fd_sc_hs__nand2_8_47/a_27_74# sky130_fd_sc_hs__nand2_8
Xsky130_fd_sc_hs__einvp_2_19 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_8_9/A sky130_fd_sc_hs__inv_4_21/Y
+ pi5_r[1] sky130_fd_sc_hs__einvp_2_19/a_263_323# sky130_fd_sc_hs__einvp_2_19/a_36_74#
+ sky130_fd_sc_hs__einvp_2_19/a_27_368# sky130_fd_sc_hs__einvp_2
Xsky130_fd_sc_hs__inv_4_14 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_15/Y osc_000
+ sky130_fd_sc_hs__inv_4
Xsky130_fd_sc_hs__inv_4_25 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_25/Y sky130_fd_sc_hs__inv_1_7/Y
+ sky130_fd_sc_hs__inv_4
Xsky130_fd_sc_hs__inv_4_36 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_36/Y delay_con_lsb[1]
+ sky130_fd_sc_hs__inv_4
Xsky130_fd_sc_hs__einvp_8_18 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_8_9/A pi5_r[3]
+ sky130_fd_sc_hs__inv_4_21/Y sky130_fd_sc_hs__einvp_8_19/a_802_323# sky130_fd_sc_hs__einvp_8_19/a_27_74#
+ sky130_fd_sc_hs__einvp_8_19/a_27_368# sky130_fd_sc_hs__einvp_8
Xsky130_fd_sc_hs__nand2_2_15 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_2_15/Y sky130_fd_sc_hs__nand2_2_7/B
+ osc_144 sky130_fd_sc_hs__nand2_2_15/a_27_74# sky130_fd_sc_hs__nand2_2
Xsky130_fd_sc_hs__nand2_2_26 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_2_27/Y sky130_fd_sc_hs__nand2_2_43/B
+ osc_108 sky130_fd_sc_hs__nand2_2_27/a_27_74# sky130_fd_sc_hs__nand2_2
Xsky130_fd_sc_hs__nand2_2_37 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_2_37/Y sky130_fd_sc_hs__nand2_2_37/B
+ osc_000 sky130_fd_sc_hs__nand2_2_37/a_27_74# sky130_fd_sc_hs__nand2_2
Xsky130_fd_sc_hs__nand2_2_48 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_2_49/Y sky130_fd_sc_hs__nand2_2_65/B
+ osc_144 sky130_fd_sc_hs__nand2_2_49/a_27_74# sky130_fd_sc_hs__nand2_2
Xsky130_fd_sc_hs__nand2_2_59 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_2_59/Y sky130_fd_sc_hs__nand2_2_61/B
+ osc_108 sky130_fd_sc_hs__nand2_2_59/a_27_74# sky130_fd_sc_hs__nand2_2
Xsky130_fd_sc_hs__nand2_4_107 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_4_107/Y delay_con_msb[1]
+ osc_108 sky130_fd_sc_hs__nand2_4_107/a_27_74# sky130_fd_sc_hs__nand2_4
Xsky130_fd_sc_hs__nand2_4_118 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_4_119/Y delay_con_msb[3]
+ osc_072 sky130_fd_sc_hs__nand2_4_119/a_27_74# sky130_fd_sc_hs__nand2_4
Xsky130_fd_sc_hs__nand2_4_129 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_4_129/Y delay_con_msb[3]
+ osc_072 sky130_fd_sc_hs__nand2_4_129/a_27_74# sky130_fd_sc_hs__nand2_4
Xsky130_fd_sc_hs__dlygate4sd3_1_0 DVSS DVDD DVSS DVDD sky130_fd_sc_hs__dlygate4sd3_1_1/A
+ sky130_fd_sc_hs__dlygate4sd3_1_1/X sky130_fd_sc_hs__dlygate4sd3_1_1/a_405_138# sky130_fd_sc_hs__dlygate4sd3_1_1/a_28_74#
+ sky130_fd_sc_hs__dlygate4sd3_1_1/a_289_74# sky130_fd_sc_hs__dlygate4sd3_1
Xsky130_fd_sc_hs__a21oi_1_5 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_31/Y sky130_fd_sc_hs__nand2_2_5/B
+ con_perb_5[0] sky130_fd_sc_hs__inv_4_29/Y sky130_fd_sc_hs__a21oi_1_5/a_117_74# sky130_fd_sc_hs__a21oi_1_5/a_29_368#
+ sky130_fd_sc_hs__a21oi_1
Xsky130_fd_sc_hs__inv_16_4 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_16_5/Y sky130_fd_sc_hs__inv_16_9/A
+ sky130_fd_sc_hs__inv_16
Xsky130_fd_sc_hs__nand2_8_14 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_8_9/B osc_108
+ osc_144 sky130_fd_sc_hs__nand2_8_15/a_27_74# sky130_fd_sc_hs__nand2_8
Xsky130_fd_sc_hs__nand2_8_25 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_8_9/B osc_108
+ osc_144 sky130_fd_sc_hs__nand2_8_25/a_27_74# sky130_fd_sc_hs__nand2_8
Xsky130_fd_sc_hs__nand2_8_36 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_8_9/B osc_000
+ osc_036 sky130_fd_sc_hs__nand2_8_37/a_27_74# sky130_fd_sc_hs__nand2_8
Xsky130_fd_sc_hs__nand2_8_47 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_8_9/B osc_000
+ osc_036 sky130_fd_sc_hs__nand2_8_47/a_27_74# sky130_fd_sc_hs__nand2_8
Xsky130_fd_sc_hs__and4_2_0 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_16_5/Y sky130_fd_sc_hs__inv_16_9/Y
+ sky130_fd_sc_hs__inv_16_1/Y sky130_fd_sc_hs__inv_16_3/Y sky130_fd_sc_hs__and4_2_1/X
+ sky130_fd_sc_hs__and4_2_1/a_335_74# sky130_fd_sc_hs__and4_2_1/a_143_74# sky130_fd_sc_hs__and4_2_1/a_221_74#
+ sky130_fd_sc_hs__and4_2_1/a_56_74# sky130_fd_sc_hs__and4_2
Xsky130_fd_sc_hs__inv_4_15 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_15/Y osc_000
+ sky130_fd_sc_hs__inv_4
Xsky130_fd_sc_hs__inv_4_26 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_27/Y sky130_fd_sc_hs__inv_1_9/Y
+ sky130_fd_sc_hs__inv_4
Xsky130_fd_sc_hs__inv_4_37 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_37/Y delay_con_lsb[2]
+ sky130_fd_sc_hs__inv_4
Xsky130_fd_sc_hs__einvp_8_19 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_8_9/A pi5_r[3]
+ sky130_fd_sc_hs__inv_4_21/Y sky130_fd_sc_hs__einvp_8_19/a_802_323# sky130_fd_sc_hs__einvp_8_19/a_27_74#
+ sky130_fd_sc_hs__einvp_8_19/a_27_368# sky130_fd_sc_hs__einvp_8
Xsky130_fd_sc_hs__nand2_1_0 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_1_1/B sky130_fd_sc_hs__nand2_1_1/Y
+ osc_144 sky130_fd_sc_hs__nand2_1_1/a_117_74# sky130_fd_sc_hs__nand2_1
Xsky130_fd_sc_hs__nand2_2_16 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_2_17/Y sky130_fd_sc_hs__nand2_2_5/B
+ osc_000 sky130_fd_sc_hs__nand2_2_17/a_27_74# sky130_fd_sc_hs__nand2_2
Xsky130_fd_sc_hs__nand2_2_27 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_2_27/Y sky130_fd_sc_hs__nand2_2_43/B
+ osc_108 sky130_fd_sc_hs__nand2_2_27/a_27_74# sky130_fd_sc_hs__nand2_2
Xsky130_fd_sc_hs__nand2_2_38 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_2_39/Y sky130_fd_sc_hs__nand2_2_61/B
+ osc_108 sky130_fd_sc_hs__nand2_2_39/a_27_74# sky130_fd_sc_hs__nand2_2
Xsky130_fd_sc_hs__nand2_2_49 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_2_49/Y sky130_fd_sc_hs__nand2_2_65/B
+ osc_144 sky130_fd_sc_hs__nand2_2_49/a_27_74# sky130_fd_sc_hs__nand2_2
Xsky130_fd_sc_hs__nand2_4_108 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_4_110/Y delay_con_msb[1]
+ osc_072 sky130_fd_sc_hs__nand2_4_110/a_27_74# sky130_fd_sc_hs__nand2_4
Xsky130_fd_sc_hs__nand2_4_119 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_4_119/Y delay_con_msb[3]
+ osc_072 sky130_fd_sc_hs__nand2_4_119/a_27_74# sky130_fd_sc_hs__nand2_4
Xsky130_fd_sc_hs__dlygate4sd3_1_1 DVSS DVDD DVSS DVDD sky130_fd_sc_hs__dlygate4sd3_1_1/A
+ sky130_fd_sc_hs__dlygate4sd3_1_1/X sky130_fd_sc_hs__dlygate4sd3_1_1/a_405_138# sky130_fd_sc_hs__dlygate4sd3_1_1/a_28_74#
+ sky130_fd_sc_hs__dlygate4sd3_1_1/a_289_74# sky130_fd_sc_hs__dlygate4sd3_1
Xsky130_fd_sc_hs__a21oi_1_6 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_39/Y sky130_fd_sc_hs__nand2_2_9/B
+ con_perb_5[3] sky130_fd_sc_hs__inv_4_29/Y sky130_fd_sc_hs__a21oi_1_7/a_117_74# sky130_fd_sc_hs__a21oi_1_7/a_29_368#
+ sky130_fd_sc_hs__a21oi_1
Xsky130_fd_sc_hs__inv_16_5 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_16_5/Y sky130_fd_sc_hs__inv_16_9/A
+ sky130_fd_sc_hs__inv_16
Xsky130_fd_sc_hs__nand2_8_15 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_8_9/B osc_108
+ osc_144 sky130_fd_sc_hs__nand2_8_15/a_27_74# sky130_fd_sc_hs__nand2_8
Xsky130_fd_sc_hs__nand2_8_26 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_8_9/B osc_000
+ osc_036 sky130_fd_sc_hs__nand2_8_27/a_27_74# sky130_fd_sc_hs__nand2_8
Xsky130_fd_sc_hs__nand2_8_37 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_8_9/B osc_000
+ osc_036 sky130_fd_sc_hs__nand2_8_37/a_27_74# sky130_fd_sc_hs__nand2_8
Xsky130_fd_sc_hs__nand2_8_48 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_8_9/B osc_144
+ osc_000 sky130_fd_sc_hs__nand2_8_49/a_27_74# sky130_fd_sc_hs__nand2_8
Xsky130_fd_sc_hs__inv_1_0 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_1_1/Y sky130_fd_sc_hs__inv_4_1/Y
+ sky130_fd_sc_hs__inv_1
Xsky130_fd_sc_hs__and4_2_1 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_16_5/Y sky130_fd_sc_hs__inv_16_9/Y
+ sky130_fd_sc_hs__inv_16_1/Y sky130_fd_sc_hs__inv_16_3/Y sky130_fd_sc_hs__and4_2_1/X
+ sky130_fd_sc_hs__and4_2_1/a_335_74# sky130_fd_sc_hs__and4_2_1/a_143_74# sky130_fd_sc_hs__and4_2_1/a_221_74#
+ sky130_fd_sc_hs__and4_2_1/a_56_74# sky130_fd_sc_hs__and4_2
Xsky130_fd_sc_hs__inv_4_16 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_17/Y osc_036
+ sky130_fd_sc_hs__inv_4
Xsky130_fd_sc_hs__inv_4_27 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_27/Y sky130_fd_sc_hs__inv_1_9/Y
+ sky130_fd_sc_hs__inv_4
Xsky130_fd_sc_hs__inv_4_38 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_39/Y delay_con_lsb[3]
+ sky130_fd_sc_hs__inv_4
Xsky130_fd_sc_hs__nand2_1_1 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_1_1/B sky130_fd_sc_hs__nand2_1_1/Y
+ osc_144 sky130_fd_sc_hs__nand2_1_1/a_117_74# sky130_fd_sc_hs__nand2_1
Xsky130_fd_sc_hs__nand2_2_17 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_2_17/Y sky130_fd_sc_hs__nand2_2_5/B
+ osc_000 sky130_fd_sc_hs__nand2_2_17/a_27_74# sky130_fd_sc_hs__nand2_2
Xsky130_fd_sc_hs__nand2_2_28 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_2_29/Y sky130_fd_sc_hs__nand2_2_43/B
+ osc_108 sky130_fd_sc_hs__nand2_2_29/a_27_74# sky130_fd_sc_hs__nand2_2
Xsky130_fd_sc_hs__nand2_2_39 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_2_39/Y sky130_fd_sc_hs__nand2_2_61/B
+ osc_108 sky130_fd_sc_hs__nand2_2_39/a_27_74# sky130_fd_sc_hs__nand2_2
Xsky130_fd_sc_hs__nand2_4_109 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_4_111/Y delay_con_msb[1]
+ osc_072 sky130_fd_sc_hs__nand2_4_111/a_27_74# sky130_fd_sc_hs__nand2_4
Xsky130_fd_sc_hs__dlygate4sd3_1_2 DVSS DVDD DVSS DVDD sky130_fd_sc_hs__dlygate4sd3_1_3/A
+ sky130_fd_sc_hs__dlygate4sd3_1_3/X sky130_fd_sc_hs__dlygate4sd3_1_3/a_405_138# sky130_fd_sc_hs__dlygate4sd3_1_3/a_28_74#
+ sky130_fd_sc_hs__dlygate4sd3_1_3/a_289_74# sky130_fd_sc_hs__dlygate4sd3_1
Xsky130_fd_sc_hs__a21oi_1_7 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_39/Y sky130_fd_sc_hs__nand2_2_9/B
+ con_perb_5[3] sky130_fd_sc_hs__inv_4_29/Y sky130_fd_sc_hs__a21oi_1_7/a_117_74# sky130_fd_sc_hs__a21oi_1_7/a_29_368#
+ sky130_fd_sc_hs__a21oi_1
Xsky130_fd_sc_hs__inv_16_6 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_16_7/Y sky130_fd_sc_hs__inv_4_23/Y
+ sky130_fd_sc_hs__inv_16
Xsky130_fd_sc_hs__nand2_8_16 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_8_9/B osc_000
+ osc_036 sky130_fd_sc_hs__nand2_8_17/a_27_74# sky130_fd_sc_hs__nand2_8
Xsky130_fd_sc_hs__nand2_8_27 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_8_9/B osc_000
+ osc_036 sky130_fd_sc_hs__nand2_8_27/a_27_74# sky130_fd_sc_hs__nand2_8
Xsky130_fd_sc_hs__nand2_8_38 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_8_9/B osc_144
+ osc_000 sky130_fd_sc_hs__nand2_8_39/a_27_74# sky130_fd_sc_hs__nand2_8
Xsky130_fd_sc_hs__nand2_8_49 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_8_9/B osc_144
+ osc_000 sky130_fd_sc_hs__nand2_8_49/a_27_74# sky130_fd_sc_hs__nand2_8
Xsky130_fd_sc_hs__inv_1_1 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_1_1/Y sky130_fd_sc_hs__inv_4_1/Y
+ sky130_fd_sc_hs__inv_1
Xsky130_fd_sc_hs__and4_2_2 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__and4_2_3/D sky130_fd_sc_hs__and4_2_3/C
+ sky130_fd_sc_hs__and4_2_3/B sky130_fd_sc_hs__and4_2_3/A sky130_fd_sc_hs__and4_2_3/X
+ sky130_fd_sc_hs__and4_2_3/a_335_74# sky130_fd_sc_hs__and4_2_3/a_143_74# sky130_fd_sc_hs__and4_2_3/a_221_74#
+ sky130_fd_sc_hs__and4_2_3/a_56_74# sky130_fd_sc_hs__and4_2
Xsky130_fd_sc_hs__inv_4_17 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_17/Y osc_036
+ sky130_fd_sc_hs__inv_4
Xsky130_fd_sc_hs__inv_4_28 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_29/Y ref_clk
+ sky130_fd_sc_hs__inv_4
Xsky130_fd_sc_hs__inv_4_39 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_39/Y delay_con_lsb[3]
+ sky130_fd_sc_hs__inv_4
Xsky130_fd_sc_hs__nand2_1_2 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_1_3/B sky130_fd_sc_hs__nand2_1_3/Y
+ osc_000 sky130_fd_sc_hs__nand2_1_3/a_117_74# sky130_fd_sc_hs__nand2_1
Xsky130_fd_sc_hs__nand3_4_0 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand3_4_3/C sky130_fd_sc_hs__and2_2_3/X
+ sky130_fd_sc_hs__and4_2_1/X sky130_fd_sc_hs__and2_2_1/A sky130_fd_sc_hs__nand3_4_1/a_456_82#
+ sky130_fd_sc_hs__nand3_4_1/a_27_82# sky130_fd_sc_hs__nand3_4
Xsky130_fd_sc_hs__nand2_2_18 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_2_19/Y sky130_fd_sc_hs__nand2_2_43/B
+ osc_108 sky130_fd_sc_hs__nand2_2_19/a_27_74# sky130_fd_sc_hs__nand2_2
Xsky130_fd_sc_hs__nand2_2_29 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_2_29/Y sky130_fd_sc_hs__nand2_2_43/B
+ osc_108 sky130_fd_sc_hs__nand2_2_29/a_27_74# sky130_fd_sc_hs__nand2_2
Xsky130_fd_sc_hs__dlygate4sd3_1_3 DVSS DVDD DVSS DVDD sky130_fd_sc_hs__dlygate4sd3_1_3/A
+ sky130_fd_sc_hs__dlygate4sd3_1_3/X sky130_fd_sc_hs__dlygate4sd3_1_3/a_405_138# sky130_fd_sc_hs__dlygate4sd3_1_3/a_28_74#
+ sky130_fd_sc_hs__dlygate4sd3_1_3/a_289_74# sky130_fd_sc_hs__dlygate4sd3_1
Xsky130_fd_sc_hs__a21oi_1_8 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_33/Y sky130_fd_sc_hs__nand2_1_3/B
+ con_perb_5[0] sky130_fd_sc_hs__inv_4_29/Y sky130_fd_sc_hs__a21oi_1_9/a_117_74# sky130_fd_sc_hs__a21oi_1_9/a_29_368#
+ sky130_fd_sc_hs__a21oi_1
Xsky130_fd_sc_hs__inv_16_7 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_16_7/Y sky130_fd_sc_hs__inv_4_23/Y
+ sky130_fd_sc_hs__inv_16
Xsky130_fd_sc_hs__clkbuf_1_0 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__clkbuf_1_1/A osc_hold
+ sky130_fd_sc_hs__clkbuf_1_1/a_27_74# sky130_fd_sc_hs__clkbuf_1
Xsky130_fd_sc_hs__nand2_8_17 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_8_9/B osc_000
+ osc_036 sky130_fd_sc_hs__nand2_8_17/a_27_74# sky130_fd_sc_hs__nand2_8
Xsky130_fd_sc_hs__nand2_8_28 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_8_9/B osc_144
+ osc_000 sky130_fd_sc_hs__nand2_8_29/a_27_74# sky130_fd_sc_hs__nand2_8
Xsky130_fd_sc_hs__nand2_8_39 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_8_9/B osc_144
+ osc_000 sky130_fd_sc_hs__nand2_8_39/a_27_74# sky130_fd_sc_hs__nand2_8
Xsky130_fd_sc_hs__inv_1_2 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_1_7/A sky130_fd_sc_hs__inv_1_5/A
+ sky130_fd_sc_hs__inv_1
Xsky130_fd_sc_hs__and4_2_3 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__and4_2_3/D sky130_fd_sc_hs__and4_2_3/C
+ sky130_fd_sc_hs__and4_2_3/B sky130_fd_sc_hs__and4_2_3/A sky130_fd_sc_hs__and4_2_3/X
+ sky130_fd_sc_hs__and4_2_3/a_335_74# sky130_fd_sc_hs__and4_2_3/a_143_74# sky130_fd_sc_hs__and4_2_3/a_221_74#
+ sky130_fd_sc_hs__and4_2_3/a_56_74# sky130_fd_sc_hs__and4_2
Xsky130_fd_sc_hs__inv_4_18 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_19/Y osc_144
+ sky130_fd_sc_hs__inv_4
Xsky130_fd_sc_hs__inv_4_29 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_29/Y ref_clk
+ sky130_fd_sc_hs__inv_4
Xsky130_fd_sc_hs__nand2_1_3 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_1_3/B sky130_fd_sc_hs__nand2_1_3/Y
+ osc_000 sky130_fd_sc_hs__nand2_1_3/a_117_74# sky130_fd_sc_hs__nand2_1
Xsky130_fd_sc_hs__a21oi_1_40 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_33/Y sky130_fd_sc_hs__nand2_1_9/B
+ con_perb_1[0] sky130_fd_sc_hs__inv_4_29/Y sky130_fd_sc_hs__a21oi_1_42/a_117_74#
+ sky130_fd_sc_hs__a21oi_1_42/a_29_368# sky130_fd_sc_hs__a21oi_1
Xsky130_fd_sc_hs__nand3_4_1 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand3_4_3/C sky130_fd_sc_hs__and2_2_3/X
+ sky130_fd_sc_hs__and4_2_1/X sky130_fd_sc_hs__and2_2_1/A sky130_fd_sc_hs__nand3_4_1/a_456_82#
+ sky130_fd_sc_hs__nand3_4_1/a_27_82# sky130_fd_sc_hs__nand3_4
Xsky130_fd_sc_hs__nand2_2_19 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_2_19/Y sky130_fd_sc_hs__nand2_2_43/B
+ osc_108 sky130_fd_sc_hs__nand2_2_19/a_27_74# sky130_fd_sc_hs__nand2_2
Xsky130_fd_sc_hs__dlygate4sd3_1_4 DVSS DVDD DVSS DVDD sky130_fd_sc_hs__dlygate4sd3_1_5/A
+ sky130_fd_sc_hs__dlygate4sd3_1_7/A sky130_fd_sc_hs__dlygate4sd3_1_5/a_405_138# sky130_fd_sc_hs__dlygate4sd3_1_5/a_28_74#
+ sky130_fd_sc_hs__dlygate4sd3_1_5/a_289_74# sky130_fd_sc_hs__dlygate4sd3_1
Xsky130_fd_sc_hs__a21oi_1_9 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_33/Y sky130_fd_sc_hs__nand2_1_3/B
+ con_perb_5[0] sky130_fd_sc_hs__inv_4_29/Y sky130_fd_sc_hs__a21oi_1_9/a_117_74# sky130_fd_sc_hs__a21oi_1_9/a_29_368#
+ sky130_fd_sc_hs__a21oi_1
Xsky130_fd_sc_hs__inv_16_8 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_16_9/Y sky130_fd_sc_hs__inv_16_9/A
+ sky130_fd_sc_hs__inv_16
Xsky130_fd_sc_hs__clkbuf_1_1 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__clkbuf_1_1/A osc_hold
+ sky130_fd_sc_hs__clkbuf_1_1/a_27_74# sky130_fd_sc_hs__clkbuf_1
Xsky130_fd_sc_hs__nand2_8_18 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_8_9/B osc_144
+ osc_000 sky130_fd_sc_hs__nand2_8_19/a_27_74# sky130_fd_sc_hs__nand2_8
Xsky130_fd_sc_hs__nand2_8_29 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_8_9/B osc_144
+ osc_000 sky130_fd_sc_hs__nand2_8_29/a_27_74# sky130_fd_sc_hs__nand2_8
Xsky130_fd_sc_hs__inv_1_3 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_1_7/A sky130_fd_sc_hs__inv_1_5/A
+ sky130_fd_sc_hs__inv_1
Xsky130_fd_sc_hs__and4_2_4 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__and4_2_5/D sky130_fd_sc_hs__and4_2_5/C
+ sky130_fd_sc_hs__and4_2_5/B sky130_fd_sc_hs__and4_2_5/A sky130_fd_sc_hs__inv_1_5/A
+ sky130_fd_sc_hs__and4_2_5/a_335_74# sky130_fd_sc_hs__and4_2_5/a_143_74# sky130_fd_sc_hs__and4_2_5/a_221_74#
+ sky130_fd_sc_hs__and4_2_5/a_56_74# sky130_fd_sc_hs__and4_2
Xsky130_fd_sc_hs__inv_4_19 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_19/Y osc_144
+ sky130_fd_sc_hs__inv_4
Xsky130_fd_sc_hs__nand2_1_4 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_1_5/B sky130_fd_sc_hs__nand2_1_5/Y
+ osc_108 sky130_fd_sc_hs__nand2_1_5/a_117_74# sky130_fd_sc_hs__nand2_1
Xsky130_fd_sc_hs__a21oi_1_30 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_37/Y sky130_fd_sc_hs__nand2_2_73/B
+ con_perb_3[2] sky130_fd_sc_hs__inv_4_29/Y sky130_fd_sc_hs__a21oi_1_32/a_117_74#
+ sky130_fd_sc_hs__a21oi_1_32/a_29_368# sky130_fd_sc_hs__a21oi_1
Xsky130_fd_sc_hs__a21oi_1_41 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_31/Y sky130_fd_sc_hs__nand2_2_97/B
+ con_perb_1[0] sky130_fd_sc_hs__inv_4_29/Y sky130_fd_sc_hs__a21oi_1_43/a_117_74#
+ sky130_fd_sc_hs__a21oi_1_43/a_29_368# sky130_fd_sc_hs__a21oi_1
Xsky130_fd_sc_hs__nand3_4_2 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand3_4_3/C sky130_fd_sc_hs__and2_2_3/X
+ sky130_fd_sc_hs__and4_2_1/X sky130_fd_sc_hs__and2_2_1/B sky130_fd_sc_hs__nand3_4_3/a_456_82#
+ sky130_fd_sc_hs__nand3_4_3/a_27_82# sky130_fd_sc_hs__nand3_4
Xsky130_fd_sc_hs__dlygate4sd3_1_5 DVSS DVDD DVSS DVDD sky130_fd_sc_hs__dlygate4sd3_1_5/A
+ sky130_fd_sc_hs__dlygate4sd3_1_7/A sky130_fd_sc_hs__dlygate4sd3_1_5/a_405_138# sky130_fd_sc_hs__dlygate4sd3_1_5/a_28_74#
+ sky130_fd_sc_hs__dlygate4sd3_1_5/a_289_74# sky130_fd_sc_hs__dlygate4sd3_1
Xsky130_fd_sc_hs__inv_16_9 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_16_9/Y sky130_fd_sc_hs__inv_16_9/A
+ sky130_fd_sc_hs__inv_16
Xsky130_fd_sc_hs__nand2_8_19 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_8_9/B osc_144
+ osc_000 sky130_fd_sc_hs__nand2_8_19/a_27_74# sky130_fd_sc_hs__nand2_8
Xsky130_fd_sc_hs__inv_1_4 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_1_9/A sky130_fd_sc_hs__inv_1_5/A
+ sky130_fd_sc_hs__inv_1
Xsky130_fd_sc_hs__and4_2_5 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__and4_2_5/D sky130_fd_sc_hs__and4_2_5/C
+ sky130_fd_sc_hs__and4_2_5/B sky130_fd_sc_hs__and4_2_5/A sky130_fd_sc_hs__inv_1_5/A
+ sky130_fd_sc_hs__and4_2_5/a_335_74# sky130_fd_sc_hs__and4_2_5/a_143_74# sky130_fd_sc_hs__and4_2_5/a_221_74#
+ sky130_fd_sc_hs__and4_2_5/a_56_74# sky130_fd_sc_hs__and4_2
Xsky130_fd_sc_hs__nand2_1_5 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_1_5/B sky130_fd_sc_hs__nand2_1_5/Y
+ osc_108 sky130_fd_sc_hs__nand2_1_5/a_117_74# sky130_fd_sc_hs__nand2_1
Xsky130_fd_sc_hs__a21oi_1_20 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_33/Y sky130_fd_sc_hs__nand2_1_5/B
+ con_perb_3[0] sky130_fd_sc_hs__inv_4_29/Y sky130_fd_sc_hs__a21oi_1_21/a_117_74#
+ sky130_fd_sc_hs__a21oi_1_21/a_29_368# sky130_fd_sc_hs__a21oi_1
Xsky130_fd_sc_hs__a21oi_1_31 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_39/Y sky130_fd_sc_hs__nand2_2_61/B
+ con_perb_3[3] sky130_fd_sc_hs__inv_4_29/Y sky130_fd_sc_hs__a21oi_1_33/a_117_74#
+ sky130_fd_sc_hs__a21oi_1_33/a_29_368# sky130_fd_sc_hs__a21oi_1
Xsky130_fd_sc_hs__a21oi_1_42 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_33/Y sky130_fd_sc_hs__nand2_1_9/B
+ con_perb_1[0] sky130_fd_sc_hs__inv_4_29/Y sky130_fd_sc_hs__a21oi_1_42/a_117_74#
+ sky130_fd_sc_hs__a21oi_1_42/a_29_368# sky130_fd_sc_hs__a21oi_1
Xsky130_fd_sc_hs__nand3_4_3 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand3_4_3/C sky130_fd_sc_hs__and2_2_3/X
+ sky130_fd_sc_hs__and4_2_1/X sky130_fd_sc_hs__and2_2_1/B sky130_fd_sc_hs__nand3_4_3/a_456_82#
+ sky130_fd_sc_hs__nand3_4_3/a_27_82# sky130_fd_sc_hs__nand3_4
Xsky130_fd_sc_hs__dlygate4sd3_1_6 DVSS DVDD DVSS DVDD sky130_fd_sc_hs__dlygate4sd3_1_7/A
+ sky130_fd_sc_hs__dlygate4sd3_1_7/X sky130_fd_sc_hs__dlygate4sd3_1_7/a_405_138# sky130_fd_sc_hs__dlygate4sd3_1_7/a_28_74#
+ sky130_fd_sc_hs__dlygate4sd3_1_7/a_289_74# sky130_fd_sc_hs__dlygate4sd3_1
Xsky130_fd_sc_hs__einvp_1_0 DVSS DVDD DVDD DVSS pi3_l[0] sky130_fd_sc_hs__inv_8_1/A
+ sky130_fd_sc_hs__inv_4_3/Y sky130_fd_sc_hs__einvp_1_1/a_44_549# sky130_fd_sc_hs__einvp_1_1/a_318_74#
+ sky130_fd_sc_hs__einvp_1_1/a_310_392# sky130_fd_sc_hs__einvp_1
Xsky130_fd_sc_hs__inv_1_5 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_1_9/A sky130_fd_sc_hs__inv_1_5/A
+ sky130_fd_sc_hs__inv_1
Xsky130_fd_sc_hs__nand2_1_6 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_1_7/B sky130_fd_sc_hs__nand2_1_7/Y
+ osc_072 sky130_fd_sc_hs__nand2_1_7/a_117_74# sky130_fd_sc_hs__nand2_1
Xsky130_fd_sc_hs__a21oi_1_10 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_37/Y sky130_fd_sc_hs__nand2_2_35/B
+ con_perb_5[2] sky130_fd_sc_hs__inv_4_29/Y sky130_fd_sc_hs__a21oi_1_11/a_117_74#
+ sky130_fd_sc_hs__a21oi_1_11/a_29_368# sky130_fd_sc_hs__a21oi_1
Xsky130_fd_sc_hs__a21oi_1_21 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_33/Y sky130_fd_sc_hs__nand2_1_5/B
+ con_perb_3[0] sky130_fd_sc_hs__inv_4_29/Y sky130_fd_sc_hs__a21oi_1_21/a_117_74#
+ sky130_fd_sc_hs__a21oi_1_21/a_29_368# sky130_fd_sc_hs__a21oi_1
Xsky130_fd_sc_hs__a21oi_1_32 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_37/Y sky130_fd_sc_hs__nand2_2_73/B
+ con_perb_3[2] sky130_fd_sc_hs__inv_4_29/Y sky130_fd_sc_hs__a21oi_1_32/a_117_74#
+ sky130_fd_sc_hs__a21oi_1_32/a_29_368# sky130_fd_sc_hs__a21oi_1
Xsky130_fd_sc_hs__a21oi_1_43 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_31/Y sky130_fd_sc_hs__nand2_2_97/B
+ con_perb_1[0] sky130_fd_sc_hs__inv_4_29/Y sky130_fd_sc_hs__a21oi_1_43/a_117_74#
+ sky130_fd_sc_hs__a21oi_1_43/a_29_368# sky130_fd_sc_hs__a21oi_1
Xsky130_fd_sc_hs__dlygate4sd3_1_7 DVSS DVDD DVSS DVDD sky130_fd_sc_hs__dlygate4sd3_1_7/A
+ sky130_fd_sc_hs__dlygate4sd3_1_7/X sky130_fd_sc_hs__dlygate4sd3_1_7/a_405_138# sky130_fd_sc_hs__dlygate4sd3_1_7/a_28_74#
+ sky130_fd_sc_hs__dlygate4sd3_1_7/a_289_74# sky130_fd_sc_hs__dlygate4sd3_1
Xsky130_fd_sc_hs__einvp_1_1 DVSS DVDD DVDD DVSS pi3_l[0] sky130_fd_sc_hs__inv_8_1/A
+ sky130_fd_sc_hs__inv_4_3/Y sky130_fd_sc_hs__einvp_1_1/a_44_549# sky130_fd_sc_hs__einvp_1_1/a_318_74#
+ sky130_fd_sc_hs__einvp_1_1/a_310_392# sky130_fd_sc_hs__einvp_1
Xsky130_fd_sc_hs__inv_1_6 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_1_7/Y sky130_fd_sc_hs__inv_1_7/A
+ sky130_fd_sc_hs__inv_1
Xsky130_fd_sc_hs__nand2_8_0 DVSS DVDD DVDD DVSS inj_out osc_072 osc_108 sky130_fd_sc_hs__nand2_8_1/a_27_74#
+ sky130_fd_sc_hs__nand2_8
Xsky130_fd_sc_hs__nand2_1_7 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_1_7/B sky130_fd_sc_hs__nand2_1_7/Y
+ osc_072 sky130_fd_sc_hs__nand2_1_7/a_117_74# sky130_fd_sc_hs__nand2_1
Xsky130_fd_sc_hs__a21oi_1_11 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_37/Y sky130_fd_sc_hs__nand2_2_35/B
+ con_perb_5[2] sky130_fd_sc_hs__inv_4_29/Y sky130_fd_sc_hs__a21oi_1_11/a_117_74#
+ sky130_fd_sc_hs__a21oi_1_11/a_29_368# sky130_fd_sc_hs__a21oi_1
Xsky130_fd_sc_hs__a21oi_1_22 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_37/Y sky130_fd_sc_hs__nand2_2_57/B
+ con_perb_4[2] sky130_fd_sc_hs__inv_4_29/Y sky130_fd_sc_hs__a21oi_1_23/a_117_74#
+ sky130_fd_sc_hs__a21oi_1_23/a_29_368# sky130_fd_sc_hs__a21oi_1
Xsky130_fd_sc_hs__a21oi_1_33 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_39/Y sky130_fd_sc_hs__nand2_2_61/B
+ con_perb_3[3] sky130_fd_sc_hs__inv_4_29/Y sky130_fd_sc_hs__a21oi_1_33/a_117_74#
+ sky130_fd_sc_hs__a21oi_1_33/a_29_368# sky130_fd_sc_hs__a21oi_1
Xsky130_fd_sc_hs__a21oi_1_44 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_36/Y sky130_fd_sc_hs__a21oi_1_45/Y
+ con_perb_1[1] sky130_fd_sc_hs__inv_4_29/Y sky130_fd_sc_hs__a21oi_1_45/a_117_74#
+ sky130_fd_sc_hs__a21oi_1_45/a_29_368# sky130_fd_sc_hs__a21oi_1
Xsky130_fd_sc_hs__dlygate4sd3_1_8 DVSS DVDD DVSS DVDD sky130_fd_sc_hs__dlygate4sd3_1_9/A
+ sky130_fd_sc_hs__dlygate4sd3_1_9/X sky130_fd_sc_hs__dlygate4sd3_1_9/a_405_138# sky130_fd_sc_hs__dlygate4sd3_1_9/a_28_74#
+ sky130_fd_sc_hs__dlygate4sd3_1_9/a_289_74# sky130_fd_sc_hs__dlygate4sd3_1
Xsky130_fd_sc_hs__einvp_1_2 DVSS DVDD DVDD DVSS pi3_r[0] sky130_fd_sc_hs__inv_8_1/A
+ sky130_fd_sc_hs__inv_4_5/Y sky130_fd_sc_hs__einvp_1_3/a_44_549# sky130_fd_sc_hs__einvp_1_3/a_318_74#
+ sky130_fd_sc_hs__einvp_1_3/a_310_392# sky130_fd_sc_hs__einvp_1
Xsky130_fd_sc_hs__inv_8_0 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_8_1/A p3 sky130_fd_sc_hs__inv_8
Xsky130_fd_sc_hs__inv_1_7 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_1_7/Y sky130_fd_sc_hs__inv_1_7/A
+ sky130_fd_sc_hs__inv_1
Xsky130_fd_sc_hs__nand2_8_1 DVSS DVDD DVDD DVSS inj_out osc_072 osc_108 sky130_fd_sc_hs__nand2_8_1/a_27_74#
+ sky130_fd_sc_hs__nand2_8
Xsky130_fd_sc_hs__nand2_1_8 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_1_9/B sky130_fd_sc_hs__nand2_1_9/Y
+ osc_036 sky130_fd_sc_hs__nand2_1_9/a_117_74# sky130_fd_sc_hs__nand2_1
Xsky130_fd_sc_hs__a21oi_1_12 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_36/Y sky130_fd_sc_hs__nand2_2_37/B
+ con_perb_5[1] sky130_fd_sc_hs__inv_4_29/Y sky130_fd_sc_hs__a21oi_1_13/a_117_74#
+ sky130_fd_sc_hs__a21oi_1_13/a_29_368# sky130_fd_sc_hs__a21oi_1
Xsky130_fd_sc_hs__a21oi_1_23 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_37/Y sky130_fd_sc_hs__nand2_2_57/B
+ con_perb_4[2] sky130_fd_sc_hs__inv_4_29/Y sky130_fd_sc_hs__a21oi_1_23/a_117_74#
+ sky130_fd_sc_hs__a21oi_1_23/a_29_368# sky130_fd_sc_hs__a21oi_1
Xsky130_fd_sc_hs__a21oi_1_34 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_36/Y sky130_fd_sc_hs__nand2_2_88/B
+ con_perb_2[1] sky130_fd_sc_hs__inv_4_29/Y sky130_fd_sc_hs__a21oi_1_35/a_117_74#
+ sky130_fd_sc_hs__a21oi_1_35/a_29_368# sky130_fd_sc_hs__a21oi_1
Xsky130_fd_sc_hs__a21oi_1_45 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_36/Y sky130_fd_sc_hs__a21oi_1_45/Y
+ con_perb_1[1] sky130_fd_sc_hs__inv_4_29/Y sky130_fd_sc_hs__a21oi_1_45/a_117_74#
+ sky130_fd_sc_hs__a21oi_1_45/a_29_368# sky130_fd_sc_hs__a21oi_1
Xsky130_fd_sc_hs__dlygate4sd3_1_9 DVSS DVDD DVSS DVDD sky130_fd_sc_hs__dlygate4sd3_1_9/A
+ sky130_fd_sc_hs__dlygate4sd3_1_9/X sky130_fd_sc_hs__dlygate4sd3_1_9/a_405_138# sky130_fd_sc_hs__dlygate4sd3_1_9/a_28_74#
+ sky130_fd_sc_hs__dlygate4sd3_1_9/a_289_74# sky130_fd_sc_hs__dlygate4sd3_1
Xsky130_fd_sc_hs__einvp_1_3 DVSS DVDD DVDD DVSS pi3_r[0] sky130_fd_sc_hs__inv_8_1/A
+ sky130_fd_sc_hs__inv_4_5/Y sky130_fd_sc_hs__einvp_1_3/a_44_549# sky130_fd_sc_hs__einvp_1_3/a_318_74#
+ sky130_fd_sc_hs__einvp_1_3/a_310_392# sky130_fd_sc_hs__einvp_1
Xsky130_fd_sc_hs__inv_8_1 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_8_1/A p3 sky130_fd_sc_hs__inv_8
Xsky130_fd_sc_hs__inv_1_8 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_1_9/Y sky130_fd_sc_hs__inv_1_9/A
+ sky130_fd_sc_hs__inv_1
Xsky130_fd_sc_hs__nand2_8_2 DVSS DVDD DVDD DVSS osc_hold osc_036 osc_072 sky130_fd_sc_hs__nand2_8_3/a_27_74#
+ sky130_fd_sc_hs__nand2_8
Xsky130_fd_sc_hs__nand2_1_9 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_1_9/B sky130_fd_sc_hs__nand2_1_9/Y
+ osc_036 sky130_fd_sc_hs__nand2_1_9/a_117_74# sky130_fd_sc_hs__nand2_1
Xsky130_fd_sc_hs__a21oi_1_13 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_36/Y sky130_fd_sc_hs__nand2_2_37/B
+ con_perb_5[1] sky130_fd_sc_hs__inv_4_29/Y sky130_fd_sc_hs__a21oi_1_13/a_117_74#
+ sky130_fd_sc_hs__a21oi_1_13/a_29_368# sky130_fd_sc_hs__a21oi_1
Xsky130_fd_sc_hs__a21oi_1_24 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_36/Y sky130_fd_sc_hs__nand2_2_45/B
+ con_perb_3[1] sky130_fd_sc_hs__inv_4_29/Y sky130_fd_sc_hs__a21oi_1_25/a_117_74#
+ sky130_fd_sc_hs__a21oi_1_25/a_29_368# sky130_fd_sc_hs__a21oi_1
Xsky130_fd_sc_hs__a21oi_1_35 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_36/Y sky130_fd_sc_hs__nand2_2_88/B
+ con_perb_2[1] sky130_fd_sc_hs__inv_4_29/Y sky130_fd_sc_hs__a21oi_1_35/a_117_74#
+ sky130_fd_sc_hs__a21oi_1_35/a_29_368# sky130_fd_sc_hs__a21oi_1
Xsky130_fd_sc_hs__a21oi_1_46 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_39/Y sky130_fd_sc_hs__nand2_2_99/B
+ con_perb_1[3] sky130_fd_sc_hs__inv_4_29/Y sky130_fd_sc_hs__a21oi_1_47/a_117_74#
+ sky130_fd_sc_hs__a21oi_1_47/a_29_368# sky130_fd_sc_hs__a21oi_1
Xsky130_fd_sc_hs__einvp_1_4 DVSS DVDD DVDD DVSS pi2_l[0] sky130_fd_sc_hs__inv_8_3/A
+ sky130_fd_sc_hs__inv_4_7/Y sky130_fd_sc_hs__einvp_1_5/a_44_549# sky130_fd_sc_hs__einvp_1_5/a_318_74#
+ sky130_fd_sc_hs__einvp_1_5/a_310_392# sky130_fd_sc_hs__einvp_1
Xsky130_fd_sc_hs__inv_8_2 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_8_3/A p2 sky130_fd_sc_hs__inv_8
Xsky130_fd_sc_hs__inv_1_9 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_1_9/Y sky130_fd_sc_hs__inv_1_9/A
+ sky130_fd_sc_hs__inv_1
Xsky130_fd_sc_hs__nand2_8_3 DVSS DVDD DVDD DVSS osc_hold osc_036 osc_072 sky130_fd_sc_hs__nand2_8_3/a_27_74#
+ sky130_fd_sc_hs__nand2_8
Xsky130_fd_sc_hs__a21oi_1_14 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_31/Y sky130_fd_sc_hs__nand2_2_43/B
+ con_perb_3[0] sky130_fd_sc_hs__inv_4_29/Y sky130_fd_sc_hs__a21oi_1_15/a_117_74#
+ sky130_fd_sc_hs__a21oi_1_15/a_29_368# sky130_fd_sc_hs__a21oi_1
Xsky130_fd_sc_hs__a21oi_1_25 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_36/Y sky130_fd_sc_hs__nand2_2_45/B
+ con_perb_3[1] sky130_fd_sc_hs__inv_4_29/Y sky130_fd_sc_hs__a21oi_1_25/a_117_74#
+ sky130_fd_sc_hs__a21oi_1_25/a_29_368# sky130_fd_sc_hs__a21oi_1
Xsky130_fd_sc_hs__a21oi_1_36 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_37/Y sky130_fd_sc_hs__nand2_2_84/B
+ con_perb_2[2] sky130_fd_sc_hs__inv_4_29/Y sky130_fd_sc_hs__a21oi_1_37/a_117_74#
+ sky130_fd_sc_hs__a21oi_1_37/a_29_368# sky130_fd_sc_hs__a21oi_1
Xsky130_fd_sc_hs__a21oi_1_47 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_39/Y sky130_fd_sc_hs__nand2_2_99/B
+ con_perb_1[3] sky130_fd_sc_hs__inv_4_29/Y sky130_fd_sc_hs__a21oi_1_47/a_117_74#
+ sky130_fd_sc_hs__a21oi_1_47/a_29_368# sky130_fd_sc_hs__a21oi_1
Xsky130_fd_sc_hs__dlygate4sd2_1_0 DVSS DVDD DVSS DVDD sky130_fd_sc_hs__dlygate4sd2_1_1/A
+ sky130_fd_sc_hs__dlygate4sd2_1_1/X sky130_fd_sc_hs__dlygate4sd2_1_1/a_405_138# sky130_fd_sc_hs__dlygate4sd2_1_1/a_28_74#
+ sky130_fd_sc_hs__dlygate4sd2_1_1/a_288_74# sky130_fd_sc_hs__dlygate4sd2_1
Xsky130_fd_sc_hs__einvp_1_5 DVSS DVDD DVDD DVSS pi2_l[0] sky130_fd_sc_hs__inv_8_3/A
+ sky130_fd_sc_hs__inv_4_7/Y sky130_fd_sc_hs__einvp_1_5/a_44_549# sky130_fd_sc_hs__einvp_1_5/a_318_74#
+ sky130_fd_sc_hs__einvp_1_5/a_310_392# sky130_fd_sc_hs__einvp_1
Xsky130_fd_sc_hs__inv_8_3 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_8_3/A p2 sky130_fd_sc_hs__inv_8
Xsky130_fd_sc_hs__nand2_4_90 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_4_91/Y delay_con_msb[1]
+ osc_108 sky130_fd_sc_hs__nand2_4_91/a_27_74# sky130_fd_sc_hs__nand2_4
Xsky130_fd_sc_hs__nand2_8_4 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_8_9/B osc_108
+ osc_144 sky130_fd_sc_hs__nand2_8_5/a_27_74# sky130_fd_sc_hs__nand2_8
Xsky130_fd_sc_hs__a21oi_1_15 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_31/Y sky130_fd_sc_hs__nand2_2_43/B
+ con_perb_3[0] sky130_fd_sc_hs__inv_4_29/Y sky130_fd_sc_hs__a21oi_1_15/a_117_74#
+ sky130_fd_sc_hs__a21oi_1_15/a_29_368# sky130_fd_sc_hs__a21oi_1
Xsky130_fd_sc_hs__a21oi_1_26 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_33/Y sky130_fd_sc_hs__nand2_1_7/B
+ con_perb_2[0] sky130_fd_sc_hs__inv_4_29/Y sky130_fd_sc_hs__a21oi_1_28/a_117_74#
+ sky130_fd_sc_hs__a21oi_1_28/a_29_368# sky130_fd_sc_hs__a21oi_1
Xsky130_fd_sc_hs__a21oi_1_37 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_37/Y sky130_fd_sc_hs__nand2_2_84/B
+ con_perb_2[2] sky130_fd_sc_hs__inv_4_29/Y sky130_fd_sc_hs__a21oi_1_37/a_117_74#
+ sky130_fd_sc_hs__a21oi_1_37/a_29_368# sky130_fd_sc_hs__a21oi_1
Xsky130_fd_sc_hs__a21oi_1_48 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_37/Y sky130_fd_sc_hs__a21oi_1_49/Y
+ con_perb_1[2] sky130_fd_sc_hs__inv_4_29/Y sky130_fd_sc_hs__a21oi_1_49/a_117_74#
+ sky130_fd_sc_hs__a21oi_1_49/a_29_368# sky130_fd_sc_hs__a21oi_1
Xsky130_fd_sc_hs__dlygate4sd3_1_70 DVSS DVDD DVSS DVDD inj_en sky130_fd_sc_hs__dlygate4sd3_1_71/X
+ sky130_fd_sc_hs__dlygate4sd3_1_71/a_405_138# sky130_fd_sc_hs__dlygate4sd3_1_71/a_28_74#
+ sky130_fd_sc_hs__dlygate4sd3_1_71/a_289_74# sky130_fd_sc_hs__dlygate4sd3_1
Xsky130_fd_sc_hs__dlygate4sd2_1_1 DVSS DVDD DVSS DVDD sky130_fd_sc_hs__dlygate4sd2_1_1/A
+ sky130_fd_sc_hs__dlygate4sd2_1_1/X sky130_fd_sc_hs__dlygate4sd2_1_1/a_405_138# sky130_fd_sc_hs__dlygate4sd2_1_1/a_28_74#
+ sky130_fd_sc_hs__dlygate4sd2_1_1/a_288_74# sky130_fd_sc_hs__dlygate4sd2_1
Xsky130_fd_sc_hs__einvp_1_6 DVSS DVDD DVDD DVSS pi2_r[0] sky130_fd_sc_hs__inv_8_3/A
+ sky130_fd_sc_hs__inv_4_9/Y sky130_fd_sc_hs__einvp_1_7/a_44_549# sky130_fd_sc_hs__einvp_1_7/a_318_74#
+ sky130_fd_sc_hs__einvp_1_7/a_310_392# sky130_fd_sc_hs__einvp_1
Xsky130_fd_sc_hs__inv_8_4 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_8_5/A p4 sky130_fd_sc_hs__inv_8
Xsky130_fd_sc_hs__nand2_4_80 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_4_81/Y delay_con_msb[2]
+ osc_108 sky130_fd_sc_hs__nand2_4_81/a_27_74# sky130_fd_sc_hs__nand2_4
Xsky130_fd_sc_hs__nand2_4_91 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_4_91/Y delay_con_msb[1]
+ osc_108 sky130_fd_sc_hs__nand2_4_91/a_27_74# sky130_fd_sc_hs__nand2_4
Xsky130_fd_sc_hs__nand2_8_5 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_8_9/B osc_108
+ osc_144 sky130_fd_sc_hs__nand2_8_5/a_27_74# sky130_fd_sc_hs__nand2_8
Xsky130_fd_sc_hs__a21oi_1_16 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_39/Y sky130_fd_sc_hs__nand2_2_65/B
+ con_perb_4[3] sky130_fd_sc_hs__inv_4_29/Y sky130_fd_sc_hs__a21oi_1_17/a_117_74#
+ sky130_fd_sc_hs__a21oi_1_17/a_29_368# sky130_fd_sc_hs__a21oi_1
Xsky130_fd_sc_hs__a21oi_1_27 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_31/Y sky130_fd_sc_hs__nand2_2_79/B
+ con_perb_2[0] sky130_fd_sc_hs__inv_4_29/Y sky130_fd_sc_hs__a21oi_1_29/a_117_74#
+ sky130_fd_sc_hs__a21oi_1_29/a_29_368# sky130_fd_sc_hs__a21oi_1
Xsky130_fd_sc_hs__a21oi_1_38 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_39/Y sky130_fd_sc_hs__nand2_2_85/B
+ con_perb_2[3] sky130_fd_sc_hs__inv_4_29/Y sky130_fd_sc_hs__a21oi_1_39/a_117_74#
+ sky130_fd_sc_hs__a21oi_1_39/a_29_368# sky130_fd_sc_hs__a21oi_1
Xsky130_fd_sc_hs__a21oi_1_49 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_37/Y sky130_fd_sc_hs__a21oi_1_49/Y
+ con_perb_1[2] sky130_fd_sc_hs__inv_4_29/Y sky130_fd_sc_hs__a21oi_1_49/a_117_74#
+ sky130_fd_sc_hs__a21oi_1_49/a_29_368# sky130_fd_sc_hs__a21oi_1
Xsky130_fd_sc_hs__dlygate4sd3_1_60 DVSS DVDD DVSS DVDD sky130_fd_sc_hs__dlygate4sd3_1_68/X
+ sky130_fd_sc_hs__dlygate4sd3_1_62/X sky130_fd_sc_hs__dlygate4sd3_1_62/a_405_138#
+ sky130_fd_sc_hs__dlygate4sd3_1_62/a_28_74# sky130_fd_sc_hs__dlygate4sd3_1_62/a_289_74#
+ sky130_fd_sc_hs__dlygate4sd3_1
Xsky130_fd_sc_hs__dlygate4sd3_1_71 DVSS DVDD DVSS DVDD inj_en sky130_fd_sc_hs__dlygate4sd3_1_71/X
+ sky130_fd_sc_hs__dlygate4sd3_1_71/a_405_138# sky130_fd_sc_hs__dlygate4sd3_1_71/a_28_74#
+ sky130_fd_sc_hs__dlygate4sd3_1_71/a_289_74# sky130_fd_sc_hs__dlygate4sd3_1
Xsky130_fd_sc_hs__einvp_8_0 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_8_1/A pi3_l[3]
+ sky130_fd_sc_hs__inv_4_3/Y sky130_fd_sc_hs__einvp_8_2/a_802_323# sky130_fd_sc_hs__einvp_8_2/a_27_74#
+ sky130_fd_sc_hs__einvp_8_2/a_27_368# sky130_fd_sc_hs__einvp_8
Xsky130_fd_sc_hs__einvp_1_7 DVSS DVDD DVDD DVSS pi2_r[0] sky130_fd_sc_hs__inv_8_3/A
+ sky130_fd_sc_hs__inv_4_9/Y sky130_fd_sc_hs__einvp_1_7/a_44_549# sky130_fd_sc_hs__einvp_1_7/a_318_74#
+ sky130_fd_sc_hs__einvp_1_7/a_310_392# sky130_fd_sc_hs__einvp_1
Xsky130_fd_sc_hs__inv_8_5 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_8_5/A p4 sky130_fd_sc_hs__inv_8
Xsky130_fd_sc_hs__nand2_4_70 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_4_71/Y delay_con_msb[1]
+ osc_108 sky130_fd_sc_hs__nand2_4_71/a_27_74# sky130_fd_sc_hs__nand2_4
Xsky130_fd_sc_hs__nand2_4_81 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_4_81/Y delay_con_msb[2]
+ osc_108 sky130_fd_sc_hs__nand2_4_81/a_27_74# sky130_fd_sc_hs__nand2_4
Xsky130_fd_sc_hs__nand2_4_92 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_4_93/Y delay_con_msb[2]
+ osc_108 sky130_fd_sc_hs__nand2_4_93/a_27_74# sky130_fd_sc_hs__nand2_4
Xsky130_fd_sc_hs__nand2_8_6 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_8_9/B osc_000
+ osc_036 sky130_fd_sc_hs__nand2_8_7/a_27_74# sky130_fd_sc_hs__nand2_8
Xsky130_fd_sc_hs__a21oi_1_17 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_39/Y sky130_fd_sc_hs__nand2_2_65/B
+ con_perb_4[3] sky130_fd_sc_hs__inv_4_29/Y sky130_fd_sc_hs__a21oi_1_17/a_117_74#
+ sky130_fd_sc_hs__a21oi_1_17/a_29_368# sky130_fd_sc_hs__a21oi_1
Xsky130_fd_sc_hs__a21oi_1_28 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_33/Y sky130_fd_sc_hs__nand2_1_7/B
+ con_perb_2[0] sky130_fd_sc_hs__inv_4_29/Y sky130_fd_sc_hs__a21oi_1_28/a_117_74#
+ sky130_fd_sc_hs__a21oi_1_28/a_29_368# sky130_fd_sc_hs__a21oi_1
Xsky130_fd_sc_hs__a21oi_1_39 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_39/Y sky130_fd_sc_hs__nand2_2_85/B
+ con_perb_2[3] sky130_fd_sc_hs__inv_4_29/Y sky130_fd_sc_hs__a21oi_1_39/a_117_74#
+ sky130_fd_sc_hs__a21oi_1_39/a_29_368# sky130_fd_sc_hs__a21oi_1
Xsky130_fd_sc_hs__bufbuf_8_0 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__clkbuf_4_3/X sky130_fd_sc_hs__bufbuf_8_1/X
+ sky130_fd_sc_hs__bufbuf_8_1/a_334_368# sky130_fd_sc_hs__bufbuf_8_1/a_27_112# sky130_fd_sc_hs__bufbuf_8_1/a_221_368#
+ sky130_fd_sc_hs__bufbuf_8
Xsky130_fd_sc_hs__dlygate4sd3_1_50 DVSS DVDD DVSS DVDD sky130_fd_sc_hs__dlygate4sd3_1_57/X
+ sky130_fd_sc_hs__dlygate4sd3_1_51/X sky130_fd_sc_hs__dlygate4sd3_1_51/a_405_138#
+ sky130_fd_sc_hs__dlygate4sd3_1_51/a_28_74# sky130_fd_sc_hs__dlygate4sd3_1_51/a_289_74#
+ sky130_fd_sc_hs__dlygate4sd3_1
Xsky130_fd_sc_hs__dlygate4sd3_1_61 DVSS DVDD DVSS DVDD sky130_fd_sc_hs__dlygate4sd3_1_63/A
+ sky130_fd_sc_hs__dlygate4sd3_1_68/A sky130_fd_sc_hs__dlygate4sd3_1_63/a_405_138#
+ sky130_fd_sc_hs__dlygate4sd3_1_63/a_28_74# sky130_fd_sc_hs__dlygate4sd3_1_63/a_289_74#
+ sky130_fd_sc_hs__dlygate4sd3_1
Xsky130_fd_sc_hs__dlygate4sd3_1_72 DVSS DVDD DVSS DVDD sky130_fd_sc_hs__dlygate4sd3_1_78/X
+ sky130_fd_sc_hs__clkbuf_4_1/A sky130_fd_sc_hs__dlygate4sd3_1_74/a_405_138# sky130_fd_sc_hs__dlygate4sd3_1_74/a_28_74#
+ sky130_fd_sc_hs__dlygate4sd3_1_74/a_289_74# sky130_fd_sc_hs__dlygate4sd3_1
Xsky130_fd_sc_hs__nand2_4_0 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_4_1/Y delay_con_msb[3]
+ osc_144 sky130_fd_sc_hs__nand2_4_1/a_27_74# sky130_fd_sc_hs__nand2_4
Xsky130_fd_sc_hs__einvp_8_1 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_8_1/A pi3_r[3]
+ sky130_fd_sc_hs__inv_4_5/Y sky130_fd_sc_hs__einvp_8_3/a_802_323# sky130_fd_sc_hs__einvp_8_3/a_27_74#
+ sky130_fd_sc_hs__einvp_8_3/a_27_368# sky130_fd_sc_hs__einvp_8
Xsky130_fd_sc_hs__einvp_1_8 DVSS DVDD DVDD DVSS pi4_l[0] sky130_fd_sc_hs__inv_8_5/A
+ sky130_fd_sc_hs__inv_4_11/Y sky130_fd_sc_hs__einvp_1_9/a_44_549# sky130_fd_sc_hs__einvp_1_9/a_318_74#
+ sky130_fd_sc_hs__einvp_1_9/a_310_392# sky130_fd_sc_hs__einvp_1
Xsky130_fd_sc_hs__einvp_1_10 DVSS DVDD DVDD DVSS pi4_r[0] sky130_fd_sc_hs__inv_8_5/A
+ sky130_fd_sc_hs__inv_4_13/Y sky130_fd_sc_hs__einvp_1_11/a_44_549# sky130_fd_sc_hs__einvp_1_11/a_318_74#
+ sky130_fd_sc_hs__einvp_1_11/a_310_392# sky130_fd_sc_hs__einvp_1
Xsky130_fd_sc_hs__inv_8_6 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_8_7/A p1 sky130_fd_sc_hs__inv_8
Xsky130_fd_sc_hs__nand2_4_60 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_4_60/Y delay_con_msb[3]
+ osc_108 sky130_fd_sc_hs__nand2_4_60/a_27_74# sky130_fd_sc_hs__nand2_4
Xsky130_fd_sc_hs__nand2_4_71 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_4_71/Y delay_con_msb[1]
+ osc_108 sky130_fd_sc_hs__nand2_4_71/a_27_74# sky130_fd_sc_hs__nand2_4
Xsky130_fd_sc_hs__nand2_4_82 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_4_83/Y delay_con_msb[2]
+ osc_108 sky130_fd_sc_hs__nand2_4_83/a_27_74# sky130_fd_sc_hs__nand2_4
Xsky130_fd_sc_hs__nand2_4_93 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_4_93/Y delay_con_msb[2]
+ osc_108 sky130_fd_sc_hs__nand2_4_93/a_27_74# sky130_fd_sc_hs__nand2_4
Xsky130_fd_sc_hs__buf_4_0 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__buf_4_1/A sky130_fd_sc_hs__buf_4_1/X
+ sky130_fd_sc_hs__buf_4_1/a_86_260# sky130_fd_sc_hs__buf_4
Xsky130_fd_sc_hs__nand2_8_7 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_8_9/B osc_000
+ osc_036 sky130_fd_sc_hs__nand2_8_7/a_27_74# sky130_fd_sc_hs__nand2_8
Xsky130_fd_sc_hs__inv_4_0 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_1/Y ref_clk sky130_fd_sc_hs__inv_4
Xsky130_fd_sc_hs__a21oi_1_18 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_36/Y sky130_fd_sc_hs__nand2_2_71/B
+ con_perb_4[1] sky130_fd_sc_hs__inv_4_29/Y sky130_fd_sc_hs__a21oi_1_19/a_117_74#
+ sky130_fd_sc_hs__a21oi_1_19/a_29_368# sky130_fd_sc_hs__a21oi_1
Xsky130_fd_sc_hs__a21oi_1_29 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_31/Y sky130_fd_sc_hs__nand2_2_79/B
+ con_perb_2[0] sky130_fd_sc_hs__inv_4_29/Y sky130_fd_sc_hs__a21oi_1_29/a_117_74#
+ sky130_fd_sc_hs__a21oi_1_29/a_29_368# sky130_fd_sc_hs__a21oi_1
Xsky130_fd_sc_hs__bufbuf_8_1 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__clkbuf_4_3/X sky130_fd_sc_hs__bufbuf_8_1/X
+ sky130_fd_sc_hs__bufbuf_8_1/a_334_368# sky130_fd_sc_hs__bufbuf_8_1/a_27_112# sky130_fd_sc_hs__bufbuf_8_1/a_221_368#
+ sky130_fd_sc_hs__bufbuf_8
Xsky130_fd_sc_hs__einvp_4_10 DVSS DVDD DVDD DVSS pi4_r[2] sky130_fd_sc_hs__inv_8_5/A
+ sky130_fd_sc_hs__inv_4_13/Y sky130_fd_sc_hs__einvp_4_11/a_27_74# sky130_fd_sc_hs__einvp_4_11/a_27_368#
+ sky130_fd_sc_hs__einvp_4_11/a_473_323# sky130_fd_sc_hs__einvp_4
Xsky130_fd_sc_hs__dlygate4sd3_1_40 DVSS DVDD DVSS DVDD sky130_fd_sc_hs__bufbuf_8_1/X
+ sky130_fd_sc_hs__dlygate4sd3_1_75/A sky130_fd_sc_hs__dlygate4sd3_1_41/a_405_138#
+ sky130_fd_sc_hs__dlygate4sd3_1_41/a_28_74# sky130_fd_sc_hs__dlygate4sd3_1_41/a_289_74#
+ sky130_fd_sc_hs__dlygate4sd3_1
Xsky130_fd_sc_hs__dlygate4sd3_1_51 DVSS DVDD DVSS DVDD sky130_fd_sc_hs__dlygate4sd3_1_57/X
+ sky130_fd_sc_hs__dlygate4sd3_1_51/X sky130_fd_sc_hs__dlygate4sd3_1_51/a_405_138#
+ sky130_fd_sc_hs__dlygate4sd3_1_51/a_28_74# sky130_fd_sc_hs__dlygate4sd3_1_51/a_289_74#
+ sky130_fd_sc_hs__dlygate4sd3_1
Xsky130_fd_sc_hs__dlygate4sd3_1_62 DVSS DVDD DVSS DVDD sky130_fd_sc_hs__dlygate4sd3_1_68/X
+ sky130_fd_sc_hs__dlygate4sd3_1_62/X sky130_fd_sc_hs__dlygate4sd3_1_62/a_405_138#
+ sky130_fd_sc_hs__dlygate4sd3_1_62/a_28_74# sky130_fd_sc_hs__dlygate4sd3_1_62/a_289_74#
+ sky130_fd_sc_hs__dlygate4sd3_1
Xsky130_fd_sc_hs__dlygate4sd3_1_73 DVSS DVDD DVSS DVDD sky130_fd_sc_hs__dlygate4sd3_1_75/A
+ sky130_fd_sc_hs__dlygate4sd3_1_75/X sky130_fd_sc_hs__dlygate4sd3_1_75/a_405_138#
+ sky130_fd_sc_hs__dlygate4sd3_1_75/a_28_74# sky130_fd_sc_hs__dlygate4sd3_1_75/a_289_74#
+ sky130_fd_sc_hs__dlygate4sd3_1
Xsky130_fd_sc_hs__nand2_4_1 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_4_1/Y delay_con_msb[3]
+ osc_144 sky130_fd_sc_hs__nand2_4_1/a_27_74# sky130_fd_sc_hs__nand2_4
Xsky130_fd_sc_hs__nand2_2_100 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_2_102/Y sky130_fd_sc_hs__nand2_2_99/B
+ osc_036 sky130_fd_sc_hs__nand2_2_102/a_27_74# sky130_fd_sc_hs__nand2_2
Xsky130_fd_sc_hs__einvp_8_2 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_8_1/A pi3_l[3]
+ sky130_fd_sc_hs__inv_4_3/Y sky130_fd_sc_hs__einvp_8_2/a_802_323# sky130_fd_sc_hs__einvp_8_2/a_27_74#
+ sky130_fd_sc_hs__einvp_8_2/a_27_368# sky130_fd_sc_hs__einvp_8
Xsky130_fd_sc_hs__einvp_1_9 DVSS DVDD DVDD DVSS pi4_l[0] sky130_fd_sc_hs__inv_8_5/A
+ sky130_fd_sc_hs__inv_4_11/Y sky130_fd_sc_hs__einvp_1_9/a_44_549# sky130_fd_sc_hs__einvp_1_9/a_318_74#
+ sky130_fd_sc_hs__einvp_1_9/a_310_392# sky130_fd_sc_hs__einvp_1
Xsky130_fd_sc_hs__einvp_1_11 DVSS DVDD DVDD DVSS pi4_r[0] sky130_fd_sc_hs__inv_8_5/A
+ sky130_fd_sc_hs__inv_4_13/Y sky130_fd_sc_hs__einvp_1_11/a_44_549# sky130_fd_sc_hs__einvp_1_11/a_318_74#
+ sky130_fd_sc_hs__einvp_1_11/a_310_392# sky130_fd_sc_hs__einvp_1
Xsky130_fd_sc_hs__inv_8_7 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_8_7/A p1 sky130_fd_sc_hs__inv_8
Xsky130_fd_sc_hs__nand2_4_50 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_4_51/Y delay_con_msb[3]
+ osc_108 sky130_fd_sc_hs__nand2_4_51/a_27_74# sky130_fd_sc_hs__nand2_4
Xsky130_fd_sc_hs__nand2_4_61 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_4_61/Y delay_con_msb[3]
+ osc_108 sky130_fd_sc_hs__nand2_4_61/a_27_74# sky130_fd_sc_hs__nand2_4
Xsky130_fd_sc_hs__nand2_4_72 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_4_73/Y delay_con_msb[2]
+ osc_108 sky130_fd_sc_hs__nand2_4_73/a_27_74# sky130_fd_sc_hs__nand2_4
Xsky130_fd_sc_hs__nand2_4_83 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_4_83/Y delay_con_msb[2]
+ osc_108 sky130_fd_sc_hs__nand2_4_83/a_27_74# sky130_fd_sc_hs__nand2_4
Xsky130_fd_sc_hs__nand2_4_94 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_4_95/Y delay_con_msb[2]
+ osc_072 sky130_fd_sc_hs__nand2_4_95/a_27_74# sky130_fd_sc_hs__nand2_4
Xsky130_fd_sc_hs__buf_4_1 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__buf_4_1/A sky130_fd_sc_hs__buf_4_1/X
+ sky130_fd_sc_hs__buf_4_1/a_86_260# sky130_fd_sc_hs__buf_4
Xsky130_fd_sc_hs__nand2_8_8 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_8_9/B osc_144
+ osc_000 sky130_fd_sc_hs__nand2_8_9/a_27_74# sky130_fd_sc_hs__nand2_8
Xsky130_fd_sc_hs__inv_4_1 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_1/Y ref_clk sky130_fd_sc_hs__inv_4
Xsky130_fd_sc_hs__a21oi_1_19 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_36/Y sky130_fd_sc_hs__nand2_2_71/B
+ con_perb_4[1] sky130_fd_sc_hs__inv_4_29/Y sky130_fd_sc_hs__a21oi_1_19/a_117_74#
+ sky130_fd_sc_hs__a21oi_1_19/a_29_368# sky130_fd_sc_hs__a21oi_1
Xsky130_fd_sc_hs__einvp_4_11 DVSS DVDD DVDD DVSS pi4_r[2] sky130_fd_sc_hs__inv_8_5/A
+ sky130_fd_sc_hs__inv_4_13/Y sky130_fd_sc_hs__einvp_4_11/a_27_74# sky130_fd_sc_hs__einvp_4_11/a_27_368#
+ sky130_fd_sc_hs__einvp_4_11/a_473_323# sky130_fd_sc_hs__einvp_4
Xsky130_fd_sc_hs__dlygate4sd3_1_41 DVSS DVDD DVSS DVDD sky130_fd_sc_hs__bufbuf_8_1/X
+ sky130_fd_sc_hs__dlygate4sd3_1_75/A sky130_fd_sc_hs__dlygate4sd3_1_41/a_405_138#
+ sky130_fd_sc_hs__dlygate4sd3_1_41/a_28_74# sky130_fd_sc_hs__dlygate4sd3_1_41/a_289_74#
+ sky130_fd_sc_hs__dlygate4sd3_1
Xsky130_fd_sc_hs__dlygate4sd3_1_52 DVSS DVDD DVSS DVDD sky130_fd_sc_hs__dlygate4sd3_1_53/A
+ sky130_fd_sc_hs__dlygate4sd3_1_53/X sky130_fd_sc_hs__dlygate4sd3_1_53/a_405_138#
+ sky130_fd_sc_hs__dlygate4sd3_1_53/a_28_74# sky130_fd_sc_hs__dlygate4sd3_1_53/a_289_74#
+ sky130_fd_sc_hs__dlygate4sd3_1
Xsky130_fd_sc_hs__dlygate4sd3_1_63 DVSS DVDD DVSS DVDD sky130_fd_sc_hs__dlygate4sd3_1_63/A
+ sky130_fd_sc_hs__dlygate4sd3_1_68/A sky130_fd_sc_hs__dlygate4sd3_1_63/a_405_138#
+ sky130_fd_sc_hs__dlygate4sd3_1_63/a_28_74# sky130_fd_sc_hs__dlygate4sd3_1_63/a_289_74#
+ sky130_fd_sc_hs__dlygate4sd3_1
Xsky130_fd_sc_hs__dlygate4sd3_1_74 DVSS DVDD DVSS DVDD sky130_fd_sc_hs__dlygate4sd3_1_78/X
+ sky130_fd_sc_hs__clkbuf_4_1/A sky130_fd_sc_hs__dlygate4sd3_1_74/a_405_138# sky130_fd_sc_hs__dlygate4sd3_1_74/a_28_74#
+ sky130_fd_sc_hs__dlygate4sd3_1_74/a_289_74# sky130_fd_sc_hs__dlygate4sd3_1
Xsky130_fd_sc_hs__dlygate4sd3_1_30 DVSS DVDD DVSS DVDD sky130_fd_sc_hs__dlygate4sd3_1_43/X
+ sky130_fd_sc_hs__dlygate4sd3_1_31/X sky130_fd_sc_hs__dlygate4sd3_1_31/a_405_138#
+ sky130_fd_sc_hs__dlygate4sd3_1_31/a_28_74# sky130_fd_sc_hs__dlygate4sd3_1_31/a_289_74#
+ sky130_fd_sc_hs__dlygate4sd3_1
Xsky130_fd_sc_hs__nand2_4_2 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_4_3/Y delay_con_msb[3]
+ osc_000 sky130_fd_sc_hs__nand2_4_3/a_27_74# sky130_fd_sc_hs__nand2_4
Xsky130_fd_sc_hs__nand2_2_101 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_2_103/Y sky130_fd_sc_hs__nand2_2_99/B
+ osc_036 sky130_fd_sc_hs__nand2_2_103/a_27_74# sky130_fd_sc_hs__nand2_2
Xsky130_fd_sc_hs__einvp_8_3 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_8_1/A pi3_r[3]
+ sky130_fd_sc_hs__inv_4_5/Y sky130_fd_sc_hs__einvp_8_3/a_802_323# sky130_fd_sc_hs__einvp_8_3/a_27_74#
+ sky130_fd_sc_hs__einvp_8_3/a_27_368# sky130_fd_sc_hs__einvp_8
Xsky130_fd_sc_hs__inv_16_30 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__and4_2_3/C sky130_fd_sc_hs__inv_16_31/A
+ sky130_fd_sc_hs__inv_16
Xsky130_fd_sc_hs__einvp_1_12 DVSS DVDD DVDD DVSS pi1_l[0] sky130_fd_sc_hs__inv_8_7/A
+ sky130_fd_sc_hs__inv_4_15/Y sky130_fd_sc_hs__einvp_1_13/a_44_549# sky130_fd_sc_hs__einvp_1_13/a_318_74#
+ sky130_fd_sc_hs__einvp_1_13/a_310_392# sky130_fd_sc_hs__einvp_1
Xsky130_fd_sc_hs__inv_8_8 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_8_9/A p5 sky130_fd_sc_hs__inv_8
Xsky130_fd_sc_hs__nand2_4_40 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_4_40/Y delay_con_msb[2]
+ osc_000 sky130_fd_sc_hs__nand2_4_40/a_27_74# sky130_fd_sc_hs__nand2_4
Xsky130_fd_sc_hs__nand2_4_51 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_4_51/Y delay_con_msb[3]
+ osc_108 sky130_fd_sc_hs__nand2_4_51/a_27_74# sky130_fd_sc_hs__nand2_4
Xsky130_fd_sc_hs__nand2_4_62 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_4_63/Y delay_con_msb[0]
+ osc_144 sky130_fd_sc_hs__nand2_4_63/a_27_74# sky130_fd_sc_hs__nand2_4
Xsky130_fd_sc_hs__nand2_4_73 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_4_73/Y delay_con_msb[2]
+ osc_108 sky130_fd_sc_hs__nand2_4_73/a_27_74# sky130_fd_sc_hs__nand2_4
Xsky130_fd_sc_hs__nand2_4_84 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_4_85/Y delay_con_msb[0]
+ osc_108 sky130_fd_sc_hs__nand2_4_85/a_27_74# sky130_fd_sc_hs__nand2_4
Xsky130_fd_sc_hs__nand2_4_95 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_4_95/Y delay_con_msb[2]
+ osc_072 sky130_fd_sc_hs__nand2_4_95/a_27_74# sky130_fd_sc_hs__nand2_4
Xsky130_fd_sc_hs__clkbuf_4_0 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__clkbuf_4_1/A sky130_fd_sc_hs__nand2_8_9/B
+ sky130_fd_sc_hs__clkbuf_4_1/a_83_270# sky130_fd_sc_hs__clkbuf_4
Xsky130_fd_sc_hs__inv_4_2 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_3/Y osc_072 sky130_fd_sc_hs__inv_4
Xsky130_fd_sc_hs__nand2_8_9 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_8_9/B osc_144
+ osc_000 sky130_fd_sc_hs__nand2_8_9/a_27_74# sky130_fd_sc_hs__nand2_8
Xsky130_fd_sc_hs__einvp_4_12 DVSS DVDD DVDD DVSS pi1_l[2] sky130_fd_sc_hs__inv_8_7/A
+ sky130_fd_sc_hs__inv_4_15/Y sky130_fd_sc_hs__einvp_4_13/a_27_74# sky130_fd_sc_hs__einvp_4_13/a_27_368#
+ sky130_fd_sc_hs__einvp_4_13/a_473_323# sky130_fd_sc_hs__einvp_4
Xsky130_fd_sc_hs__dlygate4sd3_1_20 DVSS DVDD DVSS DVDD sky130_fd_sc_hs__dlygate4sd3_1_20/A
+ sky130_fd_sc_hs__dlygate4sd3_1_9/A sky130_fd_sc_hs__dlygate4sd3_1_20/a_405_138#
+ sky130_fd_sc_hs__dlygate4sd3_1_20/a_28_74# sky130_fd_sc_hs__dlygate4sd3_1_20/a_289_74#
+ sky130_fd_sc_hs__dlygate4sd3_1
Xsky130_fd_sc_hs__dlygate4sd3_1_42 DVSS DVDD DVSS DVDD sky130_fd_sc_hs__dlygate4sd3_1_75/X
+ sky130_fd_sc_hs__dlygate4sd3_1_43/X sky130_fd_sc_hs__dlygate4sd3_1_43/a_405_138#
+ sky130_fd_sc_hs__dlygate4sd3_1_43/a_28_74# sky130_fd_sc_hs__dlygate4sd3_1_43/a_289_74#
+ sky130_fd_sc_hs__dlygate4sd3_1
Xsky130_fd_sc_hs__dlygate4sd3_1_31 DVSS DVDD DVSS DVDD sky130_fd_sc_hs__dlygate4sd3_1_43/X
+ sky130_fd_sc_hs__dlygate4sd3_1_31/X sky130_fd_sc_hs__dlygate4sd3_1_31/a_405_138#
+ sky130_fd_sc_hs__dlygate4sd3_1_31/a_28_74# sky130_fd_sc_hs__dlygate4sd3_1_31/a_289_74#
+ sky130_fd_sc_hs__dlygate4sd3_1
Xsky130_fd_sc_hs__dlygate4sd3_1_53 DVSS DVDD DVSS DVDD sky130_fd_sc_hs__dlygate4sd3_1_53/A
+ sky130_fd_sc_hs__dlygate4sd3_1_53/X sky130_fd_sc_hs__dlygate4sd3_1_53/a_405_138#
+ sky130_fd_sc_hs__dlygate4sd3_1_53/a_28_74# sky130_fd_sc_hs__dlygate4sd3_1_53/a_289_74#
+ sky130_fd_sc_hs__dlygate4sd3_1
Xsky130_fd_sc_hs__dlygate4sd3_1_64 DVSS DVDD DVSS DVDD sky130_fd_sc_hs__dlygate4sd2_1_1/X
+ sky130_fd_sc_hs__dlygate4sd3_1_65/X sky130_fd_sc_hs__dlygate4sd3_1_65/a_405_138#
+ sky130_fd_sc_hs__dlygate4sd3_1_65/a_28_74# sky130_fd_sc_hs__dlygate4sd3_1_65/a_289_74#
+ sky130_fd_sc_hs__dlygate4sd3_1
Xsky130_fd_sc_hs__dlygate4sd3_1_75 DVSS DVDD DVSS DVDD sky130_fd_sc_hs__dlygate4sd3_1_75/A
+ sky130_fd_sc_hs__dlygate4sd3_1_75/X sky130_fd_sc_hs__dlygate4sd3_1_75/a_405_138#
+ sky130_fd_sc_hs__dlygate4sd3_1_75/a_28_74# sky130_fd_sc_hs__dlygate4sd3_1_75/a_289_74#
+ sky130_fd_sc_hs__dlygate4sd3_1
Xsky130_fd_sc_hs__nand2_4_3 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_4_3/Y delay_con_msb[3]
+ osc_000 sky130_fd_sc_hs__nand2_4_3/a_27_74# sky130_fd_sc_hs__nand2_4
Xsky130_fd_sc_hs__nand2_2_102 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_2_102/Y sky130_fd_sc_hs__nand2_2_99/B
+ osc_036 sky130_fd_sc_hs__nand2_2_102/a_27_74# sky130_fd_sc_hs__nand2_2
Xsky130_fd_sc_hs__einvp_8_4 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_8_3/A pi2_l[3]
+ sky130_fd_sc_hs__inv_4_7/Y sky130_fd_sc_hs__einvp_8_5/a_802_323# sky130_fd_sc_hs__einvp_8_5/a_27_74#
+ sky130_fd_sc_hs__einvp_8_5/a_27_368# sky130_fd_sc_hs__einvp_8
Xsky130_fd_sc_hs__inv_16_20 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__and4_2_3/A sky130_fd_sc_hs__inv_16_31/A
+ sky130_fd_sc_hs__inv_16
Xsky130_fd_sc_hs__inv_16_31 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__and4_2_3/D sky130_fd_sc_hs__inv_16_31/A
+ sky130_fd_sc_hs__inv_16
Xsky130_fd_sc_hs__nand2_2_0 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_2_1/Y sky130_fd_sc_hs__nand2_2_9/B
+ osc_000 sky130_fd_sc_hs__nand2_2_1/a_27_74# sky130_fd_sc_hs__nand2_2
Xsky130_fd_sc_hs__einvp_1_13 DVSS DVDD DVDD DVSS pi1_l[0] sky130_fd_sc_hs__inv_8_7/A
+ sky130_fd_sc_hs__inv_4_15/Y sky130_fd_sc_hs__einvp_1_13/a_44_549# sky130_fd_sc_hs__einvp_1_13/a_318_74#
+ sky130_fd_sc_hs__einvp_1_13/a_310_392# sky130_fd_sc_hs__einvp_1
Xsky130_fd_sc_hs__inv_8_9 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_8_9/A p5 sky130_fd_sc_hs__inv_8
Xsky130_fd_sc_hs__nand2_4_30 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_4_31/Y delay_con_msb[2]
+ osc_000 sky130_fd_sc_hs__nand2_4_31/a_27_74# sky130_fd_sc_hs__nand2_4
Xsky130_fd_sc_hs__nand2_4_41 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_4_41/Y delay_con_msb[3]
+ osc_000 sky130_fd_sc_hs__nand2_4_41/a_27_74# sky130_fd_sc_hs__nand2_4
Xsky130_fd_sc_hs__nand2_4_52 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_4_53/Y delay_con_msb[1]
+ osc_000 sky130_fd_sc_hs__nand2_4_53/a_27_74# sky130_fd_sc_hs__nand2_4
Xsky130_fd_sc_hs__nand2_4_63 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_4_63/Y delay_con_msb[0]
+ osc_144 sky130_fd_sc_hs__nand2_4_63/a_27_74# sky130_fd_sc_hs__nand2_4
Xsky130_fd_sc_hs__nand2_4_74 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_4_75/Y delay_con_msb[0]
+ osc_108 sky130_fd_sc_hs__nand2_4_75/a_27_74# sky130_fd_sc_hs__nand2_4
Xsky130_fd_sc_hs__nand2_4_85 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_4_85/Y delay_con_msb[0]
+ osc_108 sky130_fd_sc_hs__nand2_4_85/a_27_74# sky130_fd_sc_hs__nand2_4
Xsky130_fd_sc_hs__nand2_4_96 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_4_97/Y delay_con_msb[0]
+ osc_072 sky130_fd_sc_hs__nand2_4_97/a_27_74# sky130_fd_sc_hs__nand2_4
Xsky130_fd_sc_hs__clkbuf_4_1 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__clkbuf_4_1/A sky130_fd_sc_hs__nand2_8_9/B
+ sky130_fd_sc_hs__clkbuf_4_1/a_83_270# sky130_fd_sc_hs__clkbuf_4
Xsky130_fd_sc_hs__inv_4_3 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_3/Y osc_072 sky130_fd_sc_hs__inv_4
Xsky130_fd_sc_hs__einvp_4_13 DVSS DVDD DVDD DVSS pi1_l[2] sky130_fd_sc_hs__inv_8_7/A
+ sky130_fd_sc_hs__inv_4_15/Y sky130_fd_sc_hs__einvp_4_13/a_27_74# sky130_fd_sc_hs__einvp_4_13/a_27_368#
+ sky130_fd_sc_hs__einvp_4_13/a_473_323# sky130_fd_sc_hs__einvp_4
Xsky130_fd_sc_hs__dlygate4sd3_1_10 DVSS DVDD DVSS DVDD sky130_fd_sc_hs__dlygate4sd3_1_25/X
+ sky130_fd_sc_hs__dlygate4sd3_1_5/A sky130_fd_sc_hs__dlygate4sd3_1_11/a_405_138#
+ sky130_fd_sc_hs__dlygate4sd3_1_11/a_28_74# sky130_fd_sc_hs__dlygate4sd3_1_11/a_289_74#
+ sky130_fd_sc_hs__dlygate4sd3_1
Xsky130_fd_sc_hs__dlygate4sd3_1_21 DVSS DVDD DVSS DVDD sky130_fd_sc_hs__dlygate4sd3_1_1/X
+ sky130_fd_sc_hs__dlygate4sd3_1_3/A sky130_fd_sc_hs__dlygate4sd3_1_21/a_405_138#
+ sky130_fd_sc_hs__dlygate4sd3_1_21/a_28_74# sky130_fd_sc_hs__dlygate4sd3_1_21/a_289_74#
+ sky130_fd_sc_hs__dlygate4sd3_1
Xsky130_fd_sc_hs__dlygate4sd3_1_43 DVSS DVDD DVSS DVDD sky130_fd_sc_hs__dlygate4sd3_1_75/X
+ sky130_fd_sc_hs__dlygate4sd3_1_43/X sky130_fd_sc_hs__dlygate4sd3_1_43/a_405_138#
+ sky130_fd_sc_hs__dlygate4sd3_1_43/a_28_74# sky130_fd_sc_hs__dlygate4sd3_1_43/a_289_74#
+ sky130_fd_sc_hs__dlygate4sd3_1
Xsky130_fd_sc_hs__dlygate4sd3_1_54 DVSS DVDD DVSS DVDD sky130_fd_sc_hs__dlygate4sd3_1_56/A
+ sky130_fd_sc_hs__dlygate4sd3_1_63/A sky130_fd_sc_hs__dlygate4sd3_1_56/a_405_138#
+ sky130_fd_sc_hs__dlygate4sd3_1_56/a_28_74# sky130_fd_sc_hs__dlygate4sd3_1_56/a_289_74#
+ sky130_fd_sc_hs__dlygate4sd3_1
Xsky130_fd_sc_hs__dlygate4sd3_1_65 DVSS DVDD DVSS DVDD sky130_fd_sc_hs__dlygate4sd2_1_1/X
+ sky130_fd_sc_hs__dlygate4sd3_1_65/X sky130_fd_sc_hs__dlygate4sd3_1_65/a_405_138#
+ sky130_fd_sc_hs__dlygate4sd3_1_65/a_28_74# sky130_fd_sc_hs__dlygate4sd3_1_65/a_289_74#
+ sky130_fd_sc_hs__dlygate4sd3_1
Xsky130_fd_sc_hs__dlygate4sd3_1_76 DVSS DVDD DVSS DVDD sky130_fd_sc_hs__dlygate4sd3_1_79/X
+ sky130_fd_sc_hs__dlygate4sd3_1_78/X sky130_fd_sc_hs__dlygate4sd3_1_78/a_405_138#
+ sky130_fd_sc_hs__dlygate4sd3_1_78/a_28_74# sky130_fd_sc_hs__dlygate4sd3_1_78/a_289_74#
+ sky130_fd_sc_hs__dlygate4sd3_1
Xsky130_fd_sc_hs__dlygate4sd3_1_32 DVSS DVDD DVSS DVDD sky130_fd_sc_hs__dlygate4sd3_1_33/A
+ sky130_fd_sc_hs__dlygate4sd3_1_45/A sky130_fd_sc_hs__dlygate4sd3_1_33/a_405_138#
+ sky130_fd_sc_hs__dlygate4sd3_1_33/a_28_74# sky130_fd_sc_hs__dlygate4sd3_1_33/a_289_74#
+ sky130_fd_sc_hs__dlygate4sd3_1
Xsky130_fd_sc_hs__nand2_4_4 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_4_5/Y delay_con_msb[3]
+ osc_144 sky130_fd_sc_hs__nand2_4_5/a_27_74# sky130_fd_sc_hs__nand2_4
Xsky130_fd_sc_hs__nand2_2_103 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_2_103/Y sky130_fd_sc_hs__nand2_2_99/B
+ osc_036 sky130_fd_sc_hs__nand2_2_103/a_27_74# sky130_fd_sc_hs__nand2_2
Xsky130_fd_sc_hs__einvp_8_5 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_8_3/A pi2_l[3]
+ sky130_fd_sc_hs__inv_4_7/Y sky130_fd_sc_hs__einvp_8_5/a_802_323# sky130_fd_sc_hs__einvp_8_5/a_27_74#
+ sky130_fd_sc_hs__einvp_8_5/a_27_368# sky130_fd_sc_hs__einvp_8
Xsky130_fd_sc_hs__inv_16_10 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__and4_2_5/B sky130_fd_sc_hs__inv_16_7/Y
+ sky130_fd_sc_hs__inv_16
Xsky130_fd_sc_hs__inv_16_21 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__and4_2_3/A sky130_fd_sc_hs__inv_16_31/A
+ sky130_fd_sc_hs__inv_16
Xsky130_fd_sc_hs__nand2_2_1 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_2_1/Y sky130_fd_sc_hs__nand2_2_9/B
+ osc_000 sky130_fd_sc_hs__nand2_2_1/a_27_74# sky130_fd_sc_hs__nand2_2
Xsky130_fd_sc_hs__einvp_1_14 DVSS DVDD DVDD DVSS pi1_r[0] sky130_fd_sc_hs__inv_8_7/A
+ sky130_fd_sc_hs__inv_4_17/Y sky130_fd_sc_hs__einvp_1_15/a_44_549# sky130_fd_sc_hs__einvp_1_15/a_318_74#
+ sky130_fd_sc_hs__einvp_1_15/a_310_392# sky130_fd_sc_hs__einvp_1
Xsky130_fd_sc_hs__nand2_4_20 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_4_21/Y delay_con_msb[1]
+ osc_144 sky130_fd_sc_hs__nand2_4_21/a_27_74# sky130_fd_sc_hs__nand2_4
Xsky130_fd_sc_hs__nand2_4_31 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_4_31/Y delay_con_msb[2]
+ osc_000 sky130_fd_sc_hs__nand2_4_31/a_27_74# sky130_fd_sc_hs__nand2_4
Xsky130_fd_sc_hs__nand2_4_42 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_4_43/Y delay_con_msb[3]
+ osc_144 sky130_fd_sc_hs__nand2_4_43/a_27_74# sky130_fd_sc_hs__nand2_4
Xsky130_fd_sc_hs__nand2_4_53 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_4_53/Y delay_con_msb[1]
+ osc_000 sky130_fd_sc_hs__nand2_4_53/a_27_74# sky130_fd_sc_hs__nand2_4
Xsky130_fd_sc_hs__nand2_4_64 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_4_65/Y delay_con_msb[0]
+ osc_000 sky130_fd_sc_hs__nand2_4_65/a_27_74# sky130_fd_sc_hs__nand2_4
Xsky130_fd_sc_hs__nand2_4_75 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_4_75/Y delay_con_msb[0]
+ osc_108 sky130_fd_sc_hs__nand2_4_75/a_27_74# sky130_fd_sc_hs__nand2_4
Xsky130_fd_sc_hs__nand2_4_86 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_4_87/Y delay_con_msb[0]
+ osc_108 sky130_fd_sc_hs__nand2_4_87/a_27_74# sky130_fd_sc_hs__nand2_4
Xsky130_fd_sc_hs__nand2_4_97 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_4_97/Y delay_con_msb[0]
+ osc_072 sky130_fd_sc_hs__nand2_4_97/a_27_74# sky130_fd_sc_hs__nand2_4
Xsky130_fd_sc_hs__clkbuf_4_2 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__clkbuf_4_3/A sky130_fd_sc_hs__clkbuf_4_3/X
+ sky130_fd_sc_hs__clkbuf_4_3/a_83_270# sky130_fd_sc_hs__clkbuf_4
Xsky130_fd_sc_hs__inv_4_4 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_5/Y osc_108 sky130_fd_sc_hs__inv_4
Xsky130_fd_sc_hs__clkbuf_2_10 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__buf_4_1/A sky130_fd_sc_hs__clkbuf_2_8/A
+ sky130_fd_sc_hs__clkbuf_2_8/a_43_192# sky130_fd_sc_hs__clkbuf_2
Xsky130_fd_sc_hs__einvp_4_14 DVSS DVDD DVDD DVSS pi1_r[2] sky130_fd_sc_hs__inv_8_7/A
+ sky130_fd_sc_hs__inv_4_17/Y sky130_fd_sc_hs__einvp_4_15/a_27_74# sky130_fd_sc_hs__einvp_4_15/a_27_368#
+ sky130_fd_sc_hs__einvp_4_15/a_473_323# sky130_fd_sc_hs__einvp_4
Xsky130_fd_sc_hs__dlygate4sd3_1_11 DVSS DVDD DVSS DVDD sky130_fd_sc_hs__dlygate4sd3_1_25/X
+ sky130_fd_sc_hs__dlygate4sd3_1_5/A sky130_fd_sc_hs__dlygate4sd3_1_11/a_405_138#
+ sky130_fd_sc_hs__dlygate4sd3_1_11/a_28_74# sky130_fd_sc_hs__dlygate4sd3_1_11/a_289_74#
+ sky130_fd_sc_hs__dlygate4sd3_1
Xsky130_fd_sc_hs__dlygate4sd3_1_22 DVSS DVDD DVSS DVDD sky130_fd_sc_hs__inv_16_13/Y
+ sky130_fd_sc_hs__clkbuf_2_1/A sky130_fd_sc_hs__dlygate4sd3_1_23/a_405_138# sky130_fd_sc_hs__dlygate4sd3_1_23/a_28_74#
+ sky130_fd_sc_hs__dlygate4sd3_1_23/a_289_74# sky130_fd_sc_hs__dlygate4sd3_1
Xsky130_fd_sc_hs__dlygate4sd3_1_44 DVSS DVDD DVSS DVDD sky130_fd_sc_hs__dlygate4sd3_1_45/A
+ sky130_fd_sc_hs__dlygate4sd3_1_79/A sky130_fd_sc_hs__dlygate4sd3_1_45/a_405_138#
+ sky130_fd_sc_hs__dlygate4sd3_1_45/a_28_74# sky130_fd_sc_hs__dlygate4sd3_1_45/a_289_74#
+ sky130_fd_sc_hs__dlygate4sd3_1
Xsky130_fd_sc_hs__dlygate4sd3_1_55 DVSS DVDD DVSS DVDD sky130_fd_sc_hs__dlygate4sd3_1_62/X
+ sky130_fd_sc_hs__dlygate4sd3_1_57/X sky130_fd_sc_hs__dlygate4sd3_1_57/a_405_138#
+ sky130_fd_sc_hs__dlygate4sd3_1_57/a_28_74# sky130_fd_sc_hs__dlygate4sd3_1_57/a_289_74#
+ sky130_fd_sc_hs__dlygate4sd3_1
Xsky130_fd_sc_hs__dlygate4sd3_1_66 DVSS DVDD DVSS DVDD sky130_fd_sc_hs__dlygate4sd3_1_68/A
+ sky130_fd_sc_hs__dlygate4sd3_1_68/X sky130_fd_sc_hs__dlygate4sd3_1_68/a_405_138#
+ sky130_fd_sc_hs__dlygate4sd3_1_68/a_28_74# sky130_fd_sc_hs__dlygate4sd3_1_68/a_289_74#
+ sky130_fd_sc_hs__dlygate4sd3_1
Xsky130_fd_sc_hs__dlygate4sd3_1_77 DVSS DVDD DVSS DVDD sky130_fd_sc_hs__dlygate4sd3_1_79/A
+ sky130_fd_sc_hs__dlygate4sd3_1_79/X sky130_fd_sc_hs__dlygate4sd3_1_79/a_405_138#
+ sky130_fd_sc_hs__dlygate4sd3_1_79/a_28_74# sky130_fd_sc_hs__dlygate4sd3_1_79/a_289_74#
+ sky130_fd_sc_hs__dlygate4sd3_1
Xsky130_fd_sc_hs__dlygate4sd3_1_33 DVSS DVDD DVSS DVDD sky130_fd_sc_hs__dlygate4sd3_1_33/A
+ sky130_fd_sc_hs__dlygate4sd3_1_45/A sky130_fd_sc_hs__dlygate4sd3_1_33/a_405_138#
+ sky130_fd_sc_hs__dlygate4sd3_1_33/a_28_74# sky130_fd_sc_hs__dlygate4sd3_1_33/a_289_74#
+ sky130_fd_sc_hs__dlygate4sd3_1
Xsky130_fd_sc_hs__nand2_4_5 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_4_5/Y delay_con_msb[3]
+ osc_144 sky130_fd_sc_hs__nand2_4_5/a_27_74# sky130_fd_sc_hs__nand2_4
Xsky130_fd_sc_hs__nand2_2_104 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_2_105/Y sky130_fd_sc_hs__a21oi_1_45/Y
+ osc_036 sky130_fd_sc_hs__nand2_2_105/a_27_74# sky130_fd_sc_hs__nand2_2
Xsky130_fd_sc_hs__einvp_8_6 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_8_3/A pi2_r[3]
+ sky130_fd_sc_hs__inv_4_9/Y sky130_fd_sc_hs__einvp_8_7/a_802_323# sky130_fd_sc_hs__einvp_8_7/a_27_74#
+ sky130_fd_sc_hs__einvp_8_7/a_27_368# sky130_fd_sc_hs__einvp_8
Xsky130_fd_sc_hs__inv_16_11 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__and4_2_5/B sky130_fd_sc_hs__inv_16_7/Y
+ sky130_fd_sc_hs__inv_16
Xsky130_fd_sc_hs__inv_16_22 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__and4_2_5/C sky130_fd_sc_hs__inv_16_7/Y
+ sky130_fd_sc_hs__inv_16
Xsky130_fd_sc_hs__nand2_2_2 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_2_3/Y sky130_fd_sc_hs__nand2_2_5/B
+ osc_000 sky130_fd_sc_hs__nand2_2_3/a_27_74# sky130_fd_sc_hs__nand2_2
Xsky130_fd_sc_hs__einvp_1_15 DVSS DVDD DVDD DVSS pi1_r[0] sky130_fd_sc_hs__inv_8_7/A
+ sky130_fd_sc_hs__inv_4_17/Y sky130_fd_sc_hs__einvp_1_15/a_44_549# sky130_fd_sc_hs__einvp_1_15/a_318_74#
+ sky130_fd_sc_hs__einvp_1_15/a_310_392# sky130_fd_sc_hs__einvp_1
Xsky130_fd_sc_hs__nand2_4_10 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_4_11/Y delay_con_msb[3]
+ osc_000 sky130_fd_sc_hs__nand2_4_11/a_27_74# sky130_fd_sc_hs__nand2_4
Xsky130_fd_sc_hs__nand2_4_21 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_4_21/Y delay_con_msb[1]
+ osc_144 sky130_fd_sc_hs__nand2_4_21/a_27_74# sky130_fd_sc_hs__nand2_4
Xsky130_fd_sc_hs__nand2_4_32 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_4_33/Y delay_con_msb[1]
+ osc_144 sky130_fd_sc_hs__nand2_4_33/a_27_74# sky130_fd_sc_hs__nand2_4
Xsky130_fd_sc_hs__nand2_4_43 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_4_43/Y delay_con_msb[3]
+ osc_144 sky130_fd_sc_hs__nand2_4_43/a_27_74# sky130_fd_sc_hs__nand2_4
Xsky130_fd_sc_hs__nand2_4_54 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_4_55/Y delay_con_msb[0]
+ osc_000 sky130_fd_sc_hs__nand2_4_55/a_27_74# sky130_fd_sc_hs__nand2_4
Xsky130_fd_sc_hs__nand2_4_65 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_4_65/Y delay_con_msb[0]
+ osc_000 sky130_fd_sc_hs__nand2_4_65/a_27_74# sky130_fd_sc_hs__nand2_4
Xsky130_fd_sc_hs__nand2_4_76 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_4_77/Y delay_con_msb[0]
+ osc_144 sky130_fd_sc_hs__nand2_4_77/a_27_74# sky130_fd_sc_hs__nand2_4
Xsky130_fd_sc_hs__nand2_4_87 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_4_87/Y delay_con_msb[0]
+ osc_108 sky130_fd_sc_hs__nand2_4_87/a_27_74# sky130_fd_sc_hs__nand2_4
Xsky130_fd_sc_hs__nand2_4_98 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_4_99/Y delay_con_msb[0]
+ osc_072 sky130_fd_sc_hs__nand2_4_99/a_27_74# sky130_fd_sc_hs__nand2_4
Xsky130_fd_sc_hs__einvp_4_0 DVSS DVDD DVDD DVSS pi3_l[2] sky130_fd_sc_hs__inv_8_1/A
+ sky130_fd_sc_hs__inv_4_3/Y sky130_fd_sc_hs__einvp_4_1/a_27_74# sky130_fd_sc_hs__einvp_4_1/a_27_368#
+ sky130_fd_sc_hs__einvp_4_1/a_473_323# sky130_fd_sc_hs__einvp_4
Xsky130_fd_sc_hs__clkbuf_4_3 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__clkbuf_4_3/A sky130_fd_sc_hs__clkbuf_4_3/X
+ sky130_fd_sc_hs__clkbuf_4_3/a_83_270# sky130_fd_sc_hs__clkbuf_4
Xsky130_fd_sc_hs__inv_4_5 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_5/Y osc_108 sky130_fd_sc_hs__inv_4
Xsky130_fd_sc_hs__clkbuf_2_0 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__clkbuf_2_1/X sky130_fd_sc_hs__clkbuf_2_1/A
+ sky130_fd_sc_hs__clkbuf_2_1/a_43_192# sky130_fd_sc_hs__clkbuf_2
Xsky130_fd_sc_hs__clkbuf_2_11 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__clkbuf_4_5/A sky130_fd_sc_hs__clkbuf_2_9/A
+ sky130_fd_sc_hs__clkbuf_2_9/a_43_192# sky130_fd_sc_hs__clkbuf_2
Xsky130_fd_sc_hs__einvp_4_15 DVSS DVDD DVDD DVSS pi1_r[2] sky130_fd_sc_hs__inv_8_7/A
+ sky130_fd_sc_hs__inv_4_17/Y sky130_fd_sc_hs__einvp_4_15/a_27_74# sky130_fd_sc_hs__einvp_4_15/a_27_368#
+ sky130_fd_sc_hs__einvp_4_15/a_473_323# sky130_fd_sc_hs__einvp_4
Xsky130_fd_sc_hs__dlygate4sd3_1_12 DVSS DVDD DVSS DVDD sky130_fd_sc_hs__dlygate4sd3_1_9/X
+ sky130_fd_sc_hs__clkbuf_1_1/A sky130_fd_sc_hs__dlygate4sd3_1_14/a_405_138# sky130_fd_sc_hs__dlygate4sd3_1_14/a_28_74#
+ sky130_fd_sc_hs__dlygate4sd3_1_14/a_289_74# sky130_fd_sc_hs__dlygate4sd3_1
Xsky130_fd_sc_hs__dlygate4sd3_1_23 DVSS DVDD DVSS DVDD sky130_fd_sc_hs__inv_16_13/Y
+ sky130_fd_sc_hs__clkbuf_2_1/A sky130_fd_sc_hs__dlygate4sd3_1_23/a_405_138# sky130_fd_sc_hs__dlygate4sd3_1_23/a_28_74#
+ sky130_fd_sc_hs__dlygate4sd3_1_23/a_289_74# sky130_fd_sc_hs__dlygate4sd3_1
Xsky130_fd_sc_hs__dlygate4sd3_1_34 DVSS DVDD DVSS DVDD sky130_fd_sc_hs__dlygate4sd3_1_53/X
+ sky130_fd_sc_hs__dlygate4sd3_1_35/X sky130_fd_sc_hs__dlygate4sd3_1_35/a_405_138#
+ sky130_fd_sc_hs__dlygate4sd3_1_35/a_28_74# sky130_fd_sc_hs__dlygate4sd3_1_35/a_289_74#
+ sky130_fd_sc_hs__dlygate4sd3_1
Xsky130_fd_sc_hs__dlygate4sd3_1_45 DVSS DVDD DVSS DVDD sky130_fd_sc_hs__dlygate4sd3_1_45/A
+ sky130_fd_sc_hs__dlygate4sd3_1_79/A sky130_fd_sc_hs__dlygate4sd3_1_45/a_405_138#
+ sky130_fd_sc_hs__dlygate4sd3_1_45/a_28_74# sky130_fd_sc_hs__dlygate4sd3_1_45/a_289_74#
+ sky130_fd_sc_hs__dlygate4sd3_1
Xsky130_fd_sc_hs__dlygate4sd3_1_56 DVSS DVDD DVSS DVDD sky130_fd_sc_hs__dlygate4sd3_1_56/A
+ sky130_fd_sc_hs__dlygate4sd3_1_63/A sky130_fd_sc_hs__dlygate4sd3_1_56/a_405_138#
+ sky130_fd_sc_hs__dlygate4sd3_1_56/a_28_74# sky130_fd_sc_hs__dlygate4sd3_1_56/a_289_74#
+ sky130_fd_sc_hs__dlygate4sd3_1
Xsky130_fd_sc_hs__dlygate4sd3_1_67 DVSS DVDD DVSS DVDD sky130_fd_sc_hs__dlygate4sd3_1_71/X
+ sky130_fd_sc_hs__dlygate4sd2_1_1/A sky130_fd_sc_hs__dlygate4sd3_1_69/a_405_138#
+ sky130_fd_sc_hs__dlygate4sd3_1_69/a_28_74# sky130_fd_sc_hs__dlygate4sd3_1_69/a_289_74#
+ sky130_fd_sc_hs__dlygate4sd3_1
Xsky130_fd_sc_hs__dlygate4sd3_1_78 DVSS DVDD DVSS DVDD sky130_fd_sc_hs__dlygate4sd3_1_79/X
+ sky130_fd_sc_hs__dlygate4sd3_1_78/X sky130_fd_sc_hs__dlygate4sd3_1_78/a_405_138#
+ sky130_fd_sc_hs__dlygate4sd3_1_78/a_28_74# sky130_fd_sc_hs__dlygate4sd3_1_78/a_289_74#
+ sky130_fd_sc_hs__dlygate4sd3_1
Xsky130_fd_sc_hs__nand2_4_6 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_4_7/Y delay_con_msb[3]
+ osc_000 sky130_fd_sc_hs__nand2_4_7/a_27_74# sky130_fd_sc_hs__nand2_4
Xsky130_fd_sc_hs__nand2_2_105 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_2_105/Y sky130_fd_sc_hs__a21oi_1_45/Y
+ osc_036 sky130_fd_sc_hs__nand2_2_105/a_27_74# sky130_fd_sc_hs__nand2_2
Xsky130_fd_sc_hs__einvp_8_7 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_8_3/A pi2_r[3]
+ sky130_fd_sc_hs__inv_4_9/Y sky130_fd_sc_hs__einvp_8_7/a_802_323# sky130_fd_sc_hs__einvp_8_7/a_27_74#
+ sky130_fd_sc_hs__einvp_8_7/a_27_368# sky130_fd_sc_hs__einvp_8
Xsky130_fd_sc_hs__inv_16_12 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_16_13/Y sky130_fd_sc_hs__and2_2_3/X
+ sky130_fd_sc_hs__inv_16
Xsky130_fd_sc_hs__inv_16_23 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__and4_2_5/C sky130_fd_sc_hs__inv_16_7/Y
+ sky130_fd_sc_hs__inv_16
Xsky130_fd_sc_hs__nand2_2_3 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_2_3/Y sky130_fd_sc_hs__nand2_2_5/B
+ osc_000 sky130_fd_sc_hs__nand2_2_3/a_27_74# sky130_fd_sc_hs__nand2_2
Xsky130_fd_sc_hs__einvp_1_16 DVSS DVDD DVDD DVSS pi5_l[0] sky130_fd_sc_hs__inv_8_9/A
+ sky130_fd_sc_hs__inv_4_19/Y sky130_fd_sc_hs__einvp_1_17/a_44_549# sky130_fd_sc_hs__einvp_1_17/a_318_74#
+ sky130_fd_sc_hs__einvp_1_17/a_310_392# sky130_fd_sc_hs__einvp_1
Xsky130_fd_sc_hs__nand2_4_11 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_4_11/Y delay_con_msb[3]
+ osc_000 sky130_fd_sc_hs__nand2_4_11/a_27_74# sky130_fd_sc_hs__nand2_4
Xsky130_fd_sc_hs__nand2_4_22 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_4_23/Y delay_con_msb[3]
+ osc_144 sky130_fd_sc_hs__nand2_4_23/a_27_74# sky130_fd_sc_hs__nand2_4
Xsky130_fd_sc_hs__nand2_4_33 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_4_33/Y delay_con_msb[1]
+ osc_144 sky130_fd_sc_hs__nand2_4_33/a_27_74# sky130_fd_sc_hs__nand2_4
Xsky130_fd_sc_hs__nand2_4_44 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_4_45/Y delay_con_msb[1]
+ osc_000 sky130_fd_sc_hs__nand2_4_45/a_27_74# sky130_fd_sc_hs__nand2_4
Xsky130_fd_sc_hs__nand2_4_55 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_4_55/Y delay_con_msb[0]
+ osc_000 sky130_fd_sc_hs__nand2_4_55/a_27_74# sky130_fd_sc_hs__nand2_4
Xsky130_fd_sc_hs__nand2_4_66 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_4_67/Y delay_con_msb[3]
+ osc_108 sky130_fd_sc_hs__nand2_4_67/a_27_74# sky130_fd_sc_hs__nand2_4
Xsky130_fd_sc_hs__nand2_4_77 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_4_77/Y delay_con_msb[0]
+ osc_144 sky130_fd_sc_hs__nand2_4_77/a_27_74# sky130_fd_sc_hs__nand2_4
Xsky130_fd_sc_hs__nand2_4_88 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_4_89/Y delay_con_msb[0]
+ osc_108 sky130_fd_sc_hs__nand2_4_89/a_27_74# sky130_fd_sc_hs__nand2_4
Xsky130_fd_sc_hs__nand2_4_99 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_4_99/Y delay_con_msb[0]
+ osc_072 sky130_fd_sc_hs__nand2_4_99/a_27_74# sky130_fd_sc_hs__nand2_4
Xsky130_fd_sc_hs__einvp_4_1 DVSS DVDD DVDD DVSS pi3_l[2] sky130_fd_sc_hs__inv_8_1/A
+ sky130_fd_sc_hs__inv_4_3/Y sky130_fd_sc_hs__einvp_4_1/a_27_74# sky130_fd_sc_hs__einvp_4_1/a_27_368#
+ sky130_fd_sc_hs__einvp_4_1/a_473_323# sky130_fd_sc_hs__einvp_4
Xsky130_fd_sc_hs__clkbuf_4_4 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__clkbuf_4_5/A sky130_fd_sc_hs__clkbuf_4_5/X
+ sky130_fd_sc_hs__clkbuf_4_5/a_83_270# sky130_fd_sc_hs__clkbuf_4
Xsky130_fd_sc_hs__inv_4_6 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_7/Y osc_036 sky130_fd_sc_hs__inv_4
Xsky130_fd_sc_hs__clkbuf_2_1 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__clkbuf_2_1/X sky130_fd_sc_hs__clkbuf_2_1/A
+ sky130_fd_sc_hs__clkbuf_2_1/a_43_192# sky130_fd_sc_hs__clkbuf_2
Xsky130_fd_sc_hs__clkbuf_2_12 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__clkbuf_2_8/A sky130_fd_sc_hs__clkbuf_4_5/X
+ sky130_fd_sc_hs__clkbuf_2_14/a_43_192# sky130_fd_sc_hs__clkbuf_2
Xsky130_fd_sc_hs__einvp_4_16 DVSS DVDD DVDD DVSS pi5_l[2] sky130_fd_sc_hs__inv_8_9/A
+ sky130_fd_sc_hs__inv_4_19/Y sky130_fd_sc_hs__einvp_4_17/a_27_74# sky130_fd_sc_hs__einvp_4_17/a_27_368#
+ sky130_fd_sc_hs__einvp_4_17/a_473_323# sky130_fd_sc_hs__einvp_4
Xsky130_fd_sc_hs__dlygate4sd3_1_13 DVSS DVDD DVSS DVDD sky130_fd_sc_hs__dlygate4sd3_1_7/X
+ sky130_fd_sc_hs__dlygate4sd3_1_20/A sky130_fd_sc_hs__dlygate4sd3_1_15/a_405_138#
+ sky130_fd_sc_hs__dlygate4sd3_1_15/a_28_74# sky130_fd_sc_hs__dlygate4sd3_1_15/a_289_74#
+ sky130_fd_sc_hs__dlygate4sd3_1
Xsky130_fd_sc_hs__dlygate4sd3_1_24 DVSS DVDD DVSS DVDD sky130_fd_sc_hs__dlygate4sd3_1_3/X
+ sky130_fd_sc_hs__dlygate4sd3_1_25/X sky130_fd_sc_hs__dlygate4sd3_1_25/a_405_138#
+ sky130_fd_sc_hs__dlygate4sd3_1_25/a_28_74# sky130_fd_sc_hs__dlygate4sd3_1_25/a_289_74#
+ sky130_fd_sc_hs__dlygate4sd3_1
Xsky130_fd_sc_hs__dlygate4sd3_1_35 DVSS DVDD DVSS DVDD sky130_fd_sc_hs__dlygate4sd3_1_53/X
+ sky130_fd_sc_hs__dlygate4sd3_1_35/X sky130_fd_sc_hs__dlygate4sd3_1_35/a_405_138#
+ sky130_fd_sc_hs__dlygate4sd3_1_35/a_28_74# sky130_fd_sc_hs__dlygate4sd3_1_35/a_289_74#
+ sky130_fd_sc_hs__dlygate4sd3_1
Xsky130_fd_sc_hs__dlygate4sd3_1_46 DVSS DVDD DVSS DVDD sky130_fd_sc_hs__dlygate4sd3_1_49/X
+ sky130_fd_sc_hs__nand3_4_3/C sky130_fd_sc_hs__dlygate4sd3_1_47/a_405_138# sky130_fd_sc_hs__dlygate4sd3_1_47/a_28_74#
+ sky130_fd_sc_hs__dlygate4sd3_1_47/a_289_74# sky130_fd_sc_hs__dlygate4sd3_1
Xsky130_fd_sc_hs__dlygate4sd3_1_57 DVSS DVDD DVSS DVDD sky130_fd_sc_hs__dlygate4sd3_1_62/X
+ sky130_fd_sc_hs__dlygate4sd3_1_57/X sky130_fd_sc_hs__dlygate4sd3_1_57/a_405_138#
+ sky130_fd_sc_hs__dlygate4sd3_1_57/a_28_74# sky130_fd_sc_hs__dlygate4sd3_1_57/a_289_74#
+ sky130_fd_sc_hs__dlygate4sd3_1
Xsky130_fd_sc_hs__dlygate4sd3_1_68 DVSS DVDD DVSS DVDD sky130_fd_sc_hs__dlygate4sd3_1_68/A
+ sky130_fd_sc_hs__dlygate4sd3_1_68/X sky130_fd_sc_hs__dlygate4sd3_1_68/a_405_138#
+ sky130_fd_sc_hs__dlygate4sd3_1_68/a_28_74# sky130_fd_sc_hs__dlygate4sd3_1_68/a_289_74#
+ sky130_fd_sc_hs__dlygate4sd3_1
Xsky130_fd_sc_hs__dlygate4sd3_1_79 DVSS DVDD DVSS DVDD sky130_fd_sc_hs__dlygate4sd3_1_79/A
+ sky130_fd_sc_hs__dlygate4sd3_1_79/X sky130_fd_sc_hs__dlygate4sd3_1_79/a_405_138#
+ sky130_fd_sc_hs__dlygate4sd3_1_79/a_28_74# sky130_fd_sc_hs__dlygate4sd3_1_79/a_289_74#
+ sky130_fd_sc_hs__dlygate4sd3_1
Xsky130_fd_sc_hs__nand2_4_7 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_4_7/Y delay_con_msb[3]
+ osc_000 sky130_fd_sc_hs__nand2_4_7/a_27_74# sky130_fd_sc_hs__nand2_4
Xsky130_fd_sc_hs__nand2_2_106 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_2_108/Y sky130_fd_sc_hs__a21oi_1_49/Y
+ osc_036 sky130_fd_sc_hs__nand2_2_108/a_27_74# sky130_fd_sc_hs__nand2_2
Xsky130_fd_sc_hs__einvp_8_8 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_8_5/A pi4_l[3]
+ sky130_fd_sc_hs__inv_4_11/Y sky130_fd_sc_hs__einvp_8_8/a_802_323# sky130_fd_sc_hs__einvp_8_8/a_27_74#
+ sky130_fd_sc_hs__einvp_8_8/a_27_368# sky130_fd_sc_hs__einvp_8
Xsky130_fd_sc_hs__inv_16_13 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_16_13/Y sky130_fd_sc_hs__and2_2_3/X
+ sky130_fd_sc_hs__inv_16
Xsky130_fd_sc_hs__inv_16_24 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_16_31/A sky130_fd_sc_hs__inv_4_27/Y
+ sky130_fd_sc_hs__inv_16
Xsky130_fd_sc_hs__nand2_2_4 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_2_5/Y sky130_fd_sc_hs__nand2_2_5/B
+ osc_000 sky130_fd_sc_hs__nand2_2_5/a_27_74# sky130_fd_sc_hs__nand2_2
Xsky130_fd_sc_hs__einvp_1_17 DVSS DVDD DVDD DVSS pi5_l[0] sky130_fd_sc_hs__inv_8_9/A
+ sky130_fd_sc_hs__inv_4_19/Y sky130_fd_sc_hs__einvp_1_17/a_44_549# sky130_fd_sc_hs__einvp_1_17/a_318_74#
+ sky130_fd_sc_hs__einvp_1_17/a_310_392# sky130_fd_sc_hs__einvp_1
Xsky130_fd_sc_hs__nand2_4_12 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_4_13/Y delay_con_msb[2]
+ osc_144 sky130_fd_sc_hs__nand2_4_13/a_27_74# sky130_fd_sc_hs__nand2_4
Xsky130_fd_sc_hs__nand2_4_23 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_4_23/Y delay_con_msb[3]
+ osc_144 sky130_fd_sc_hs__nand2_4_23/a_27_74# sky130_fd_sc_hs__nand2_4
Xsky130_fd_sc_hs__nand2_4_34 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_4_35/Y delay_con_msb[2]
+ osc_144 sky130_fd_sc_hs__nand2_4_35/a_27_74# sky130_fd_sc_hs__nand2_4
Xsky130_fd_sc_hs__nand2_4_45 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_4_45/Y delay_con_msb[1]
+ osc_000 sky130_fd_sc_hs__nand2_4_45/a_27_74# sky130_fd_sc_hs__nand2_4
Xsky130_fd_sc_hs__nand2_4_56 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_4_57/Y delay_con_msb[0]
+ osc_000 sky130_fd_sc_hs__nand2_4_57/a_27_74# sky130_fd_sc_hs__nand2_4
Xsky130_fd_sc_hs__nand2_4_67 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_4_67/Y delay_con_msb[3]
+ osc_108 sky130_fd_sc_hs__nand2_4_67/a_27_74# sky130_fd_sc_hs__nand2_4
Xsky130_fd_sc_hs__nand2_4_78 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_4_79/Y delay_con_msb[1]
+ osc_108 sky130_fd_sc_hs__nand2_4_79/a_27_74# sky130_fd_sc_hs__nand2_4
Xsky130_fd_sc_hs__nand2_4_89 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_4_89/Y delay_con_msb[0]
+ osc_108 sky130_fd_sc_hs__nand2_4_89/a_27_74# sky130_fd_sc_hs__nand2_4
Xsky130_fd_sc_hs__einvp_4_2 DVSS DVDD DVDD DVSS pi3_r[2] sky130_fd_sc_hs__inv_8_1/A
+ sky130_fd_sc_hs__inv_4_5/Y sky130_fd_sc_hs__einvp_4_3/a_27_74# sky130_fd_sc_hs__einvp_4_3/a_27_368#
+ sky130_fd_sc_hs__einvp_4_3/a_473_323# sky130_fd_sc_hs__einvp_4
Xsky130_fd_sc_hs__clkbuf_4_5 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__clkbuf_4_5/A sky130_fd_sc_hs__clkbuf_4_5/X
+ sky130_fd_sc_hs__clkbuf_4_5/a_83_270# sky130_fd_sc_hs__clkbuf_4
Xsky130_fd_sc_hs__inv_4_7 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_7/Y osc_036 sky130_fd_sc_hs__inv_4
Xsky130_fd_sc_hs__clkbuf_2_13 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__clkbuf_2_17/A sky130_fd_sc_hs__buf_4_1/X
+ sky130_fd_sc_hs__clkbuf_2_15/a_43_192# sky130_fd_sc_hs__clkbuf_2
Xsky130_fd_sc_hs__clkbuf_2_2 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__clkbuf_4_3/A sky130_fd_sc_hs__clkbuf_2_3/A
+ sky130_fd_sc_hs__clkbuf_2_3/a_43_192# sky130_fd_sc_hs__clkbuf_2
Xsky130_fd_sc_hs__einvp_4_17 DVSS DVDD DVDD DVSS pi5_l[2] sky130_fd_sc_hs__inv_8_9/A
+ sky130_fd_sc_hs__inv_4_19/Y sky130_fd_sc_hs__einvp_4_17/a_27_74# sky130_fd_sc_hs__einvp_4_17/a_27_368#
+ sky130_fd_sc_hs__einvp_4_17/a_473_323# sky130_fd_sc_hs__einvp_4
Xsky130_fd_sc_hs__dlygate4sd3_1_14 DVSS DVDD DVSS DVDD sky130_fd_sc_hs__dlygate4sd3_1_9/X
+ sky130_fd_sc_hs__clkbuf_1_1/A sky130_fd_sc_hs__dlygate4sd3_1_14/a_405_138# sky130_fd_sc_hs__dlygate4sd3_1_14/a_28_74#
+ sky130_fd_sc_hs__dlygate4sd3_1_14/a_289_74# sky130_fd_sc_hs__dlygate4sd3_1
Xsky130_fd_sc_hs__dlygate4sd3_1_25 DVSS DVDD DVSS DVDD sky130_fd_sc_hs__dlygate4sd3_1_3/X
+ sky130_fd_sc_hs__dlygate4sd3_1_25/X sky130_fd_sc_hs__dlygate4sd3_1_25/a_405_138#
+ sky130_fd_sc_hs__dlygate4sd3_1_25/a_28_74# sky130_fd_sc_hs__dlygate4sd3_1_25/a_289_74#
+ sky130_fd_sc_hs__dlygate4sd3_1
Xsky130_fd_sc_hs__dlygate4sd3_1_36 DVSS DVDD DVSS DVDD sky130_fd_sc_hs__dlygate4sd3_1_37/A
+ sky130_fd_sc_hs__dlygate4sd3_1_56/A sky130_fd_sc_hs__dlygate4sd3_1_37/a_405_138#
+ sky130_fd_sc_hs__dlygate4sd3_1_37/a_28_74# sky130_fd_sc_hs__dlygate4sd3_1_37/a_289_74#
+ sky130_fd_sc_hs__dlygate4sd3_1
Xsky130_fd_sc_hs__dlygate4sd3_1_47 DVSS DVDD DVSS DVDD sky130_fd_sc_hs__dlygate4sd3_1_49/X
+ sky130_fd_sc_hs__nand3_4_3/C sky130_fd_sc_hs__dlygate4sd3_1_47/a_405_138# sky130_fd_sc_hs__dlygate4sd3_1_47/a_28_74#
+ sky130_fd_sc_hs__dlygate4sd3_1_47/a_289_74# sky130_fd_sc_hs__dlygate4sd3_1
Xsky130_fd_sc_hs__dlygate4sd3_1_58 DVSS DVDD DVSS DVDD sky130_fd_sc_hs__dlygate4sd3_1_65/X
+ sky130_fd_sc_hs__dlygate4sd3_1_59/X sky130_fd_sc_hs__dlygate4sd3_1_59/a_405_138#
+ sky130_fd_sc_hs__dlygate4sd3_1_59/a_28_74# sky130_fd_sc_hs__dlygate4sd3_1_59/a_289_74#
+ sky130_fd_sc_hs__dlygate4sd3_1
Xsky130_fd_sc_hs__dlygate4sd3_1_69 DVSS DVDD DVSS DVDD sky130_fd_sc_hs__dlygate4sd3_1_71/X
+ sky130_fd_sc_hs__dlygate4sd2_1_1/A sky130_fd_sc_hs__dlygate4sd3_1_69/a_405_138#
+ sky130_fd_sc_hs__dlygate4sd3_1_69/a_28_74# sky130_fd_sc_hs__dlygate4sd3_1_69/a_289_74#
+ sky130_fd_sc_hs__dlygate4sd3_1
Xsky130_fd_sc_hs__nand2_4_8 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_4_9/Y delay_con_msb[2]
+ osc_144 sky130_fd_sc_hs__nand2_4_9/a_27_74# sky130_fd_sc_hs__nand2_4
Xsky130_fd_sc_hs__nand2_2_107 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_2_109/Y sky130_fd_sc_hs__a21oi_1_49/Y
+ osc_036 sky130_fd_sc_hs__nand2_2_109/a_27_74# sky130_fd_sc_hs__nand2_2
Xsky130_fd_sc_hs__einvp_8_9 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_8_5/A pi4_r[3]
+ sky130_fd_sc_hs__inv_4_13/Y sky130_fd_sc_hs__einvp_8_9/a_802_323# sky130_fd_sc_hs__einvp_8_9/a_27_74#
+ sky130_fd_sc_hs__einvp_8_9/a_27_368# sky130_fd_sc_hs__einvp_8
Xsky130_fd_sc_hs__inv_16_14 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__and4_2_5/A sky130_fd_sc_hs__inv_16_7/Y
+ sky130_fd_sc_hs__inv_16
Xsky130_fd_sc_hs__inv_16_25 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_16_9/A sky130_fd_sc_hs__inv_4_25/Y
+ sky130_fd_sc_hs__inv_16
Xsky130_fd_sc_hs__nand2_2_5 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__nand2_2_5/Y sky130_fd_sc_hs__nand2_2_5/B
+ osc_000 sky130_fd_sc_hs__nand2_2_5/a_27_74# sky130_fd_sc_hs__nand2_2
Xsky130_fd_sc_hs__einvp_1_18 DVSS DVDD DVDD DVSS pi5_r[0] sky130_fd_sc_hs__inv_8_9/A
+ sky130_fd_sc_hs__inv_4_21/Y sky130_fd_sc_hs__einvp_1_19/a_44_549# sky130_fd_sc_hs__einvp_1_19/a_318_74#
+ sky130_fd_sc_hs__einvp_1_19/a_310_392# sky130_fd_sc_hs__einvp_1
.ends

.subckt sky130_fd_sc_hs__clkinv_8 VNB VPB VPWR VGND A Y
X0 VPWR A Y VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X1 VGND A Y VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 VPWR A Y VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X3 Y A VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X4 VGND A Y VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 Y A VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X6 Y A VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7 VPWR A Y VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X8 VPWR A Y VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X9 Y A VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X10 Y A VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11 VGND A Y VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12 VGND A Y VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13 VPWR A Y VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X14 Y A VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15 Y A VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X16 VPWR A Y VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X17 Y A VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X18 Y A VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X19 Y A VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
.ends

.subckt sky130_fd_sc_hs__einvn_4 VNB VPB VPWR VGND TE_B A Z a_114_74# a_241_368# a_281_74#
X0 Z A a_241_368# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X1 a_281_74# A Z VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X2 a_114_74# TE_B VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X3 a_241_368# TE_B VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X4 VGND a_114_74# a_281_74# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X5 a_114_74# TE_B VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X6 Z A a_281_74# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X7 VPWR TE_B a_241_368# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X8 a_241_368# TE_B VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X9 Z A a_281_74# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X10 VGND a_114_74# a_281_74# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X11 a_281_74# A Z VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X12 VPWR TE_B a_241_368# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X13 a_281_74# a_114_74# VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X14 a_241_368# A Z VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X15 a_281_74# a_114_74# VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X16 Z A a_241_368# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X17 a_241_368# A Z VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
.ends

.subckt sky130_fd_sc_hs__buf_8 VNB VPB VPWR VGND X A a_27_74#
X0 VPWR a_27_74# X VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X1 X a_27_74# VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X2 VGND A a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X3 VPWR A a_27_74# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X4 X a_27_74# VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X5 VGND a_27_74# X VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X6 VGND A a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X7 a_27_74# A VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X8 VPWR a_27_74# X VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X9 VGND a_27_74# X VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X10 VPWR a_27_74# X VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X11 X a_27_74# VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X12 X a_27_74# VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X13 VPWR a_27_74# X VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X14 X a_27_74# VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X15 VPWR A a_27_74# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X16 X a_27_74# VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X17 a_27_74# A VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X18 X a_27_74# VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X19 X a_27_74# VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X20 VGND a_27_74# X VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X21 VGND a_27_74# X VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
.ends

.subckt sky130_fd_sc_hs__einvn_2 VNB VPB VPWR VGND TE_B A Z a_227_368# a_231_74# a_115_464#
X0 a_231_74# a_115_464# VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X1 VPWR TE_B a_227_368# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X2 a_115_464# TE_B VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X3 a_115_464# TE_B VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4 VGND a_115_464# a_231_74# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X5 Z A a_231_74# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X6 a_231_74# A Z VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X7 a_227_368# A Z VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X8 Z A a_227_368# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X9 a_227_368# TE_B VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
.ends

.subckt sky130_fd_sc_hs__or4_2 VNB VPB VPWR VGND X D A B C a_174_392# a_258_392# a_342_392#
+ a_85_392#
X0 a_174_392# D a_85_392# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 VGND A a_85_392# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X2 X a_85_392# VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X3 VPWR A a_342_392# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 a_85_392# B VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X5 a_85_392# D VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X6 VGND C a_85_392# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X7 a_342_392# B a_258_392# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 VGND a_85_392# X VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X9 VPWR a_85_392# X VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X10 a_258_392# C a_174_392# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 X a_85_392# VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
.ends

.subckt hr_16t4_mux_top clk din[15] din[14] din[13] din[12] din[11] din[10] din[9]
+ din[8] din[7] din[6] din[5] din[4] din[3] din[2] din[1] din[0] rst clk_prbs dout[3]
+ dout[2] dout[1] dout[0] DVSS DVDD sky130_fd_sc_hs__dfxtp_4_31/D sky130_fd_sc_hs__dfxtp_4_15/a_735_102#
+ sky130_fd_sc_hs__dfxtp_4_23/Q sky130_fd_sc_hs__clkbuf_4_1/X sky130_fd_sc_hs__inv_4_11/A
+ sky130_fd_sc_hs__clkbuf_2_25/a_43_192# sky130_fd_sc_hs__inv_4_19/A sky130_fd_sc_hs__dfrtp_4_3/a_890_138#
+ sky130_fd_sc_hs__buf_2_11/a_21_260# sky130_fd_sc_hs__dfxtp_4_1/a_1141_508# sky130_fd_sc_hs__dfxtp_4_5/Q
+ sky130_fd_sc_hs__dfxtp_4_29/a_544_485# sky130_fd_sc_hs__dfxtp_4_39/a_696_458# sky130_fd_sc_hs__dfxtp_4_46/a_735_102#
+ sky130_fd_sc_hs__dfxtp_4_47/a_1034_424# sky130_fd_sc_hs__dfxtp_4_24/D sky130_fd_sc_hs__a22o_1_9/A2
+ sky130_fd_sc_hs__a22o_1_9/B1 sky130_fd_sc_hs__dfxtp_4_8/a_27_74# sky130_fd_sc_hs__a22o_1_5/X
+ sky130_fd_sc_hs__dfxtp_4_19/a_651_503# sky130_fd_sc_hs__a22o_1_7/X sky130_fd_sc_hs__dfxtp_4_33/a_735_102#
+ sky130_fd_sc_hs__dfxtp_4_31/a_27_74# sky130_fd_sc_hs__dfxtp_4_46/a_1034_424# sky130_fd_sc_hs__clkinv_4_1/Y
+ sky130_fd_sc_hs__dfxtp_4_25/a_1141_508# sky130_fd_sc_hs__dfxtp_4_46/Q sky130_fd_sc_hs__dfxtp_4_46/D
+ sky130_fd_sc_hs__dfxtp_4_35/a_1226_296# sky130_fd_sc_hs__dfxtp_4_5/a_696_458# sky130_fd_sc_hs__dfxtp_4_41/Q
+ sky130_fd_sc_hs__dfxtp_4_45/a_1034_424# sky130_fd_sc_hs__dfxtp_4_24/a_1141_508#
+ sky130_fd_sc_hs__clkbuf_2_11/a_43_192# sky130_fd_sc_hs__dfxtp_4_33/a_1226_296# sky130_fd_sc_hs__a22o_1_15/a_230_79#
+ sky130_fd_sc_hs__dfxtp_4_47/a_206_368# sky130_fd_sc_hs__dfxtp_4_39/a_544_485# sky130_fd_sc_hs__dfxtp_4_13/a_735_102#
+ sky130_fd_sc_hs__dfxtp_4_33/Q sky130_fd_sc_hs__dfxtp_4_23/a_1141_508# sky130_fd_sc_hs__clkbuf_2_15/a_43_192#
+ sky130_fd_sc_hs__dfxtp_4_45/D sky130_fd_sc_hs__dfxtp_4_29/Q sky130_fd_sc_hs__dfxtp_4_35/a_206_368#
+ sky130_fd_sc_hs__dfxtp_4_47/a_437_503# sky130_fd_sc_hs__dfxtp_4_27/a_651_503# sky130_fd_sc_hs__inv_4_1/Y
+ sky130_fd_sc_hs__a22o_1_17/X sky130_fd_sc_hs__dfxtp_4_45/a_735_102# sky130_fd_sc_hs__dfxtp_4_37/a_696_458#
+ sky130_fd_sc_hs__dfxtp_4_41/a_1034_424# sky130_fd_sc_hs__a22o_1_15/a_222_392# sky130_fd_sc_hs__dfxtp_4_39/a_1141_508#
+ sky130_fd_sc_hs__a22o_1_15/a_52_123# sky130_fd_sc_hs__dfxtp_4_3/a_651_503# sky130_fd_sc_hs__dfxtp_4_15/D
+ sky130_fd_sc_hs__dfxtp_4_5/a_544_485# sky130_fd_sc_hs__clkbuf_2_19/a_43_192# sky130_fd_sc_hs__dfxtp_4_19/a_1178_124#
+ sky130_fd_sc_hs__dfxtp_4_35/a_437_503# sky130_fd_sc_hs__dfxtp_4_18/a_651_503# sky130_fd_sc_hs__inv_4_5/Y
+ sky130_fd_sc_hs__dfxtp_4_37/a_1141_508# sky130_fd_sc_hs__dfxtp_4_31/a_1226_296#
+ sky130_fd_sc_hs__dfxtp_4_47/D sky130_fd_sc_hs__dfxtp_4_1/a_206_368# sky130_fd_sc_hs__dfxtp_4_33/a_27_74#
+ sky130_fd_sc_hs__dfxtp_4_18/a_1178_124# sky130_fd_sc_hs__dfxtp_4_15/a_206_368# sky130_fd_sc_hs__a22o_1_23/a_132_392#
+ sky130_fd_sc_hs__dfxtp_4_5/D sky130_fd_sc_hs__dfxtp_4_19/a_696_458# sky130_fd_sc_hs__dfrtp_4_3/a_313_74#
+ sky130_fd_sc_hs__dfxtp_4_25/a_735_102# sky130_fd_sc_hs__buf_2_5/X sky130_fd_sc_hs__a22o_1_5/B2
+ sky130_fd_sc_hs__dfxtp_4_35/Q sky130_fd_sc_hs__dfrtp_4_3/a_494_366# sky130_fd_sc_hs__dfxtp_4_1/a_437_503#
+ sky130_fd_sc_hs__clkbuf_4_3/a_83_270# sky130_fd_sc_hs__clkbuf_2_9/a_43_192# sky130_fd_sc_hs__a22o_1_19/X
+ sky130_fd_sc_hs__dfxtp_4_9/a_735_102# sky130_fd_sc_hs__dfxtp_4_15/a_437_503# sky130_fd_sc_hs__dfxtp_4_46/a_206_368#
+ sky130_fd_sc_hs__dfxtp_4_37/a_544_485# sky130_fd_sc_hs__dfrtp_4_1/a_1647_81# sky130_fd_sc_hs__dfxtp_4_8/Q
+ sky130_fd_sc_hs__dfrtp_4_1/a_890_138# sky130_fd_sc_hs__dfxtp_4_15/a_1178_124# sky130_fd_sc_hs__a22o_1_21/a_230_79#
+ sky130_fd_sc_hs__dfxtp_4_33/a_206_368# sky130_fd_sc_hs__a22o_1_1/a_222_392# sky130_fd_sc_hs__dfxtp_4_46/a_437_503#
+ sky130_fd_sc_hs__clkinv_2_1/Y sky130_fd_sc_hs__dfxtp_4_45/a_27_74# sky130_fd_sc_hs__a22o_1_14/a_222_392#
+ sky130_fd_sc_hs__dfxtp_4_35/a_1141_508# sky130_fd_sc_hs__dfxtp_4_9/a_1178_124# sky130_fd_sc_hs__dfxtp_4_13/a_1178_124#
+ sky130_fd_sc_hs__dfxtp_4_33/a_437_503# sky130_fd_sc_hs__dfxtp_4_19/a_544_485# sky130_fd_sc_hs__dfxtp_4_27/D
+ sky130_fd_sc_hs__dfxtp_4_27/a_696_458# sky130_fd_sc_hs__dfxtp_4_33/a_1141_508# sky130_fd_sc_hs__dfxtp_4_8/a_1178_124#
+ sky130_fd_sc_hs__dfxtp_4_5/a_27_74# sky130_fd_sc_hs__buf_2_15/X sky130_fd_sc_hs__inv_4_11/Y
+ sky130_fd_sc_hs__dfxtp_4_18/Q sky130_fd_sc_hs__dfxtp_4_3/a_696_458# sky130_fd_sc_hs__dfxtp_4_13/a_206_368#
+ sky130_fd_sc_hs__a22o_1_21/a_52_123# sky130_fd_sc_hs__dfxtp_4_47/a_651_503# sky130_fd_sc_hs__dfxtp_4_3/D
+ sky130_fd_sc_hs__dfxtp_4_18/a_696_458# sky130_fd_sc_hs__dfxtp_4_24/a_735_102# sky130_fd_sc_hs__clkbuf_2_23/a_43_192#
+ sky130_fd_sc_hs__dfxtp_4_7/a_1178_124# sky130_fd_sc_hs__dfxtp_4_47/a_1226_296# sky130_fd_sc_hs__a22o_1_9/a_132_392#
+ sky130_fd_sc_hs__dfxtp_4_8/a_735_102# sky130_fd_sc_hs__dfxtp_4_45/a_206_368# sky130_fd_sc_hs__dfxtp_4_13/a_437_503#
+ sky130_fd_sc_hs__dfxtp_4_35/a_651_503# sky130_fd_sc_hs__dfrtp_4_3/a_2010_409# sky130_fd_sc_hs__dfxtp_4_46/a_1226_296#
+ sky130_fd_sc_hs__a22o_1_1/a_230_79# sky130_fd_sc_hs__dfxtp_4_45/Q sky130_fd_sc_hs__dfxtp_4_23/a_27_74#
+ sky130_fd_sc_hs__a22o_1_11/a_230_79# sky130_fd_sc_hs__dfxtp_4_29/a_1178_124# sky130_fd_sc_hs__dfxtp_4_45/a_437_503#
+ sky130_fd_sc_hs__dfxtp_4_27/a_544_485# sky130_fd_sc_hs__dfxtp_4_37/Q sky130_fd_sc_hs__dfxtp_4_41/a_735_102#
+ sky130_fd_sc_hs__dfxtp_4_31/a_1141_508# sky130_fd_sc_hs__inv_4_9/Y sky130_fd_sc_hs__dfxtp_4_45/a_1226_296#
+ sky130_fd_sc_hs__dfrtp_4_1/a_37_78# sky130_fd_sc_hs__dfxtp_4_1/a_651_503# sky130_fd_sc_hs__dfxtp_4_3/a_544_485#
+ sky130_fd_sc_hs__a22o_1_1/X sky130_fd_sc_hs__dfxtp_4_25/a_206_368# sky130_fd_sc_hs__a22o_1_5/a_230_79#
+ sky130_fd_sc_hs__dfxtp_4_15/a_651_503# sky130_fd_sc_hs__dfxtp_4_18/a_544_485# sky130_fd_sc_hs__a22o_1_14/a_230_79#
+ sky130_fd_sc_hs__dfrtp_4_1/a_2010_409# sky130_fd_sc_hs__dfxtp_4_31/a_735_102# sky130_fd_sc_hs__a22o_1_23/X
+ sky130_fd_sc_hs__dfxtp_4_5/a_1178_124# sky130_fd_sc_hs__buf_2_11/X sky130_fd_sc_hs__inv_4_19/Y
+ sky130_fd_sc_hs__dfxtp_4_9/a_206_368# sky130_fd_sc_hs__a22o_1_1/a_52_123# sky130_fd_sc_hs__dfxtp_4_15/a_27_74#
+ sky130_fd_sc_hs__a22o_1_21/a_132_392# sky130_fd_sc_hs__dfxtp_4_7/a_27_74# sky130_fd_sc_hs__dfxtp_4_1/D
+ sky130_fd_sc_hs__a22o_1_11/a_52_123# sky130_fd_sc_hs__dfxtp_4_25/a_437_503# sky130_fd_sc_hs__dfxtp_4_46/a_651_503#
+ sky130_fd_sc_hs__dfxtp_4_23/a_735_102# sky130_fd_sc_hs__a22o_1_9/a_230_79# sky130_fd_sc_hs__clkbuf_2_13/a_43_192#
+ sky130_fd_sc_hs__dfxtp_4_31/Q sky130_fd_sc_hs__a22o_1_19/a_230_79# sky130_fd_sc_hs__dfxtp_4_41/a_1226_296#
+ sky130_fd_sc_hs__dfrtp_4_1/a_494_366# sky130_fd_sc_hs__dfxtp_4_19/a_1034_424# sky130_fd_sc_hs__a22o_1_21/X
+ sky130_fd_sc_hs__dfxtp_4_9/a_437_503# sky130_fd_sc_hs__dfxtp_4_7/a_735_102# sky130_fd_sc_hs__dfxtp_4_27/a_1178_124#
+ sky130_fd_sc_hs__a22o_1_11/a_132_392# sky130_fd_sc_hs__clkbuf_2_1/a_43_192# sky130_fd_sc_hs__dfxtp_4_33/a_651_503#
+ sky130_fd_sc_hs__a22o_1_5/a_52_123# sky130_fd_sc_hs__dfxtp_4_47/a_696_458# sky130_fd_sc_hs__a22o_1_14/a_52_123#
+ sky130_fd_sc_hs__dfxtp_4_3/a_1178_124# sky130_fd_sc_hs__a22o_1_23/a_222_392# sky130_fd_sc_hs__dfxtp_4_39/D
+ sky130_fd_sc_hs__dfxtp_4_18/a_1034_424# sky130_fd_sc_hs__clkbuf_2_17/a_43_192# sky130_fd_sc_hs__dfrtp_4_1/Q
+ sky130_fd_sc_hs__dfxtp_4_35/a_696_458# sky130_fd_sc_hs__clkbuf_2_5/a_43_192# sky130_fd_sc_hs__inv_4_7/Y
+ sky130_fd_sc_hs__a22o_1_9/a_52_123# sky130_fd_sc_hs__a22o_1_19/a_52_123# sky130_fd_sc_hs__dfrtp_4_3/a_699_463#
+ sky130_fd_sc_hs__dfxtp_4_24/a_206_368# sky130_fd_sc_hs__dfxtp_4_13/a_651_503# sky130_fd_sc_hs__inv_4_21/Y
+ sky130_fd_sc_hs__dfxtp_4_47/a_1141_508# sky130_fd_sc_hs__dfxtp_4_1/a_1178_124# sky130_fd_sc_hs__inv_4_13/Y
+ sky130_fd_sc_hs__dfxtp_4_15/a_1034_424# sky130_fd_sc_hs__dfxtp_4_8/a_206_368# sky130_fd_sc_hs__dfxtp_4_1/a_696_458#
+ sky130_fd_sc_hs__dfxtp_4_19/Q sky130_fd_sc_hs__dfxtp_4_9/a_1034_424# sky130_fd_sc_hs__dfxtp_4_24/a_437_503#
+ sky130_fd_sc_hs__dfxtp_4_1/a_27_74# sky130_fd_sc_hs__dfxtp_4_45/a_651_503# sky130_fd_sc_hs__dfxtp_4_47/a_544_485#
+ sky130_fd_sc_hs__dfxtp_4_15/a_696_458# sky130_fd_sc_hs__dfxtp_4_46/a_1141_508# sky130_fd_sc_hs__buf_2_14/X
+ sky130_fd_sc_hs__dfxtp_4_9/D sky130_fd_sc_hs__dfxtp_4_13/a_1034_424# sky130_fd_sc_hs__dfxtp_4_19/a_27_74#
+ sky130_fd_sc_hs__a22o_1_7/a_132_392# sky130_fd_sc_hs__dfxtp_4_8/a_437_503# sky130_fd_sc_hs__dfxtp_4_27/Q
+ sky130_fd_sc_hs__buf_2_9/X sky130_fd_sc_hs__dfxtp_4_25/a_1178_124# sky130_fd_sc_hs__dfxtp_4_8/a_1034_424#
+ sky130_fd_sc_hs__dfxtp_4_41/a_206_368# sky130_fd_sc_hs__dfxtp_4_35/a_544_485# sky130_fd_sc_hs__dfxtp_4_46/a_696_458#
+ sky130_fd_sc_hs__dfxtp_4_45/a_1141_508# sky130_fd_sc_hs__dfxtp_4_24/a_1178_124#
+ sky130_fd_sc_hs__a22o_1_9/a_222_392# sky130_fd_sc_hs__dfxtp_4_7/a_1034_424# sky130_fd_sc_hs__dfxtp_4_31/a_206_368#
+ sky130_fd_sc_hs__dfxtp_4_25/a_651_503# sky130_fd_sc_hs__dfxtp_4_41/a_437_503# sky130_fd_sc_hs__dfxtp_4_33/a_696_458#
+ sky130_fd_sc_hs__buf_2_3/a_21_260# sky130_fd_sc_hs__dfxtp_4_25/D sky130_fd_sc_hs__a22o_1_7/A2
+ sky130_fd_sc_hs__dfxtp_4_9/a_651_503# sky130_fd_sc_hs__clkbuf_1_1/a_27_74# sky130_fd_sc_hs__dfxtp_4_1/a_544_485#
+ sky130_fd_sc_hs__dfxtp_4_23/a_1178_124# sky130_fd_sc_hs__dfxtp_4_27/a_27_74# sky130_fd_sc_hs__dfxtp_4_23/a_206_368#
+ sky130_fd_sc_hs__dfxtp_4_31/a_437_503# sky130_fd_sc_hs__dfxtp_4_15/a_544_485# sky130_fd_sc_hs__dfxtp_4_41/a_1141_508#
+ sky130_fd_sc_hs__dfrtp_4_3/a_124_78# sky130_fd_sc_hs__dfxtp_4_47/Q sky130_fd_sc_hs__dfxtp_4_29/a_1034_424#
+ sky130_fd_sc_hs__buf_2_7/a_21_260# sky130_fd_sc_hs__dfxtp_4_7/a_206_368# sky130_fd_sc_hs__dfxtp_4_39/a_1178_124#
+ sky130_fd_sc_hs__dfxtp_4_23/a_437_503# sky130_fd_sc_hs__dfxtp_4_7/Q sky130_fd_sc_hs__dfxtp_4_46/a_544_485#
+ sky130_fd_sc_hs__dfxtp_4_13/a_696_458# sky130_fd_sc_hs__dfxtp_4_29/a_735_102# sky130_fd_sc_hs__clkbuf_2_27/a_43_192#
+ sky130_fd_sc_hs__a22o_1_3/X sky130_fd_sc_hs__buf_2_15/a_21_260# sky130_fd_sc_hs__dfxtp_4_7/a_437_503#
+ sky130_fd_sc_hs__dfxtp_4_37/a_1178_124# sky130_fd_sc_hs__dfxtp_4_5/a_1034_424# sky130_fd_sc_hs__dfxtp_4_33/a_544_485#
+ sky130_fd_sc_hs__dfxtp_4_45/a_696_458# sky130_fd_sc_hs__dfrtp_4_3/a_1827_81# sky130_fd_sc_hs__a22o_1_21/a_222_392#
+ sky130_fd_sc_hs__a22o_1_3/a_230_79# sky130_fd_sc_hs__inv_4_17/Y sky130_fd_sc_hs__dfxtp_4_24/a_651_503#
+ sky130_fd_sc_hs__inv_4_3/Y sky130_fd_sc_hs__a22o_1_11/a_222_392# sky130_fd_sc_hs__dfxtp_4_27/a_1034_424#
+ sky130_fd_sc_hs__dfxtp_4_19/a_1226_296# sky130_fd_sc_hs__dfxtp_4_8/a_651_503# sky130_fd_sc_hs__dfrtp_4_1/a_699_463#
+ sky130_fd_sc_hs__buf_2_7/X sky130_fd_sc_hs__dfxtp_4_3/a_1034_424# sky130_fd_sc_hs__a22o_1_17/a_230_79#
+ sky130_fd_sc_hs__dfxtp_4_13/a_544_485# sky130_fd_sc_hs__dfxtp_4_25/a_696_458# sky130_fd_sc_hs__dfxtp_4_39/a_735_102#
+ sky130_fd_sc_hs__dfxtp_4_29/a_27_74# sky130_fd_sc_hs__dfxtp_4_18/a_1226_296# sky130_fd_sc_hs__dfxtp_4_9/a_696_458#
+ sky130_fd_sc_hs__a22o_1_3/a_52_123# sky130_fd_sc_hs__dfxtp_4_35/a_1178_124# sky130_fd_sc_hs__dfxtp_4_47/a_27_74#
+ sky130_fd_sc_hs__dfxtp_4_3/Q sky130_fd_sc_hs__dfxtp_4_41/a_651_503# sky130_fd_sc_hs__dfxtp_4_45/a_544_485#
+ sky130_fd_sc_hs__dfxtp_4_35/D sky130_fd_sc_hs__dfrtp_4_3/a_789_463# sky130_fd_sc_hs__a22o_1_5/a_132_392#
+ sky130_fd_sc_hs__dfxtp_4_33/a_1178_124# sky130_fd_sc_hs__dfxtp_4_5/a_735_102# sky130_fd_sc_hs__dfxtp_4_1/a_1034_424#
+ sky130_fd_sc_hs__a22o_1_19/a_132_392# sky130_fd_sc_hs__dfxtp_4_13/a_27_74# sky130_fd_sc_hs__dfxtp_4_31/a_651_503#
+ sky130_fd_sc_hs__a22o_1_17/a_52_123# sky130_fd_sc_hs__dfrtp_4_1/a_313_74# sky130_fd_sc_hs__dfxtp_4_23/D
+ sky130_fd_sc_hs__dfxtp_4_15/a_1226_296# sky130_fd_sc_hs__clkbuf_2_31/a_43_192# sky130_fd_sc_hs__inv_4_15/Y
+ sky130_fd_sc_hs__dfxtp_4_39/a_27_74# sky130_fd_sc_hs__a22o_1_7/a_222_392# sky130_fd_sc_hs__clkbuf_4_1/a_83_270#
+ sky130_fd_sc_hs__dfxtp_4_23/a_651_503# sky130_fd_sc_hs__dfxtp_4_25/a_544_485# sky130_fd_sc_hs__clkbuf_2_7/a_43_192#
+ sky130_fd_sc_hs__dfxtp_4_9/a_1226_296# sky130_fd_sc_hs__dfxtp_4_8/D sky130_fd_sc_hs__dfxtp_4_25/a_1034_424#
+ sky130_fd_sc_hs__dfrtp_4_3/a_834_355# sky130_fd_sc_hs__dfxtp_4_13/a_1226_296# sky130_fd_sc_hs__dfxtp_4_7/a_651_503#
+ sky130_fd_sc_hs__dfrtp_4_3/a_1627_493# sky130_fd_sc_hs__dfxtp_4_9/a_544_485# sky130_fd_sc_hs__dfxtp_4_29/a_206_368#
+ sky130_fd_sc_hs__dfrtp_4_3/a_812_138# sky130_fd_sc_hs__dfxtp_4_24/a_696_458# sky130_fd_sc_hs__dfxtp_4_8/a_1226_296#
+ sky130_fd_sc_hs__dfxtp_4_37/a_735_102# sky130_fd_sc_hs__dfxtp_4_24/a_1034_424# sky130_fd_sc_hs__dfxtp_4_25/a_27_74#
+ sky130_fd_sc_hs__dfxtp_4_31/a_1178_124# sky130_fd_sc_hs__dfxtp_4_8/a_696_458# sky130_fd_sc_hs__dfxtp_4_1/Q
+ sky130_fd_sc_hs__dfxtp_4_29/a_437_503# sky130_fd_sc_hs__dfxtp_4_7/a_1226_296# sky130_fd_sc_hs__dfrtp_4_3/a_37_78#
+ sky130_fd_sc_hs__dfxtp_4_23/a_1034_424# sky130_fd_sc_hs__a22o_1_23/a_230_79# sky130_fd_sc_hs__a22o_1_3/a_132_392#
+ sky130_fd_sc_hs__dfrtp_4_1/a_1627_493# sky130_fd_sc_hs__a22o_1_17/a_132_392# sky130_fd_sc_hs__dfxtp_4_19/a_735_102#
+ sky130_fd_sc_hs__dfxtp_4_41/a_696_458# sky130_fd_sc_hs__dfrtp_4_1/a_1827_81# sky130_fd_sc_hs__dfxtp_4_39/a_1034_424#
+ sky130_fd_sc_hs__dfxtp_4_19/a_1141_508# sky130_fd_sc_hs__dfxtp_4_9/a_27_74# sky130_fd_sc_hs__dfxtp_4_29/a_1226_296#
+ sky130_fd_sc_hs__dfxtp_4_18/a_27_74# sky130_fd_sc_hs__dfxtp_4_39/a_206_368# sky130_fd_sc_hs__dfxtp_4_24/a_544_485#
+ sky130_fd_sc_hs__dfxtp_4_31/a_696_458# sky130_fd_sc_hs__dfxtp_4_37/a_1034_424# sky130_fd_sc_hs__dfxtp_4_18/a_1141_508#
+ sky130_fd_sc_hs__dfxtp_4_9/Q sky130_fd_sc_hs__a22o_1_23/a_52_123# sky130_fd_sc_hs__dfxtp_4_8/a_544_485#
+ sky130_fd_sc_hs__buf_2_3/X sky130_fd_sc_hs__buf_2_14/a_21_260# sky130_fd_sc_hs__dfxtp_4_5/a_1226_296#
+ sky130_fd_sc_hs__dfxtp_4_39/a_437_503# sky130_fd_sc_hs__dfxtp_4_23/a_696_458# sky130_fd_sc_hs__buf_2_9/a_21_260#
+ sky130_fd_sc_hs__dfxtp_4_5/a_206_368# sky130_fd_sc_hs__dfxtp_4_7/a_696_458# sky130_fd_sc_hs__dfxtp_4_39/Q
+ sky130_fd_sc_hs__dfrtp_4_3/a_1678_395# sky130_fd_sc_hs__dfxtp_4_41/a_544_485# sky130_fd_sc_hs__clkbuf_2_29/a_43_192#
+ sky130_fd_sc_hs__dfxtp_4_27/a_735_102# sky130_fd_sc_hs__dfrtp_4_1/a_789_463# sky130_fd_sc_hs__dfxtp_4_15/a_1141_508#
+ sky130_fd_sc_hs__buf_2_1/X sky130_fd_sc_hs__dfxtp_4_41/a_27_74# sky130_fd_sc_hs__dfxtp_4_5/a_437_503#
+ sky130_fd_sc_hs__dfxtp_4_27/a_1226_296# sky130_fd_sc_hs__dfxtp_4_3/a_735_102# sky130_fd_sc_hs__dfxtp_4_47/a_1178_124#
+ sky130_fd_sc_hs__dfxtp_4_9/a_1141_508# sky130_fd_sc_hs__dfxtp_4_3/a_1226_296# sky130_fd_sc_hs__dfxtp_4_18/a_735_102#
+ sky130_fd_sc_hs__dfxtp_4_31/a_544_485# sky130_fd_sc_hs__dfxtp_4_35/a_1034_424# sky130_fd_sc_hs__dfxtp_4_13/a_1141_508#
+ sky130_fd_sc_hs__a22o_1_7/a_230_79# sky130_fd_sc_hs__dfxtp_4_3/a_27_74# sky130_fd_sc_hs__dfxtp_4_46/a_1178_124#
+ sky130_fd_sc_hs__dfxtp_4_8/a_1141_508# sky130_fd_sc_hs__dfrtp_4_1/a_1678_395# sky130_fd_sc_hs__a22o_1_5/a_222_392#
+ sky130_fd_sc_hs__dfxtp_4_37/a_206_368# sky130_fd_sc_hs__dfxtp_4_23/a_544_485# sky130_fd_sc_hs__dfxtp_4_29/a_651_503#
+ sky130_fd_sc_hs__a22o_1_7/B2 sky130_fd_sc_hs__a22o_1_19/a_222_392# sky130_fd_sc_hs__dfxtp_4_33/a_1034_424#
+ sky130_fd_sc_hs__dfrtp_4_1/a_834_355# sky130_fd_sc_hs__dfxtp_4_35/a_27_74# sky130_fd_sc_hs__dfxtp_4_7/a_544_485#
+ sky130_fd_sc_hs__dfxtp_4_45/a_1178_124# sky130_fd_sc_hs__dfxtp_4_7/a_1141_508# sky130_fd_sc_hs__dfrtp_4_1/a_812_138#
+ sky130_fd_sc_hs__dfxtp_4_1/a_1226_296# sky130_fd_sc_hs__dfxtp_4_37/a_437_503# sky130_fd_sc_hs__clkbuf_2_3/a_43_192#
+ sky130_fd_sc_hs__a22o_1_7/a_52_123# sky130_fd_sc_hs__dfrtp_4_3/a_1350_392# sky130_fd_sc_hs__dfxtp_4_19/a_206_368#
+ sky130_fd_sc_hs__dfxtp_4_29/a_1141_508# sky130_fd_sc_hs__dfxtp_4_25/a_1226_296#
+ sky130_fd_sc_hs__dfxtp_4_41/a_1178_124# sky130_fd_sc_hs__a22o_1_15/a_132_392# sky130_fd_sc_hs__dfxtp_4_19/a_437_503#
+ sky130_fd_sc_hs__dfxtp_4_46/a_27_74# sky130_fd_sc_hs__dfxtp_4_39/a_651_503# sky130_fd_sc_hs__dfxtp_4_31/a_1034_424#
+ sky130_fd_sc_hs__dfxtp_4_24/a_1226_296# sky130_fd_sc_hs__dfrtp_4_1/a_1350_392# sky130_fd_sc_hs__dfxtp_4_5/a_1141_508#
+ sky130_fd_sc_hs__a22o_1_3/a_222_392# sky130_fd_sc_hs__clkbuf_16_1/a_114_74# sky130_fd_sc_hs__dfxtp_4_47/a_735_102#
+ sky130_fd_sc_hs__a22o_1_17/a_222_392# sky130_fd_sc_hs__dfxtp_4_23/a_1226_296# sky130_fd_sc_hs__dfxtp_4_5/a_651_503#
+ sky130_fd_sc_hs__dfxtp_4_27/a_206_368# sky130_fd_sc_hs__dfxtp_4_37/a_27_74# sky130_fd_sc_hs__dfxtp_4_29/a_696_458#
+ sky130_fd_sc_hs__dfxtp_4_35/a_735_102# sky130_fd_sc_hs__dfxtp_4_27/a_1141_508# sky130_fd_sc_hs__dfxtp_4_3/a_206_368#
+ sky130_fd_sc_hs__dfxtp_4_39/a_1226_296# sky130_fd_sc_hs__buf_2_1/a_21_260# sky130_fd_sc_hs__dfxtp_4_3/a_1141_508#
+ sky130_fd_sc_hs__dfxtp_4_18/a_206_368# sky130_fd_sc_hs__dfxtp_4_27/a_437_503# sky130_fd_sc_hs__clkbuf_2_21/a_43_192#
+ sky130_fd_sc_hs__a22o_1_1/a_132_392# sky130_fd_sc_hs__dfxtp_4_3/a_437_503# sky130_fd_sc_hs__dfrtp_4_1/a_124_78#
+ sky130_fd_sc_hs__dfxtp_4_37/a_1226_296# sky130_fd_sc_hs__dfxtp_4_24/a_27_74# sky130_fd_sc_hs__dfxtp_4_1/a_735_102#
+ sky130_fd_sc_hs__buf_2_5/a_21_260# sky130_fd_sc_hs__a22o_1_14/a_132_392# sky130_fd_sc_hs__dfxtp_4_37/a_651_503#
+ sky130_fd_sc_hs__dfxtp_4_18/a_437_503# sky130_fd_sc_hs__dfrtp_4_3/a_1647_81#
Xsky130_fd_sc_hs__clkbuf_2_3 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__dfxtp_4_3/D din[15]
+ sky130_fd_sc_hs__clkbuf_2_3/a_43_192# sky130_fd_sc_hs__clkbuf_2
Xsky130_fd_sc_hs__clkbuf_2_25 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__dfxtp_4_35/D din[4]
+ sky130_fd_sc_hs__clkbuf_2_25/a_43_192# sky130_fd_sc_hs__clkbuf_2
Xsky130_fd_sc_hs__a22o_1_14 DVSS DVDD DVDD DVSS dout[2] sky130_fd_sc_hs__dfxtp_4_19/Q
+ sky130_fd_sc_hs__a22o_1_9/B1 sky130_fd_sc_hs__dfxtp_4_18/Q sky130_fd_sc_hs__inv_4_19/A
+ sky130_fd_sc_hs__a22o_1_14/a_222_392# sky130_fd_sc_hs__a22o_1_14/a_230_79# sky130_fd_sc_hs__a22o_1_14/a_52_123#
+ sky130_fd_sc_hs__a22o_1_14/a_132_392# sky130_fd_sc_hs__a22o_1
Xsky130_fd_sc_hs__clkbuf_2_14 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__dfxtp_4_25/D din[8]
+ sky130_fd_sc_hs__clkbuf_2_15/a_43_192# sky130_fd_sc_hs__clkbuf_2
Xsky130_fd_sc_hs__inv_4_8 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_9/Y clk_prbs
+ sky130_fd_sc_hs__inv_4
Xsky130_fd_sc_hs__buf_2_5 DVSS DVDD DVDD DVSS clk_prbs sky130_fd_sc_hs__buf_2_5/X
+ sky130_fd_sc_hs__buf_2_5/a_21_260# sky130_fd_sc_hs__buf_2
Xsky130_fd_sc_hs__dfxtp_4_4 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__dfxtp_4_5/Q sky130_fd_sc_hs__dfxtp_4_5/D
+ sky130_fd_sc_hs__clkbuf_4_1/X sky130_fd_sc_hs__dfxtp_4_5/a_1226_296# sky130_fd_sc_hs__dfxtp_4_5/a_735_102#
+ sky130_fd_sc_hs__dfxtp_4_5/a_1141_508# sky130_fd_sc_hs__dfxtp_4_5/a_206_368# sky130_fd_sc_hs__dfxtp_4_5/a_437_503#
+ sky130_fd_sc_hs__dfxtp_4_5/a_27_74# sky130_fd_sc_hs__dfxtp_4_5/a_651_503# sky130_fd_sc_hs__dfxtp_4_5/a_696_458#
+ sky130_fd_sc_hs__dfxtp_4_5/a_544_485# sky130_fd_sc_hs__dfxtp_4_5/a_1178_124# sky130_fd_sc_hs__dfxtp_4_5/a_1034_424#
+ sky130_fd_sc_hs__dfxtp_4
Xsky130_fd_sc_hs__buf_2_10 DVSS DVDD DVDD DVSS clk_prbs sky130_fd_sc_hs__buf_2_11/X
+ sky130_fd_sc_hs__buf_2_11/a_21_260# sky130_fd_sc_hs__buf_2
Xsky130_fd_sc_hs__inv_4_9 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_9/Y clk_prbs
+ sky130_fd_sc_hs__inv_4
Xsky130_fd_sc_hs__clkbuf_2_4 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__dfxtp_4_5/D din[13]
+ sky130_fd_sc_hs__clkbuf_2_5/a_43_192# sky130_fd_sc_hs__clkbuf_2
Xsky130_fd_sc_hs__clkbuf_2_26 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__dfxtp_4_46/D din[0]
+ sky130_fd_sc_hs__clkbuf_2_27/a_43_192# sky130_fd_sc_hs__clkbuf_2
Xsky130_fd_sc_hs__a22o_1_15 DVSS DVDD DVDD DVSS dout[1] sky130_fd_sc_hs__dfxtp_4_37/Q
+ sky130_fd_sc_hs__a22o_1_9/B1 sky130_fd_sc_hs__dfxtp_4_29/Q sky130_fd_sc_hs__inv_4_19/A
+ sky130_fd_sc_hs__a22o_1_15/a_222_392# sky130_fd_sc_hs__a22o_1_15/a_230_79# sky130_fd_sc_hs__a22o_1_15/a_52_123#
+ sky130_fd_sc_hs__a22o_1_15/a_132_392# sky130_fd_sc_hs__a22o_1
Xsky130_fd_sc_hs__clkbuf_2_15 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__dfxtp_4_25/D din[8]
+ sky130_fd_sc_hs__clkbuf_2_15/a_43_192# sky130_fd_sc_hs__clkbuf_2
Xsky130_fd_sc_hs__buf_2_6 DVSS DVDD DVDD DVSS clk_prbs sky130_fd_sc_hs__buf_2_7/X
+ sky130_fd_sc_hs__buf_2_7/a_21_260# sky130_fd_sc_hs__buf_2
Xsky130_fd_sc_hs__dfxtp_4_5 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__dfxtp_4_5/Q sky130_fd_sc_hs__dfxtp_4_5/D
+ sky130_fd_sc_hs__clkbuf_4_1/X sky130_fd_sc_hs__dfxtp_4_5/a_1226_296# sky130_fd_sc_hs__dfxtp_4_5/a_735_102#
+ sky130_fd_sc_hs__dfxtp_4_5/a_1141_508# sky130_fd_sc_hs__dfxtp_4_5/a_206_368# sky130_fd_sc_hs__dfxtp_4_5/a_437_503#
+ sky130_fd_sc_hs__dfxtp_4_5/a_27_74# sky130_fd_sc_hs__dfxtp_4_5/a_651_503# sky130_fd_sc_hs__dfxtp_4_5/a_696_458#
+ sky130_fd_sc_hs__dfxtp_4_5/a_544_485# sky130_fd_sc_hs__dfxtp_4_5/a_1178_124# sky130_fd_sc_hs__dfxtp_4_5/a_1034_424#
+ sky130_fd_sc_hs__dfxtp_4
Xsky130_fd_sc_hs__buf_2_11 DVSS DVDD DVDD DVSS clk_prbs sky130_fd_sc_hs__buf_2_11/X
+ sky130_fd_sc_hs__buf_2_11/a_21_260# sky130_fd_sc_hs__buf_2
Xsky130_fd_sc_hs__clkbuf_2_5 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__dfxtp_4_5/D din[13]
+ sky130_fd_sc_hs__clkbuf_2_5/a_43_192# sky130_fd_sc_hs__clkbuf_2
Xsky130_fd_sc_hs__clkbuf_2_27 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__dfxtp_4_46/D din[0]
+ sky130_fd_sc_hs__clkbuf_2_27/a_43_192# sky130_fd_sc_hs__clkbuf_2
Xsky130_fd_sc_hs__a22o_1_16 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__a22o_1_17/X sky130_fd_sc_hs__dfxtp_4_27/Q
+ sky130_fd_sc_hs__inv_4_13/Y sky130_fd_sc_hs__dfxtp_4_23/Q sky130_fd_sc_hs__buf_2_9/X
+ sky130_fd_sc_hs__a22o_1_17/a_222_392# sky130_fd_sc_hs__a22o_1_17/a_230_79# sky130_fd_sc_hs__a22o_1_17/a_52_123#
+ sky130_fd_sc_hs__a22o_1_17/a_132_392# sky130_fd_sc_hs__a22o_1
Xsky130_fd_sc_hs__clkbuf_2_16 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__dfxtp_4_23/D din[7]
+ sky130_fd_sc_hs__clkbuf_2_17/a_43_192# sky130_fd_sc_hs__clkbuf_2
Xsky130_fd_sc_hs__buf_2_7 DVSS DVDD DVDD DVSS clk_prbs sky130_fd_sc_hs__buf_2_7/X
+ sky130_fd_sc_hs__buf_2_7/a_21_260# sky130_fd_sc_hs__buf_2
Xsky130_fd_sc_hs__dfxtp_4_6 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__dfxtp_4_7/Q sky130_fd_sc_hs__a22o_1_3/X
+ sky130_fd_sc_hs__inv_4_19/A sky130_fd_sc_hs__dfxtp_4_7/a_1226_296# sky130_fd_sc_hs__dfxtp_4_7/a_735_102#
+ sky130_fd_sc_hs__dfxtp_4_7/a_1141_508# sky130_fd_sc_hs__dfxtp_4_7/a_206_368# sky130_fd_sc_hs__dfxtp_4_7/a_437_503#
+ sky130_fd_sc_hs__dfxtp_4_7/a_27_74# sky130_fd_sc_hs__dfxtp_4_7/a_651_503# sky130_fd_sc_hs__dfxtp_4_7/a_696_458#
+ sky130_fd_sc_hs__dfxtp_4_7/a_544_485# sky130_fd_sc_hs__dfxtp_4_7/a_1178_124# sky130_fd_sc_hs__dfxtp_4_7/a_1034_424#
+ sky130_fd_sc_hs__dfxtp_4
Xsky130_fd_sc_hs__buf_2_12 DVSS DVDD DVDD DVSS clk_prbs sky130_fd_sc_hs__buf_2_14/X
+ sky130_fd_sc_hs__buf_2_14/a_21_260# sky130_fd_sc_hs__buf_2
Xsky130_fd_sc_hs__clkbuf_2_6 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__dfxtp_4_9/D din[12]
+ sky130_fd_sc_hs__clkbuf_2_7/a_43_192# sky130_fd_sc_hs__clkbuf_2
Xsky130_fd_sc_hs__clkbuf_2_28 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__dfxtp_4_45/D din[1]
+ sky130_fd_sc_hs__clkbuf_2_29/a_43_192# sky130_fd_sc_hs__clkbuf_2
Xsky130_fd_sc_hs__a22o_1_17 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__a22o_1_17/X sky130_fd_sc_hs__dfxtp_4_27/Q
+ sky130_fd_sc_hs__inv_4_13/Y sky130_fd_sc_hs__dfxtp_4_23/Q sky130_fd_sc_hs__buf_2_9/X
+ sky130_fd_sc_hs__a22o_1_17/a_222_392# sky130_fd_sc_hs__a22o_1_17/a_230_79# sky130_fd_sc_hs__a22o_1_17/a_52_123#
+ sky130_fd_sc_hs__a22o_1_17/a_132_392# sky130_fd_sc_hs__a22o_1
Xsky130_fd_sc_hs__clkbuf_2_17 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__dfxtp_4_23/D din[7]
+ sky130_fd_sc_hs__clkbuf_2_17/a_43_192# sky130_fd_sc_hs__clkbuf_2
Xsky130_fd_sc_hs__buf_2_8 DVSS DVDD DVDD DVSS clk_prbs sky130_fd_sc_hs__buf_2_9/X
+ sky130_fd_sc_hs__buf_2_9/a_21_260# sky130_fd_sc_hs__buf_2
Xsky130_fd_sc_hs__dfxtp_4_7 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__dfxtp_4_7/Q sky130_fd_sc_hs__a22o_1_3/X
+ sky130_fd_sc_hs__inv_4_19/A sky130_fd_sc_hs__dfxtp_4_7/a_1226_296# sky130_fd_sc_hs__dfxtp_4_7/a_735_102#
+ sky130_fd_sc_hs__dfxtp_4_7/a_1141_508# sky130_fd_sc_hs__dfxtp_4_7/a_206_368# sky130_fd_sc_hs__dfxtp_4_7/a_437_503#
+ sky130_fd_sc_hs__dfxtp_4_7/a_27_74# sky130_fd_sc_hs__dfxtp_4_7/a_651_503# sky130_fd_sc_hs__dfxtp_4_7/a_696_458#
+ sky130_fd_sc_hs__dfxtp_4_7/a_544_485# sky130_fd_sc_hs__dfxtp_4_7/a_1178_124# sky130_fd_sc_hs__dfxtp_4_7/a_1034_424#
+ sky130_fd_sc_hs__dfxtp_4
Xsky130_fd_sc_hs__buf_2_13 DVSS DVDD DVDD DVSS clk_prbs sky130_fd_sc_hs__buf_2_15/X
+ sky130_fd_sc_hs__buf_2_15/a_21_260# sky130_fd_sc_hs__buf_2
Xsky130_fd_sc_hs__dfrtp_4_0 DVSS DVDD sky130_fd_sc_hs__clkinv_2_1/Y DVDD DVSS sky130_fd_sc_hs__inv_4_19/Y
+ clk sky130_fd_sc_hs__dfrtp_4_1/Q sky130_fd_sc_hs__dfrtp_4_1/a_37_78# sky130_fd_sc_hs__dfrtp_4_1/a_494_366#
+ sky130_fd_sc_hs__dfrtp_4_1/a_699_463# sky130_fd_sc_hs__dfrtp_4_1/a_313_74# sky130_fd_sc_hs__dfrtp_4_1/a_1627_493#
+ sky130_fd_sc_hs__dfrtp_4_1/a_1678_395# sky130_fd_sc_hs__dfrtp_4_1/a_1827_81# sky130_fd_sc_hs__dfrtp_4_1/a_789_463#
+ sky130_fd_sc_hs__dfrtp_4_1/a_1350_392# sky130_fd_sc_hs__dfrtp_4_1/a_834_355# sky130_fd_sc_hs__dfrtp_4_1/a_812_138#
+ sky130_fd_sc_hs__dfrtp_4_1/a_124_78# sky130_fd_sc_hs__dfrtp_4_1/a_1647_81# sky130_fd_sc_hs__dfrtp_4_1/a_2010_409#
+ sky130_fd_sc_hs__dfrtp_4_1/a_890_138# sky130_fd_sc_hs__dfrtp_4
Xsky130_fd_sc_hs__clkbuf_2_7 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__dfxtp_4_9/D din[12]
+ sky130_fd_sc_hs__clkbuf_2_7/a_43_192# sky130_fd_sc_hs__clkbuf_2
Xsky130_fd_sc_hs__clkbuf_2_29 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__dfxtp_4_45/D din[1]
+ sky130_fd_sc_hs__clkbuf_2_29/a_43_192# sky130_fd_sc_hs__clkbuf_2
Xsky130_fd_sc_hs__a22o_1_18 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__a22o_1_19/X sky130_fd_sc_hs__dfxtp_4_35/Q
+ sky130_fd_sc_hs__inv_4_15/Y sky130_fd_sc_hs__dfxtp_4_31/Q sky130_fd_sc_hs__buf_2_11/X
+ sky130_fd_sc_hs__a22o_1_19/a_222_392# sky130_fd_sc_hs__a22o_1_19/a_230_79# sky130_fd_sc_hs__a22o_1_19/a_52_123#
+ sky130_fd_sc_hs__a22o_1_19/a_132_392# sky130_fd_sc_hs__a22o_1
Xsky130_fd_sc_hs__clkbuf_2_18 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__dfxtp_4_27/D din[6]
+ sky130_fd_sc_hs__clkbuf_2_19/a_43_192# sky130_fd_sc_hs__clkbuf_2
Xsky130_fd_sc_hs__dfxtp_4_8 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__dfxtp_4_8/Q sky130_fd_sc_hs__dfxtp_4_8/D
+ sky130_fd_sc_hs__clkbuf_4_1/X sky130_fd_sc_hs__dfxtp_4_8/a_1226_296# sky130_fd_sc_hs__dfxtp_4_8/a_735_102#
+ sky130_fd_sc_hs__dfxtp_4_8/a_1141_508# sky130_fd_sc_hs__dfxtp_4_8/a_206_368# sky130_fd_sc_hs__dfxtp_4_8/a_437_503#
+ sky130_fd_sc_hs__dfxtp_4_8/a_27_74# sky130_fd_sc_hs__dfxtp_4_8/a_651_503# sky130_fd_sc_hs__dfxtp_4_8/a_696_458#
+ sky130_fd_sc_hs__dfxtp_4_8/a_544_485# sky130_fd_sc_hs__dfxtp_4_8/a_1178_124# sky130_fd_sc_hs__dfxtp_4_8/a_1034_424#
+ sky130_fd_sc_hs__dfxtp_4
Xsky130_fd_sc_hs__buf_2_9 DVSS DVDD DVDD DVSS clk_prbs sky130_fd_sc_hs__buf_2_9/X
+ sky130_fd_sc_hs__buf_2_9/a_21_260# sky130_fd_sc_hs__buf_2
Xsky130_fd_sc_hs__buf_2_14 DVSS DVDD DVDD DVSS clk_prbs sky130_fd_sc_hs__buf_2_14/X
+ sky130_fd_sc_hs__buf_2_14/a_21_260# sky130_fd_sc_hs__buf_2
Xsky130_fd_sc_hs__dfrtp_4_1 DVSS DVDD sky130_fd_sc_hs__clkinv_2_1/Y DVDD DVSS sky130_fd_sc_hs__inv_4_19/Y
+ clk sky130_fd_sc_hs__dfrtp_4_1/Q sky130_fd_sc_hs__dfrtp_4_1/a_37_78# sky130_fd_sc_hs__dfrtp_4_1/a_494_366#
+ sky130_fd_sc_hs__dfrtp_4_1/a_699_463# sky130_fd_sc_hs__dfrtp_4_1/a_313_74# sky130_fd_sc_hs__dfrtp_4_1/a_1627_493#
+ sky130_fd_sc_hs__dfrtp_4_1/a_1678_395# sky130_fd_sc_hs__dfrtp_4_1/a_1827_81# sky130_fd_sc_hs__dfrtp_4_1/a_789_463#
+ sky130_fd_sc_hs__dfrtp_4_1/a_1350_392# sky130_fd_sc_hs__dfrtp_4_1/a_834_355# sky130_fd_sc_hs__dfrtp_4_1/a_812_138#
+ sky130_fd_sc_hs__dfrtp_4_1/a_124_78# sky130_fd_sc_hs__dfrtp_4_1/a_1647_81# sky130_fd_sc_hs__dfrtp_4_1/a_2010_409#
+ sky130_fd_sc_hs__dfrtp_4_1/a_890_138# sky130_fd_sc_hs__dfrtp_4
Xsky130_fd_sc_hs__clkbuf_2_8 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__dfxtp_4_15/D din[9]
+ sky130_fd_sc_hs__clkbuf_2_9/a_43_192# sky130_fd_sc_hs__clkbuf_2
Xsky130_fd_sc_hs__a22o_1_19 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__a22o_1_19/X sky130_fd_sc_hs__dfxtp_4_35/Q
+ sky130_fd_sc_hs__inv_4_15/Y sky130_fd_sc_hs__dfxtp_4_31/Q sky130_fd_sc_hs__buf_2_11/X
+ sky130_fd_sc_hs__a22o_1_19/a_222_392# sky130_fd_sc_hs__a22o_1_19/a_230_79# sky130_fd_sc_hs__a22o_1_19/a_52_123#
+ sky130_fd_sc_hs__a22o_1_19/a_132_392# sky130_fd_sc_hs__a22o_1
Xsky130_fd_sc_hs__clkbuf_2_19 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__dfxtp_4_27/D din[6]
+ sky130_fd_sc_hs__clkbuf_2_19/a_43_192# sky130_fd_sc_hs__clkbuf_2
Xsky130_fd_sc_hs__dfxtp_4_9 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__dfxtp_4_9/Q sky130_fd_sc_hs__dfxtp_4_9/D
+ sky130_fd_sc_hs__clkbuf_4_1/X sky130_fd_sc_hs__dfxtp_4_9/a_1226_296# sky130_fd_sc_hs__dfxtp_4_9/a_735_102#
+ sky130_fd_sc_hs__dfxtp_4_9/a_1141_508# sky130_fd_sc_hs__dfxtp_4_9/a_206_368# sky130_fd_sc_hs__dfxtp_4_9/a_437_503#
+ sky130_fd_sc_hs__dfxtp_4_9/a_27_74# sky130_fd_sc_hs__dfxtp_4_9/a_651_503# sky130_fd_sc_hs__dfxtp_4_9/a_696_458#
+ sky130_fd_sc_hs__dfxtp_4_9/a_544_485# sky130_fd_sc_hs__dfxtp_4_9/a_1178_124# sky130_fd_sc_hs__dfxtp_4_9/a_1034_424#
+ sky130_fd_sc_hs__dfxtp_4
Xsky130_fd_sc_hs__buf_2_15 DVSS DVDD DVDD DVSS clk_prbs sky130_fd_sc_hs__buf_2_15/X
+ sky130_fd_sc_hs__buf_2_15/a_21_260# sky130_fd_sc_hs__buf_2
Xsky130_fd_sc_hs__dfrtp_4_2 DVSS DVDD sky130_fd_sc_hs__inv_4_7/Y DVDD DVSS sky130_fd_sc_hs__inv_4_11/Y
+ sky130_fd_sc_hs__clkinv_4_1/Y sky130_fd_sc_hs__inv_4_11/A sky130_fd_sc_hs__dfrtp_4_3/a_37_78#
+ sky130_fd_sc_hs__dfrtp_4_3/a_494_366# sky130_fd_sc_hs__dfrtp_4_3/a_699_463# sky130_fd_sc_hs__dfrtp_4_3/a_313_74#
+ sky130_fd_sc_hs__dfrtp_4_3/a_1627_493# sky130_fd_sc_hs__dfrtp_4_3/a_1678_395# sky130_fd_sc_hs__dfrtp_4_3/a_1827_81#
+ sky130_fd_sc_hs__dfrtp_4_3/a_789_463# sky130_fd_sc_hs__dfrtp_4_3/a_1350_392# sky130_fd_sc_hs__dfrtp_4_3/a_834_355#
+ sky130_fd_sc_hs__dfrtp_4_3/a_812_138# sky130_fd_sc_hs__dfrtp_4_3/a_124_78# sky130_fd_sc_hs__dfrtp_4_3/a_1647_81#
+ sky130_fd_sc_hs__dfrtp_4_3/a_2010_409# sky130_fd_sc_hs__dfrtp_4_3/a_890_138# sky130_fd_sc_hs__dfrtp_4
Xsky130_fd_sc_hs__clkbuf_2_9 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__dfxtp_4_15/D din[9]
+ sky130_fd_sc_hs__clkbuf_2_9/a_43_192# sky130_fd_sc_hs__clkbuf_2
Xsky130_fd_sc_hs__dfrtp_4_3 DVSS DVDD sky130_fd_sc_hs__inv_4_7/Y DVDD DVSS sky130_fd_sc_hs__inv_4_11/Y
+ sky130_fd_sc_hs__clkinv_4_1/Y sky130_fd_sc_hs__inv_4_11/A sky130_fd_sc_hs__dfrtp_4_3/a_37_78#
+ sky130_fd_sc_hs__dfrtp_4_3/a_494_366# sky130_fd_sc_hs__dfrtp_4_3/a_699_463# sky130_fd_sc_hs__dfrtp_4_3/a_313_74#
+ sky130_fd_sc_hs__dfrtp_4_3/a_1627_493# sky130_fd_sc_hs__dfrtp_4_3/a_1678_395# sky130_fd_sc_hs__dfrtp_4_3/a_1827_81#
+ sky130_fd_sc_hs__dfrtp_4_3/a_789_463# sky130_fd_sc_hs__dfrtp_4_3/a_1350_392# sky130_fd_sc_hs__dfrtp_4_3/a_834_355#
+ sky130_fd_sc_hs__dfrtp_4_3/a_812_138# sky130_fd_sc_hs__dfrtp_4_3/a_124_78# sky130_fd_sc_hs__dfrtp_4_3/a_1647_81#
+ sky130_fd_sc_hs__dfrtp_4_3/a_2010_409# sky130_fd_sc_hs__dfrtp_4_3/a_890_138# sky130_fd_sc_hs__dfrtp_4
Xsky130_fd_sc_hs__inv_4_20 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_21/Y clk_prbs
+ sky130_fd_sc_hs__inv_4
Xsky130_fd_sc_hs__inv_4_21 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_21/Y clk_prbs
+ sky130_fd_sc_hs__inv_4
Xsky130_fd_sc_hs__inv_4_10 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_11/Y sky130_fd_sc_hs__inv_4_11/A
+ sky130_fd_sc_hs__inv_4
Xsky130_fd_sc_hs__inv_4_11 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_11/Y sky130_fd_sc_hs__inv_4_11/A
+ sky130_fd_sc_hs__inv_4
Xsky130_fd_sc_hs__inv_4_12 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_13/Y clk_prbs
+ sky130_fd_sc_hs__inv_4
Xsky130_fd_sc_hs__inv_4_13 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_13/Y clk_prbs
+ sky130_fd_sc_hs__inv_4
Xsky130_fd_sc_hs__inv_4_14 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_15/Y clk_prbs
+ sky130_fd_sc_hs__inv_4
Xsky130_fd_sc_hs__a22o_1_0 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__a22o_1_1/X sky130_fd_sc_hs__dfxtp_4_1/Q
+ sky130_fd_sc_hs__inv_4_1/Y sky130_fd_sc_hs__dfxtp_4_3/Q sky130_fd_sc_hs__buf_2_1/X
+ sky130_fd_sc_hs__a22o_1_1/a_222_392# sky130_fd_sc_hs__a22o_1_1/a_230_79# sky130_fd_sc_hs__a22o_1_1/a_52_123#
+ sky130_fd_sc_hs__a22o_1_1/a_132_392# sky130_fd_sc_hs__a22o_1
Xsky130_fd_sc_hs__inv_4_15 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_15/Y clk_prbs
+ sky130_fd_sc_hs__inv_4
Xsky130_fd_sc_hs__inv_4_16 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_17/Y clk_prbs
+ sky130_fd_sc_hs__inv_4
Xsky130_fd_sc_hs__a22o_1_1 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__a22o_1_1/X sky130_fd_sc_hs__dfxtp_4_1/Q
+ sky130_fd_sc_hs__inv_4_1/Y sky130_fd_sc_hs__dfxtp_4_3/Q sky130_fd_sc_hs__buf_2_1/X
+ sky130_fd_sc_hs__a22o_1_1/a_222_392# sky130_fd_sc_hs__a22o_1_1/a_230_79# sky130_fd_sc_hs__a22o_1_1/a_52_123#
+ sky130_fd_sc_hs__a22o_1_1/a_132_392# sky130_fd_sc_hs__a22o_1
Xsky130_fd_sc_hs__inv_4_17 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_17/Y clk_prbs
+ sky130_fd_sc_hs__inv_4
Xsky130_fd_sc_hs__a22o_1_2 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__a22o_1_3/X sky130_fd_sc_hs__dfxtp_4_9/Q
+ sky130_fd_sc_hs__inv_4_3/Y sky130_fd_sc_hs__dfxtp_4_5/Q sky130_fd_sc_hs__buf_2_3/X
+ sky130_fd_sc_hs__a22o_1_3/a_222_392# sky130_fd_sc_hs__a22o_1_3/a_230_79# sky130_fd_sc_hs__a22o_1_3/a_52_123#
+ sky130_fd_sc_hs__a22o_1_3/a_132_392# sky130_fd_sc_hs__a22o_1
Xsky130_fd_sc_hs__clkbuf_1_0 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__clkinv_4_1/Y sky130_fd_sc_hs__a22o_1_9/B1
+ sky130_fd_sc_hs__clkbuf_1_1/a_27_74# sky130_fd_sc_hs__clkbuf_1
Xsky130_fd_sc_hs__inv_4_18 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_19/Y sky130_fd_sc_hs__inv_4_19/A
+ sky130_fd_sc_hs__inv_4
Xsky130_fd_sc_hs__a22o_1_3 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__a22o_1_3/X sky130_fd_sc_hs__dfxtp_4_9/Q
+ sky130_fd_sc_hs__inv_4_3/Y sky130_fd_sc_hs__dfxtp_4_5/Q sky130_fd_sc_hs__buf_2_3/X
+ sky130_fd_sc_hs__a22o_1_3/a_222_392# sky130_fd_sc_hs__a22o_1_3/a_230_79# sky130_fd_sc_hs__a22o_1_3/a_52_123#
+ sky130_fd_sc_hs__a22o_1_3/a_132_392# sky130_fd_sc_hs__a22o_1
Xsky130_fd_sc_hs__clkbuf_1_1 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__clkinv_4_1/Y sky130_fd_sc_hs__a22o_1_9/B1
+ sky130_fd_sc_hs__clkbuf_1_1/a_27_74# sky130_fd_sc_hs__clkbuf_1
Xsky130_fd_sc_hs__inv_4_19 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_19/Y sky130_fd_sc_hs__inv_4_19/A
+ sky130_fd_sc_hs__inv_4
Xsky130_fd_sc_hs__a22o_1_4 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__a22o_1_5/X sky130_fd_sc_hs__a22o_1_5/B2
+ sky130_fd_sc_hs__inv_4_5/Y sky130_fd_sc_hs__dfxtp_4_8/Q sky130_fd_sc_hs__buf_2_5/X
+ sky130_fd_sc_hs__a22o_1_5/a_222_392# sky130_fd_sc_hs__a22o_1_5/a_230_79# sky130_fd_sc_hs__a22o_1_5/a_52_123#
+ sky130_fd_sc_hs__a22o_1_5/a_132_392# sky130_fd_sc_hs__a22o_1
Xsky130_fd_sc_hs__a22o_1_5 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__a22o_1_5/X sky130_fd_sc_hs__a22o_1_5/B2
+ sky130_fd_sc_hs__inv_4_5/Y sky130_fd_sc_hs__dfxtp_4_8/Q sky130_fd_sc_hs__buf_2_5/X
+ sky130_fd_sc_hs__a22o_1_5/a_222_392# sky130_fd_sc_hs__a22o_1_5/a_230_79# sky130_fd_sc_hs__a22o_1_5/a_52_123#
+ sky130_fd_sc_hs__a22o_1_5/a_132_392# sky130_fd_sc_hs__a22o_1
Xsky130_fd_sc_hs__a22o_1_6 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__a22o_1_7/X sky130_fd_sc_hs__a22o_1_7/B2
+ sky130_fd_sc_hs__inv_4_9/Y sky130_fd_sc_hs__a22o_1_7/A2 sky130_fd_sc_hs__buf_2_7/X
+ sky130_fd_sc_hs__a22o_1_7/a_222_392# sky130_fd_sc_hs__a22o_1_7/a_230_79# sky130_fd_sc_hs__a22o_1_7/a_52_123#
+ sky130_fd_sc_hs__a22o_1_7/a_132_392# sky130_fd_sc_hs__a22o_1
Xsky130_fd_sc_hs__a22o_1_7 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__a22o_1_7/X sky130_fd_sc_hs__a22o_1_7/B2
+ sky130_fd_sc_hs__inv_4_9/Y sky130_fd_sc_hs__a22o_1_7/A2 sky130_fd_sc_hs__buf_2_7/X
+ sky130_fd_sc_hs__a22o_1_7/a_222_392# sky130_fd_sc_hs__a22o_1_7/a_230_79# sky130_fd_sc_hs__a22o_1_7/a_52_123#
+ sky130_fd_sc_hs__a22o_1_7/a_132_392# sky130_fd_sc_hs__a22o_1
Xsky130_fd_sc_hs__clkbuf_16_0 DVSS DVDD DVDD DVSS clk_prbs sky130_fd_sc_hs__inv_4_11/A
+ sky130_fd_sc_hs__clkbuf_16_1/a_114_74# sky130_fd_sc_hs__clkbuf_16
Xsky130_fd_sc_hs__a22o_1_8 DVSS DVDD DVDD DVSS dout[3] sky130_fd_sc_hs__dfxtp_4_7/Q
+ sky130_fd_sc_hs__a22o_1_9/B1 sky130_fd_sc_hs__a22o_1_9/A2 sky130_fd_sc_hs__inv_4_19/A
+ sky130_fd_sc_hs__a22o_1_9/a_222_392# sky130_fd_sc_hs__a22o_1_9/a_230_79# sky130_fd_sc_hs__a22o_1_9/a_52_123#
+ sky130_fd_sc_hs__a22o_1_9/a_132_392# sky130_fd_sc_hs__a22o_1
Xsky130_fd_sc_hs__clkbuf_16_1 DVSS DVDD DVDD DVSS clk_prbs sky130_fd_sc_hs__inv_4_11/A
+ sky130_fd_sc_hs__clkbuf_16_1/a_114_74# sky130_fd_sc_hs__clkbuf_16
Xsky130_fd_sc_hs__dfxtp_4_40 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__dfxtp_4_41/Q sky130_fd_sc_hs__a22o_1_23/X
+ sky130_fd_sc_hs__inv_4_19/A sky130_fd_sc_hs__dfxtp_4_41/a_1226_296# sky130_fd_sc_hs__dfxtp_4_41/a_735_102#
+ sky130_fd_sc_hs__dfxtp_4_41/a_1141_508# sky130_fd_sc_hs__dfxtp_4_41/a_206_368# sky130_fd_sc_hs__dfxtp_4_41/a_437_503#
+ sky130_fd_sc_hs__dfxtp_4_41/a_27_74# sky130_fd_sc_hs__dfxtp_4_41/a_651_503# sky130_fd_sc_hs__dfxtp_4_41/a_696_458#
+ sky130_fd_sc_hs__dfxtp_4_41/a_544_485# sky130_fd_sc_hs__dfxtp_4_41/a_1178_124# sky130_fd_sc_hs__dfxtp_4_41/a_1034_424#
+ sky130_fd_sc_hs__dfxtp_4
Xsky130_fd_sc_hs__a22o_1_9 DVSS DVDD DVDD DVSS dout[3] sky130_fd_sc_hs__dfxtp_4_7/Q
+ sky130_fd_sc_hs__a22o_1_9/B1 sky130_fd_sc_hs__a22o_1_9/A2 sky130_fd_sc_hs__inv_4_19/A
+ sky130_fd_sc_hs__a22o_1_9/a_222_392# sky130_fd_sc_hs__a22o_1_9/a_230_79# sky130_fd_sc_hs__a22o_1_9/a_52_123#
+ sky130_fd_sc_hs__a22o_1_9/a_132_392# sky130_fd_sc_hs__a22o_1
Xsky130_fd_sc_hs__dfxtp_4_41 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__dfxtp_4_41/Q sky130_fd_sc_hs__a22o_1_23/X
+ sky130_fd_sc_hs__inv_4_19/A sky130_fd_sc_hs__dfxtp_4_41/a_1226_296# sky130_fd_sc_hs__dfxtp_4_41/a_735_102#
+ sky130_fd_sc_hs__dfxtp_4_41/a_1141_508# sky130_fd_sc_hs__dfxtp_4_41/a_206_368# sky130_fd_sc_hs__dfxtp_4_41/a_437_503#
+ sky130_fd_sc_hs__dfxtp_4_41/a_27_74# sky130_fd_sc_hs__dfxtp_4_41/a_651_503# sky130_fd_sc_hs__dfxtp_4_41/a_696_458#
+ sky130_fd_sc_hs__dfxtp_4_41/a_544_485# sky130_fd_sc_hs__dfxtp_4_41/a_1178_124# sky130_fd_sc_hs__dfxtp_4_41/a_1034_424#
+ sky130_fd_sc_hs__dfxtp_4
Xsky130_fd_sc_hs__dfxtp_4_30 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__dfxtp_4_31/Q sky130_fd_sc_hs__dfxtp_4_31/D
+ sky130_fd_sc_hs__clkbuf_4_1/X sky130_fd_sc_hs__dfxtp_4_31/a_1226_296# sky130_fd_sc_hs__dfxtp_4_31/a_735_102#
+ sky130_fd_sc_hs__dfxtp_4_31/a_1141_508# sky130_fd_sc_hs__dfxtp_4_31/a_206_368# sky130_fd_sc_hs__dfxtp_4_31/a_437_503#
+ sky130_fd_sc_hs__dfxtp_4_31/a_27_74# sky130_fd_sc_hs__dfxtp_4_31/a_651_503# sky130_fd_sc_hs__dfxtp_4_31/a_696_458#
+ sky130_fd_sc_hs__dfxtp_4_31/a_544_485# sky130_fd_sc_hs__dfxtp_4_31/a_1178_124# sky130_fd_sc_hs__dfxtp_4_31/a_1034_424#
+ sky130_fd_sc_hs__dfxtp_4
Xsky130_fd_sc_hs__dfxtp_4_42 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__dfxtp_4_45/Q sky130_fd_sc_hs__dfxtp_4_45/D
+ sky130_fd_sc_hs__clkbuf_4_1/X sky130_fd_sc_hs__dfxtp_4_45/a_1226_296# sky130_fd_sc_hs__dfxtp_4_45/a_735_102#
+ sky130_fd_sc_hs__dfxtp_4_45/a_1141_508# sky130_fd_sc_hs__dfxtp_4_45/a_206_368# sky130_fd_sc_hs__dfxtp_4_45/a_437_503#
+ sky130_fd_sc_hs__dfxtp_4_45/a_27_74# sky130_fd_sc_hs__dfxtp_4_45/a_651_503# sky130_fd_sc_hs__dfxtp_4_45/a_696_458#
+ sky130_fd_sc_hs__dfxtp_4_45/a_544_485# sky130_fd_sc_hs__dfxtp_4_45/a_1178_124# sky130_fd_sc_hs__dfxtp_4_45/a_1034_424#
+ sky130_fd_sc_hs__dfxtp_4
Xsky130_fd_sc_hs__dfxtp_4_31 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__dfxtp_4_31/Q sky130_fd_sc_hs__dfxtp_4_31/D
+ sky130_fd_sc_hs__clkbuf_4_1/X sky130_fd_sc_hs__dfxtp_4_31/a_1226_296# sky130_fd_sc_hs__dfxtp_4_31/a_735_102#
+ sky130_fd_sc_hs__dfxtp_4_31/a_1141_508# sky130_fd_sc_hs__dfxtp_4_31/a_206_368# sky130_fd_sc_hs__dfxtp_4_31/a_437_503#
+ sky130_fd_sc_hs__dfxtp_4_31/a_27_74# sky130_fd_sc_hs__dfxtp_4_31/a_651_503# sky130_fd_sc_hs__dfxtp_4_31/a_696_458#
+ sky130_fd_sc_hs__dfxtp_4_31/a_544_485# sky130_fd_sc_hs__dfxtp_4_31/a_1178_124# sky130_fd_sc_hs__dfxtp_4_31/a_1034_424#
+ sky130_fd_sc_hs__dfxtp_4
Xsky130_fd_sc_hs__dfxtp_4_20 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__dfxtp_4_23/Q sky130_fd_sc_hs__dfxtp_4_23/D
+ sky130_fd_sc_hs__clkbuf_4_1/X sky130_fd_sc_hs__dfxtp_4_23/a_1226_296# sky130_fd_sc_hs__dfxtp_4_23/a_735_102#
+ sky130_fd_sc_hs__dfxtp_4_23/a_1141_508# sky130_fd_sc_hs__dfxtp_4_23/a_206_368# sky130_fd_sc_hs__dfxtp_4_23/a_437_503#
+ sky130_fd_sc_hs__dfxtp_4_23/a_27_74# sky130_fd_sc_hs__dfxtp_4_23/a_651_503# sky130_fd_sc_hs__dfxtp_4_23/a_696_458#
+ sky130_fd_sc_hs__dfxtp_4_23/a_544_485# sky130_fd_sc_hs__dfxtp_4_23/a_1178_124# sky130_fd_sc_hs__dfxtp_4_23/a_1034_424#
+ sky130_fd_sc_hs__dfxtp_4
Xsky130_fd_sc_hs__dfxtp_4_10 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__dfxtp_4_8/Q sky130_fd_sc_hs__dfxtp_4_8/D
+ sky130_fd_sc_hs__clkbuf_4_1/X sky130_fd_sc_hs__dfxtp_4_8/a_1226_296# sky130_fd_sc_hs__dfxtp_4_8/a_735_102#
+ sky130_fd_sc_hs__dfxtp_4_8/a_1141_508# sky130_fd_sc_hs__dfxtp_4_8/a_206_368# sky130_fd_sc_hs__dfxtp_4_8/a_437_503#
+ sky130_fd_sc_hs__dfxtp_4_8/a_27_74# sky130_fd_sc_hs__dfxtp_4_8/a_651_503# sky130_fd_sc_hs__dfxtp_4_8/a_696_458#
+ sky130_fd_sc_hs__dfxtp_4_8/a_544_485# sky130_fd_sc_hs__dfxtp_4_8/a_1178_124# sky130_fd_sc_hs__dfxtp_4_8/a_1034_424#
+ sky130_fd_sc_hs__dfxtp_4
Xsky130_fd_sc_hs__dfxtp_4_43 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__dfxtp_4_46/Q sky130_fd_sc_hs__dfxtp_4_46/D
+ sky130_fd_sc_hs__clkbuf_4_1/X sky130_fd_sc_hs__dfxtp_4_46/a_1226_296# sky130_fd_sc_hs__dfxtp_4_46/a_735_102#
+ sky130_fd_sc_hs__dfxtp_4_46/a_1141_508# sky130_fd_sc_hs__dfxtp_4_46/a_206_368# sky130_fd_sc_hs__dfxtp_4_46/a_437_503#
+ sky130_fd_sc_hs__dfxtp_4_46/a_27_74# sky130_fd_sc_hs__dfxtp_4_46/a_651_503# sky130_fd_sc_hs__dfxtp_4_46/a_696_458#
+ sky130_fd_sc_hs__dfxtp_4_46/a_544_485# sky130_fd_sc_hs__dfxtp_4_46/a_1178_124# sky130_fd_sc_hs__dfxtp_4_46/a_1034_424#
+ sky130_fd_sc_hs__dfxtp_4
Xsky130_fd_sc_hs__dfxtp_4_32 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__dfxtp_4_33/Q sky130_fd_sc_hs__a22o_1_21/X
+ sky130_fd_sc_hs__inv_4_19/A sky130_fd_sc_hs__dfxtp_4_33/a_1226_296# sky130_fd_sc_hs__dfxtp_4_33/a_735_102#
+ sky130_fd_sc_hs__dfxtp_4_33/a_1141_508# sky130_fd_sc_hs__dfxtp_4_33/a_206_368# sky130_fd_sc_hs__dfxtp_4_33/a_437_503#
+ sky130_fd_sc_hs__dfxtp_4_33/a_27_74# sky130_fd_sc_hs__dfxtp_4_33/a_651_503# sky130_fd_sc_hs__dfxtp_4_33/a_696_458#
+ sky130_fd_sc_hs__dfxtp_4_33/a_544_485# sky130_fd_sc_hs__dfxtp_4_33/a_1178_124# sky130_fd_sc_hs__dfxtp_4_33/a_1034_424#
+ sky130_fd_sc_hs__dfxtp_4
Xsky130_fd_sc_hs__dfxtp_4_21 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__a22o_1_5/B2 sky130_fd_sc_hs__dfxtp_4_24/D
+ sky130_fd_sc_hs__clkbuf_4_1/X sky130_fd_sc_hs__dfxtp_4_24/a_1226_296# sky130_fd_sc_hs__dfxtp_4_24/a_735_102#
+ sky130_fd_sc_hs__dfxtp_4_24/a_1141_508# sky130_fd_sc_hs__dfxtp_4_24/a_206_368# sky130_fd_sc_hs__dfxtp_4_24/a_437_503#
+ sky130_fd_sc_hs__dfxtp_4_24/a_27_74# sky130_fd_sc_hs__dfxtp_4_24/a_651_503# sky130_fd_sc_hs__dfxtp_4_24/a_696_458#
+ sky130_fd_sc_hs__dfxtp_4_24/a_544_485# sky130_fd_sc_hs__dfxtp_4_24/a_1178_124# sky130_fd_sc_hs__dfxtp_4_24/a_1034_424#
+ sky130_fd_sc_hs__dfxtp_4
Xsky130_fd_sc_hs__dfxtp_4_11 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__dfxtp_4_9/Q sky130_fd_sc_hs__dfxtp_4_9/D
+ sky130_fd_sc_hs__clkbuf_4_1/X sky130_fd_sc_hs__dfxtp_4_9/a_1226_296# sky130_fd_sc_hs__dfxtp_4_9/a_735_102#
+ sky130_fd_sc_hs__dfxtp_4_9/a_1141_508# sky130_fd_sc_hs__dfxtp_4_9/a_206_368# sky130_fd_sc_hs__dfxtp_4_9/a_437_503#
+ sky130_fd_sc_hs__dfxtp_4_9/a_27_74# sky130_fd_sc_hs__dfxtp_4_9/a_651_503# sky130_fd_sc_hs__dfxtp_4_9/a_696_458#
+ sky130_fd_sc_hs__dfxtp_4_9/a_544_485# sky130_fd_sc_hs__dfxtp_4_9/a_1178_124# sky130_fd_sc_hs__dfxtp_4_9/a_1034_424#
+ sky130_fd_sc_hs__dfxtp_4
Xsky130_fd_sc_hs__dfxtp_4_44 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__dfxtp_4_47/Q sky130_fd_sc_hs__dfxtp_4_47/D
+ sky130_fd_sc_hs__clkbuf_4_1/X sky130_fd_sc_hs__dfxtp_4_47/a_1226_296# sky130_fd_sc_hs__dfxtp_4_47/a_735_102#
+ sky130_fd_sc_hs__dfxtp_4_47/a_1141_508# sky130_fd_sc_hs__dfxtp_4_47/a_206_368# sky130_fd_sc_hs__dfxtp_4_47/a_437_503#
+ sky130_fd_sc_hs__dfxtp_4_47/a_27_74# sky130_fd_sc_hs__dfxtp_4_47/a_651_503# sky130_fd_sc_hs__dfxtp_4_47/a_696_458#
+ sky130_fd_sc_hs__dfxtp_4_47/a_544_485# sky130_fd_sc_hs__dfxtp_4_47/a_1178_124# sky130_fd_sc_hs__dfxtp_4_47/a_1034_424#
+ sky130_fd_sc_hs__dfxtp_4
Xsky130_fd_sc_hs__dfxtp_4_33 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__dfxtp_4_33/Q sky130_fd_sc_hs__a22o_1_21/X
+ sky130_fd_sc_hs__inv_4_19/A sky130_fd_sc_hs__dfxtp_4_33/a_1226_296# sky130_fd_sc_hs__dfxtp_4_33/a_735_102#
+ sky130_fd_sc_hs__dfxtp_4_33/a_1141_508# sky130_fd_sc_hs__dfxtp_4_33/a_206_368# sky130_fd_sc_hs__dfxtp_4_33/a_437_503#
+ sky130_fd_sc_hs__dfxtp_4_33/a_27_74# sky130_fd_sc_hs__dfxtp_4_33/a_651_503# sky130_fd_sc_hs__dfxtp_4_33/a_696_458#
+ sky130_fd_sc_hs__dfxtp_4_33/a_544_485# sky130_fd_sc_hs__dfxtp_4_33/a_1178_124# sky130_fd_sc_hs__dfxtp_4_33/a_1034_424#
+ sky130_fd_sc_hs__dfxtp_4
Xsky130_fd_sc_hs__dfxtp_4_22 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__a22o_1_7/B2 sky130_fd_sc_hs__dfxtp_4_25/D
+ sky130_fd_sc_hs__clkbuf_4_1/X sky130_fd_sc_hs__dfxtp_4_25/a_1226_296# sky130_fd_sc_hs__dfxtp_4_25/a_735_102#
+ sky130_fd_sc_hs__dfxtp_4_25/a_1141_508# sky130_fd_sc_hs__dfxtp_4_25/a_206_368# sky130_fd_sc_hs__dfxtp_4_25/a_437_503#
+ sky130_fd_sc_hs__dfxtp_4_25/a_27_74# sky130_fd_sc_hs__dfxtp_4_25/a_651_503# sky130_fd_sc_hs__dfxtp_4_25/a_696_458#
+ sky130_fd_sc_hs__dfxtp_4_25/a_544_485# sky130_fd_sc_hs__dfxtp_4_25/a_1178_124# sky130_fd_sc_hs__dfxtp_4_25/a_1034_424#
+ sky130_fd_sc_hs__dfxtp_4
Xsky130_fd_sc_hs__dfxtp_4_12 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__a22o_1_9/A2 sky130_fd_sc_hs__a22o_1_1/X
+ sky130_fd_sc_hs__inv_4_19/A sky130_fd_sc_hs__dfxtp_4_13/a_1226_296# sky130_fd_sc_hs__dfxtp_4_13/a_735_102#
+ sky130_fd_sc_hs__dfxtp_4_13/a_1141_508# sky130_fd_sc_hs__dfxtp_4_13/a_206_368# sky130_fd_sc_hs__dfxtp_4_13/a_437_503#
+ sky130_fd_sc_hs__dfxtp_4_13/a_27_74# sky130_fd_sc_hs__dfxtp_4_13/a_651_503# sky130_fd_sc_hs__dfxtp_4_13/a_696_458#
+ sky130_fd_sc_hs__dfxtp_4_13/a_544_485# sky130_fd_sc_hs__dfxtp_4_13/a_1178_124# sky130_fd_sc_hs__dfxtp_4_13/a_1034_424#
+ sky130_fd_sc_hs__dfxtp_4
Xsky130_fd_sc_hs__dfxtp_4_45 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__dfxtp_4_45/Q sky130_fd_sc_hs__dfxtp_4_45/D
+ sky130_fd_sc_hs__clkbuf_4_1/X sky130_fd_sc_hs__dfxtp_4_45/a_1226_296# sky130_fd_sc_hs__dfxtp_4_45/a_735_102#
+ sky130_fd_sc_hs__dfxtp_4_45/a_1141_508# sky130_fd_sc_hs__dfxtp_4_45/a_206_368# sky130_fd_sc_hs__dfxtp_4_45/a_437_503#
+ sky130_fd_sc_hs__dfxtp_4_45/a_27_74# sky130_fd_sc_hs__dfxtp_4_45/a_651_503# sky130_fd_sc_hs__dfxtp_4_45/a_696_458#
+ sky130_fd_sc_hs__dfxtp_4_45/a_544_485# sky130_fd_sc_hs__dfxtp_4_45/a_1178_124# sky130_fd_sc_hs__dfxtp_4_45/a_1034_424#
+ sky130_fd_sc_hs__dfxtp_4
Xsky130_fd_sc_hs__dfxtp_4_34 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__dfxtp_4_35/Q sky130_fd_sc_hs__dfxtp_4_35/D
+ sky130_fd_sc_hs__clkbuf_4_1/X sky130_fd_sc_hs__dfxtp_4_35/a_1226_296# sky130_fd_sc_hs__dfxtp_4_35/a_735_102#
+ sky130_fd_sc_hs__dfxtp_4_35/a_1141_508# sky130_fd_sc_hs__dfxtp_4_35/a_206_368# sky130_fd_sc_hs__dfxtp_4_35/a_437_503#
+ sky130_fd_sc_hs__dfxtp_4_35/a_27_74# sky130_fd_sc_hs__dfxtp_4_35/a_651_503# sky130_fd_sc_hs__dfxtp_4_35/a_696_458#
+ sky130_fd_sc_hs__dfxtp_4_35/a_544_485# sky130_fd_sc_hs__dfxtp_4_35/a_1178_124# sky130_fd_sc_hs__dfxtp_4_35/a_1034_424#
+ sky130_fd_sc_hs__dfxtp_4
Xsky130_fd_sc_hs__dfxtp_4_23 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__dfxtp_4_23/Q sky130_fd_sc_hs__dfxtp_4_23/D
+ sky130_fd_sc_hs__clkbuf_4_1/X sky130_fd_sc_hs__dfxtp_4_23/a_1226_296# sky130_fd_sc_hs__dfxtp_4_23/a_735_102#
+ sky130_fd_sc_hs__dfxtp_4_23/a_1141_508# sky130_fd_sc_hs__dfxtp_4_23/a_206_368# sky130_fd_sc_hs__dfxtp_4_23/a_437_503#
+ sky130_fd_sc_hs__dfxtp_4_23/a_27_74# sky130_fd_sc_hs__dfxtp_4_23/a_651_503# sky130_fd_sc_hs__dfxtp_4_23/a_696_458#
+ sky130_fd_sc_hs__dfxtp_4_23/a_544_485# sky130_fd_sc_hs__dfxtp_4_23/a_1178_124# sky130_fd_sc_hs__dfxtp_4_23/a_1034_424#
+ sky130_fd_sc_hs__dfxtp_4
Xsky130_fd_sc_hs__inv_4_0 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_1/Y clk_prbs
+ sky130_fd_sc_hs__inv_4
Xsky130_fd_sc_hs__dfxtp_4_13 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__a22o_1_9/A2 sky130_fd_sc_hs__a22o_1_1/X
+ sky130_fd_sc_hs__inv_4_19/A sky130_fd_sc_hs__dfxtp_4_13/a_1226_296# sky130_fd_sc_hs__dfxtp_4_13/a_735_102#
+ sky130_fd_sc_hs__dfxtp_4_13/a_1141_508# sky130_fd_sc_hs__dfxtp_4_13/a_206_368# sky130_fd_sc_hs__dfxtp_4_13/a_437_503#
+ sky130_fd_sc_hs__dfxtp_4_13/a_27_74# sky130_fd_sc_hs__dfxtp_4_13/a_651_503# sky130_fd_sc_hs__dfxtp_4_13/a_696_458#
+ sky130_fd_sc_hs__dfxtp_4_13/a_544_485# sky130_fd_sc_hs__dfxtp_4_13/a_1178_124# sky130_fd_sc_hs__dfxtp_4_13/a_1034_424#
+ sky130_fd_sc_hs__dfxtp_4
Xsky130_fd_sc_hs__dfxtp_4_46 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__dfxtp_4_46/Q sky130_fd_sc_hs__dfxtp_4_46/D
+ sky130_fd_sc_hs__clkbuf_4_1/X sky130_fd_sc_hs__dfxtp_4_46/a_1226_296# sky130_fd_sc_hs__dfxtp_4_46/a_735_102#
+ sky130_fd_sc_hs__dfxtp_4_46/a_1141_508# sky130_fd_sc_hs__dfxtp_4_46/a_206_368# sky130_fd_sc_hs__dfxtp_4_46/a_437_503#
+ sky130_fd_sc_hs__dfxtp_4_46/a_27_74# sky130_fd_sc_hs__dfxtp_4_46/a_651_503# sky130_fd_sc_hs__dfxtp_4_46/a_696_458#
+ sky130_fd_sc_hs__dfxtp_4_46/a_544_485# sky130_fd_sc_hs__dfxtp_4_46/a_1178_124# sky130_fd_sc_hs__dfxtp_4_46/a_1034_424#
+ sky130_fd_sc_hs__dfxtp_4
Xsky130_fd_sc_hs__dfxtp_4_35 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__dfxtp_4_35/Q sky130_fd_sc_hs__dfxtp_4_35/D
+ sky130_fd_sc_hs__clkbuf_4_1/X sky130_fd_sc_hs__dfxtp_4_35/a_1226_296# sky130_fd_sc_hs__dfxtp_4_35/a_735_102#
+ sky130_fd_sc_hs__dfxtp_4_35/a_1141_508# sky130_fd_sc_hs__dfxtp_4_35/a_206_368# sky130_fd_sc_hs__dfxtp_4_35/a_437_503#
+ sky130_fd_sc_hs__dfxtp_4_35/a_27_74# sky130_fd_sc_hs__dfxtp_4_35/a_651_503# sky130_fd_sc_hs__dfxtp_4_35/a_696_458#
+ sky130_fd_sc_hs__dfxtp_4_35/a_544_485# sky130_fd_sc_hs__dfxtp_4_35/a_1178_124# sky130_fd_sc_hs__dfxtp_4_35/a_1034_424#
+ sky130_fd_sc_hs__dfxtp_4
Xsky130_fd_sc_hs__dfxtp_4_24 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__a22o_1_5/B2 sky130_fd_sc_hs__dfxtp_4_24/D
+ sky130_fd_sc_hs__clkbuf_4_1/X sky130_fd_sc_hs__dfxtp_4_24/a_1226_296# sky130_fd_sc_hs__dfxtp_4_24/a_735_102#
+ sky130_fd_sc_hs__dfxtp_4_24/a_1141_508# sky130_fd_sc_hs__dfxtp_4_24/a_206_368# sky130_fd_sc_hs__dfxtp_4_24/a_437_503#
+ sky130_fd_sc_hs__dfxtp_4_24/a_27_74# sky130_fd_sc_hs__dfxtp_4_24/a_651_503# sky130_fd_sc_hs__dfxtp_4_24/a_696_458#
+ sky130_fd_sc_hs__dfxtp_4_24/a_544_485# sky130_fd_sc_hs__dfxtp_4_24/a_1178_124# sky130_fd_sc_hs__dfxtp_4_24/a_1034_424#
+ sky130_fd_sc_hs__dfxtp_4
Xsky130_fd_sc_hs__inv_4_1 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_1/Y clk_prbs
+ sky130_fd_sc_hs__inv_4
Xsky130_fd_sc_hs__dfxtp_4_14 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__a22o_1_7/A2 sky130_fd_sc_hs__dfxtp_4_15/D
+ sky130_fd_sc_hs__clkbuf_4_1/X sky130_fd_sc_hs__dfxtp_4_15/a_1226_296# sky130_fd_sc_hs__dfxtp_4_15/a_735_102#
+ sky130_fd_sc_hs__dfxtp_4_15/a_1141_508# sky130_fd_sc_hs__dfxtp_4_15/a_206_368# sky130_fd_sc_hs__dfxtp_4_15/a_437_503#
+ sky130_fd_sc_hs__dfxtp_4_15/a_27_74# sky130_fd_sc_hs__dfxtp_4_15/a_651_503# sky130_fd_sc_hs__dfxtp_4_15/a_696_458#
+ sky130_fd_sc_hs__dfxtp_4_15/a_544_485# sky130_fd_sc_hs__dfxtp_4_15/a_1178_124# sky130_fd_sc_hs__dfxtp_4_15/a_1034_424#
+ sky130_fd_sc_hs__dfxtp_4
Xsky130_fd_sc_hs__dfxtp_4_47 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__dfxtp_4_47/Q sky130_fd_sc_hs__dfxtp_4_47/D
+ sky130_fd_sc_hs__clkbuf_4_1/X sky130_fd_sc_hs__dfxtp_4_47/a_1226_296# sky130_fd_sc_hs__dfxtp_4_47/a_735_102#
+ sky130_fd_sc_hs__dfxtp_4_47/a_1141_508# sky130_fd_sc_hs__dfxtp_4_47/a_206_368# sky130_fd_sc_hs__dfxtp_4_47/a_437_503#
+ sky130_fd_sc_hs__dfxtp_4_47/a_27_74# sky130_fd_sc_hs__dfxtp_4_47/a_651_503# sky130_fd_sc_hs__dfxtp_4_47/a_696_458#
+ sky130_fd_sc_hs__dfxtp_4_47/a_544_485# sky130_fd_sc_hs__dfxtp_4_47/a_1178_124# sky130_fd_sc_hs__dfxtp_4_47/a_1034_424#
+ sky130_fd_sc_hs__dfxtp_4
Xsky130_fd_sc_hs__dfxtp_4_36 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__dfxtp_4_37/Q sky130_fd_sc_hs__a22o_1_19/X
+ sky130_fd_sc_hs__inv_4_19/A sky130_fd_sc_hs__dfxtp_4_37/a_1226_296# sky130_fd_sc_hs__dfxtp_4_37/a_735_102#
+ sky130_fd_sc_hs__dfxtp_4_37/a_1141_508# sky130_fd_sc_hs__dfxtp_4_37/a_206_368# sky130_fd_sc_hs__dfxtp_4_37/a_437_503#
+ sky130_fd_sc_hs__dfxtp_4_37/a_27_74# sky130_fd_sc_hs__dfxtp_4_37/a_651_503# sky130_fd_sc_hs__dfxtp_4_37/a_696_458#
+ sky130_fd_sc_hs__dfxtp_4_37/a_544_485# sky130_fd_sc_hs__dfxtp_4_37/a_1178_124# sky130_fd_sc_hs__dfxtp_4_37/a_1034_424#
+ sky130_fd_sc_hs__dfxtp_4
Xsky130_fd_sc_hs__dfxtp_4_25 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__a22o_1_7/B2 sky130_fd_sc_hs__dfxtp_4_25/D
+ sky130_fd_sc_hs__clkbuf_4_1/X sky130_fd_sc_hs__dfxtp_4_25/a_1226_296# sky130_fd_sc_hs__dfxtp_4_25/a_735_102#
+ sky130_fd_sc_hs__dfxtp_4_25/a_1141_508# sky130_fd_sc_hs__dfxtp_4_25/a_206_368# sky130_fd_sc_hs__dfxtp_4_25/a_437_503#
+ sky130_fd_sc_hs__dfxtp_4_25/a_27_74# sky130_fd_sc_hs__dfxtp_4_25/a_651_503# sky130_fd_sc_hs__dfxtp_4_25/a_696_458#
+ sky130_fd_sc_hs__dfxtp_4_25/a_544_485# sky130_fd_sc_hs__dfxtp_4_25/a_1178_124# sky130_fd_sc_hs__dfxtp_4_25/a_1034_424#
+ sky130_fd_sc_hs__dfxtp_4
Xsky130_fd_sc_hs__clkinv_4_0 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__clkinv_4_1/Y sky130_fd_sc_hs__dfrtp_4_1/Q
+ sky130_fd_sc_hs__clkinv_4
Xsky130_fd_sc_hs__clkbuf_4_0 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_11/A sky130_fd_sc_hs__clkbuf_4_1/X
+ sky130_fd_sc_hs__clkbuf_4_1/a_83_270# sky130_fd_sc_hs__clkbuf_4
Xsky130_fd_sc_hs__inv_4_2 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_3/Y clk_prbs
+ sky130_fd_sc_hs__inv_4
Xsky130_fd_sc_hs__clkbuf_2_30 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__dfxtp_4_47/D din[2]
+ sky130_fd_sc_hs__clkbuf_2_31/a_43_192# sky130_fd_sc_hs__clkbuf_2
Xsky130_fd_sc_hs__dfxtp_4_15 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__a22o_1_7/A2 sky130_fd_sc_hs__dfxtp_4_15/D
+ sky130_fd_sc_hs__clkbuf_4_1/X sky130_fd_sc_hs__dfxtp_4_15/a_1226_296# sky130_fd_sc_hs__dfxtp_4_15/a_735_102#
+ sky130_fd_sc_hs__dfxtp_4_15/a_1141_508# sky130_fd_sc_hs__dfxtp_4_15/a_206_368# sky130_fd_sc_hs__dfxtp_4_15/a_437_503#
+ sky130_fd_sc_hs__dfxtp_4_15/a_27_74# sky130_fd_sc_hs__dfxtp_4_15/a_651_503# sky130_fd_sc_hs__dfxtp_4_15/a_696_458#
+ sky130_fd_sc_hs__dfxtp_4_15/a_544_485# sky130_fd_sc_hs__dfxtp_4_15/a_1178_124# sky130_fd_sc_hs__dfxtp_4_15/a_1034_424#
+ sky130_fd_sc_hs__dfxtp_4
Xsky130_fd_sc_hs__dfxtp_4_37 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__dfxtp_4_37/Q sky130_fd_sc_hs__a22o_1_19/X
+ sky130_fd_sc_hs__inv_4_19/A sky130_fd_sc_hs__dfxtp_4_37/a_1226_296# sky130_fd_sc_hs__dfxtp_4_37/a_735_102#
+ sky130_fd_sc_hs__dfxtp_4_37/a_1141_508# sky130_fd_sc_hs__dfxtp_4_37/a_206_368# sky130_fd_sc_hs__dfxtp_4_37/a_437_503#
+ sky130_fd_sc_hs__dfxtp_4_37/a_27_74# sky130_fd_sc_hs__dfxtp_4_37/a_651_503# sky130_fd_sc_hs__dfxtp_4_37/a_696_458#
+ sky130_fd_sc_hs__dfxtp_4_37/a_544_485# sky130_fd_sc_hs__dfxtp_4_37/a_1178_124# sky130_fd_sc_hs__dfxtp_4_37/a_1034_424#
+ sky130_fd_sc_hs__dfxtp_4
Xsky130_fd_sc_hs__dfxtp_4_26 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__dfxtp_4_27/Q sky130_fd_sc_hs__dfxtp_4_27/D
+ sky130_fd_sc_hs__clkbuf_4_1/X sky130_fd_sc_hs__dfxtp_4_27/a_1226_296# sky130_fd_sc_hs__dfxtp_4_27/a_735_102#
+ sky130_fd_sc_hs__dfxtp_4_27/a_1141_508# sky130_fd_sc_hs__dfxtp_4_27/a_206_368# sky130_fd_sc_hs__dfxtp_4_27/a_437_503#
+ sky130_fd_sc_hs__dfxtp_4_27/a_27_74# sky130_fd_sc_hs__dfxtp_4_27/a_651_503# sky130_fd_sc_hs__dfxtp_4_27/a_696_458#
+ sky130_fd_sc_hs__dfxtp_4_27/a_544_485# sky130_fd_sc_hs__dfxtp_4_27/a_1178_124# sky130_fd_sc_hs__dfxtp_4_27/a_1034_424#
+ sky130_fd_sc_hs__dfxtp_4
Xsky130_fd_sc_hs__clkinv_4_1 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__clkinv_4_1/Y sky130_fd_sc_hs__dfrtp_4_1/Q
+ sky130_fd_sc_hs__clkinv_4
Xsky130_fd_sc_hs__clkbuf_4_1 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_11/A sky130_fd_sc_hs__clkbuf_4_1/X
+ sky130_fd_sc_hs__clkbuf_4_1/a_83_270# sky130_fd_sc_hs__clkbuf_4
Xsky130_fd_sc_hs__inv_4_3 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_3/Y clk_prbs
+ sky130_fd_sc_hs__inv_4
Xsky130_fd_sc_hs__clkbuf_2_31 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__dfxtp_4_47/D din[2]
+ sky130_fd_sc_hs__clkbuf_2_31/a_43_192# sky130_fd_sc_hs__clkbuf_2
Xsky130_fd_sc_hs__a22o_1_20 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__a22o_1_21/X sky130_fd_sc_hs__dfxtp_4_47/Q
+ sky130_fd_sc_hs__inv_4_17/Y sky130_fd_sc_hs__dfxtp_4_39/Q sky130_fd_sc_hs__buf_2_15/X
+ sky130_fd_sc_hs__a22o_1_21/a_222_392# sky130_fd_sc_hs__a22o_1_21/a_230_79# sky130_fd_sc_hs__a22o_1_21/a_52_123#
+ sky130_fd_sc_hs__a22o_1_21/a_132_392# sky130_fd_sc_hs__a22o_1
Xsky130_fd_sc_hs__clkbuf_2_20 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__dfxtp_4_31/D din[5]
+ sky130_fd_sc_hs__clkbuf_2_21/a_43_192# sky130_fd_sc_hs__clkbuf_2
Xsky130_fd_sc_hs__buf_2_0 DVSS DVDD DVDD DVSS clk_prbs sky130_fd_sc_hs__buf_2_1/X
+ sky130_fd_sc_hs__buf_2_1/a_21_260# sky130_fd_sc_hs__buf_2
Xsky130_fd_sc_hs__dfxtp_4_38 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__dfxtp_4_39/Q sky130_fd_sc_hs__dfxtp_4_39/D
+ sky130_fd_sc_hs__clkbuf_4_1/X sky130_fd_sc_hs__dfxtp_4_39/a_1226_296# sky130_fd_sc_hs__dfxtp_4_39/a_735_102#
+ sky130_fd_sc_hs__dfxtp_4_39/a_1141_508# sky130_fd_sc_hs__dfxtp_4_39/a_206_368# sky130_fd_sc_hs__dfxtp_4_39/a_437_503#
+ sky130_fd_sc_hs__dfxtp_4_39/a_27_74# sky130_fd_sc_hs__dfxtp_4_39/a_651_503# sky130_fd_sc_hs__dfxtp_4_39/a_696_458#
+ sky130_fd_sc_hs__dfxtp_4_39/a_544_485# sky130_fd_sc_hs__dfxtp_4_39/a_1178_124# sky130_fd_sc_hs__dfxtp_4_39/a_1034_424#
+ sky130_fd_sc_hs__dfxtp_4
Xsky130_fd_sc_hs__dfxtp_4_27 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__dfxtp_4_27/Q sky130_fd_sc_hs__dfxtp_4_27/D
+ sky130_fd_sc_hs__clkbuf_4_1/X sky130_fd_sc_hs__dfxtp_4_27/a_1226_296# sky130_fd_sc_hs__dfxtp_4_27/a_735_102#
+ sky130_fd_sc_hs__dfxtp_4_27/a_1141_508# sky130_fd_sc_hs__dfxtp_4_27/a_206_368# sky130_fd_sc_hs__dfxtp_4_27/a_437_503#
+ sky130_fd_sc_hs__dfxtp_4_27/a_27_74# sky130_fd_sc_hs__dfxtp_4_27/a_651_503# sky130_fd_sc_hs__dfxtp_4_27/a_696_458#
+ sky130_fd_sc_hs__dfxtp_4_27/a_544_485# sky130_fd_sc_hs__dfxtp_4_27/a_1178_124# sky130_fd_sc_hs__dfxtp_4_27/a_1034_424#
+ sky130_fd_sc_hs__dfxtp_4
Xsky130_fd_sc_hs__dfxtp_4_16 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__dfxtp_4_18/Q sky130_fd_sc_hs__a22o_1_5/X
+ sky130_fd_sc_hs__inv_4_19/A sky130_fd_sc_hs__dfxtp_4_18/a_1226_296# sky130_fd_sc_hs__dfxtp_4_18/a_735_102#
+ sky130_fd_sc_hs__dfxtp_4_18/a_1141_508# sky130_fd_sc_hs__dfxtp_4_18/a_206_368# sky130_fd_sc_hs__dfxtp_4_18/a_437_503#
+ sky130_fd_sc_hs__dfxtp_4_18/a_27_74# sky130_fd_sc_hs__dfxtp_4_18/a_651_503# sky130_fd_sc_hs__dfxtp_4_18/a_696_458#
+ sky130_fd_sc_hs__dfxtp_4_18/a_544_485# sky130_fd_sc_hs__dfxtp_4_18/a_1178_124# sky130_fd_sc_hs__dfxtp_4_18/a_1034_424#
+ sky130_fd_sc_hs__dfxtp_4
Xsky130_fd_sc_hs__clkbuf_4_2 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__dfrtp_4_1/Q sky130_fd_sc_hs__inv_4_19/A
+ sky130_fd_sc_hs__clkbuf_4_3/a_83_270# sky130_fd_sc_hs__clkbuf_4
Xsky130_fd_sc_hs__inv_4_4 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_5/Y clk_prbs
+ sky130_fd_sc_hs__inv_4
Xsky130_fd_sc_hs__clkbuf_2_10 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__dfxtp_4_8/D din[11]
+ sky130_fd_sc_hs__clkbuf_2_11/a_43_192# sky130_fd_sc_hs__clkbuf_2
Xsky130_fd_sc_hs__a22o_1_21 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__a22o_1_21/X sky130_fd_sc_hs__dfxtp_4_47/Q
+ sky130_fd_sc_hs__inv_4_17/Y sky130_fd_sc_hs__dfxtp_4_39/Q sky130_fd_sc_hs__buf_2_15/X
+ sky130_fd_sc_hs__a22o_1_21/a_222_392# sky130_fd_sc_hs__a22o_1_21/a_230_79# sky130_fd_sc_hs__a22o_1_21/a_52_123#
+ sky130_fd_sc_hs__a22o_1_21/a_132_392# sky130_fd_sc_hs__a22o_1
Xsky130_fd_sc_hs__clkbuf_2_21 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__dfxtp_4_31/D din[5]
+ sky130_fd_sc_hs__clkbuf_2_21/a_43_192# sky130_fd_sc_hs__clkbuf_2
Xsky130_fd_sc_hs__a22o_1_10 DVSS DVDD DVDD DVSS dout[0] sky130_fd_sc_hs__dfxtp_4_41/Q
+ sky130_fd_sc_hs__a22o_1_9/B1 sky130_fd_sc_hs__dfxtp_4_33/Q sky130_fd_sc_hs__inv_4_19/A
+ sky130_fd_sc_hs__a22o_1_11/a_222_392# sky130_fd_sc_hs__a22o_1_11/a_230_79# sky130_fd_sc_hs__a22o_1_11/a_52_123#
+ sky130_fd_sc_hs__a22o_1_11/a_132_392# sky130_fd_sc_hs__a22o_1
Xsky130_fd_sc_hs__buf_2_1 DVSS DVDD DVDD DVSS clk_prbs sky130_fd_sc_hs__buf_2_1/X
+ sky130_fd_sc_hs__buf_2_1/a_21_260# sky130_fd_sc_hs__buf_2
Xsky130_fd_sc_hs__dfxtp_4_0 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__dfxtp_4_1/Q sky130_fd_sc_hs__dfxtp_4_1/D
+ sky130_fd_sc_hs__clkbuf_4_1/X sky130_fd_sc_hs__dfxtp_4_1/a_1226_296# sky130_fd_sc_hs__dfxtp_4_1/a_735_102#
+ sky130_fd_sc_hs__dfxtp_4_1/a_1141_508# sky130_fd_sc_hs__dfxtp_4_1/a_206_368# sky130_fd_sc_hs__dfxtp_4_1/a_437_503#
+ sky130_fd_sc_hs__dfxtp_4_1/a_27_74# sky130_fd_sc_hs__dfxtp_4_1/a_651_503# sky130_fd_sc_hs__dfxtp_4_1/a_696_458#
+ sky130_fd_sc_hs__dfxtp_4_1/a_544_485# sky130_fd_sc_hs__dfxtp_4_1/a_1178_124# sky130_fd_sc_hs__dfxtp_4_1/a_1034_424#
+ sky130_fd_sc_hs__dfxtp_4
Xsky130_fd_sc_hs__dfxtp_4_28 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__dfxtp_4_29/Q sky130_fd_sc_hs__a22o_1_17/X
+ sky130_fd_sc_hs__inv_4_19/A sky130_fd_sc_hs__dfxtp_4_29/a_1226_296# sky130_fd_sc_hs__dfxtp_4_29/a_735_102#
+ sky130_fd_sc_hs__dfxtp_4_29/a_1141_508# sky130_fd_sc_hs__dfxtp_4_29/a_206_368# sky130_fd_sc_hs__dfxtp_4_29/a_437_503#
+ sky130_fd_sc_hs__dfxtp_4_29/a_27_74# sky130_fd_sc_hs__dfxtp_4_29/a_651_503# sky130_fd_sc_hs__dfxtp_4_29/a_696_458#
+ sky130_fd_sc_hs__dfxtp_4_29/a_544_485# sky130_fd_sc_hs__dfxtp_4_29/a_1178_124# sky130_fd_sc_hs__dfxtp_4_29/a_1034_424#
+ sky130_fd_sc_hs__dfxtp_4
Xsky130_fd_sc_hs__dfxtp_4_17 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__dfxtp_4_19/Q sky130_fd_sc_hs__a22o_1_7/X
+ sky130_fd_sc_hs__inv_4_19/A sky130_fd_sc_hs__dfxtp_4_19/a_1226_296# sky130_fd_sc_hs__dfxtp_4_19/a_735_102#
+ sky130_fd_sc_hs__dfxtp_4_19/a_1141_508# sky130_fd_sc_hs__dfxtp_4_19/a_206_368# sky130_fd_sc_hs__dfxtp_4_19/a_437_503#
+ sky130_fd_sc_hs__dfxtp_4_19/a_27_74# sky130_fd_sc_hs__dfxtp_4_19/a_651_503# sky130_fd_sc_hs__dfxtp_4_19/a_696_458#
+ sky130_fd_sc_hs__dfxtp_4_19/a_544_485# sky130_fd_sc_hs__dfxtp_4_19/a_1178_124# sky130_fd_sc_hs__dfxtp_4_19/a_1034_424#
+ sky130_fd_sc_hs__dfxtp_4
Xsky130_fd_sc_hs__dfxtp_4_39 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__dfxtp_4_39/Q sky130_fd_sc_hs__dfxtp_4_39/D
+ sky130_fd_sc_hs__clkbuf_4_1/X sky130_fd_sc_hs__dfxtp_4_39/a_1226_296# sky130_fd_sc_hs__dfxtp_4_39/a_735_102#
+ sky130_fd_sc_hs__dfxtp_4_39/a_1141_508# sky130_fd_sc_hs__dfxtp_4_39/a_206_368# sky130_fd_sc_hs__dfxtp_4_39/a_437_503#
+ sky130_fd_sc_hs__dfxtp_4_39/a_27_74# sky130_fd_sc_hs__dfxtp_4_39/a_651_503# sky130_fd_sc_hs__dfxtp_4_39/a_696_458#
+ sky130_fd_sc_hs__dfxtp_4_39/a_544_485# sky130_fd_sc_hs__dfxtp_4_39/a_1178_124# sky130_fd_sc_hs__dfxtp_4_39/a_1034_424#
+ sky130_fd_sc_hs__dfxtp_4
Xsky130_fd_sc_hs__clkbuf_4_3 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__dfrtp_4_1/Q sky130_fd_sc_hs__inv_4_19/A
+ sky130_fd_sc_hs__clkbuf_4_3/a_83_270# sky130_fd_sc_hs__clkbuf_4
Xsky130_fd_sc_hs__inv_4_5 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_5/Y clk_prbs
+ sky130_fd_sc_hs__inv_4
Xsky130_fd_sc_hs__clkbuf_2_0 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__dfxtp_4_1/D din[14]
+ sky130_fd_sc_hs__clkbuf_2_1/a_43_192# sky130_fd_sc_hs__clkbuf_2
Xsky130_fd_sc_hs__clkbuf_2_11 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__dfxtp_4_8/D din[11]
+ sky130_fd_sc_hs__clkbuf_2_11/a_43_192# sky130_fd_sc_hs__clkbuf_2
Xsky130_fd_sc_hs__a22o_1_22 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__a22o_1_23/X sky130_fd_sc_hs__dfxtp_4_46/Q
+ sky130_fd_sc_hs__inv_4_21/Y sky130_fd_sc_hs__dfxtp_4_45/Q sky130_fd_sc_hs__buf_2_14/X
+ sky130_fd_sc_hs__a22o_1_23/a_222_392# sky130_fd_sc_hs__a22o_1_23/a_230_79# sky130_fd_sc_hs__a22o_1_23/a_52_123#
+ sky130_fd_sc_hs__a22o_1_23/a_132_392# sky130_fd_sc_hs__a22o_1
Xsky130_fd_sc_hs__clkbuf_2_22 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__dfxtp_4_39/D din[3]
+ sky130_fd_sc_hs__clkbuf_2_23/a_43_192# sky130_fd_sc_hs__clkbuf_2
Xsky130_fd_sc_hs__a22o_1_11 DVSS DVDD DVDD DVSS dout[0] sky130_fd_sc_hs__dfxtp_4_41/Q
+ sky130_fd_sc_hs__a22o_1_9/B1 sky130_fd_sc_hs__dfxtp_4_33/Q sky130_fd_sc_hs__inv_4_19/A
+ sky130_fd_sc_hs__a22o_1_11/a_222_392# sky130_fd_sc_hs__a22o_1_11/a_230_79# sky130_fd_sc_hs__a22o_1_11/a_52_123#
+ sky130_fd_sc_hs__a22o_1_11/a_132_392# sky130_fd_sc_hs__a22o_1
Xsky130_fd_sc_hs__clkinv_2_0 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__clkinv_2_1/Y rst
+ sky130_fd_sc_hs__clkinv_2
Xsky130_fd_sc_hs__buf_2_2 DVSS DVDD DVDD DVSS clk_prbs sky130_fd_sc_hs__buf_2_3/X
+ sky130_fd_sc_hs__buf_2_3/a_21_260# sky130_fd_sc_hs__buf_2
Xsky130_fd_sc_hs__dfxtp_4_1 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__dfxtp_4_1/Q sky130_fd_sc_hs__dfxtp_4_1/D
+ sky130_fd_sc_hs__clkbuf_4_1/X sky130_fd_sc_hs__dfxtp_4_1/a_1226_296# sky130_fd_sc_hs__dfxtp_4_1/a_735_102#
+ sky130_fd_sc_hs__dfxtp_4_1/a_1141_508# sky130_fd_sc_hs__dfxtp_4_1/a_206_368# sky130_fd_sc_hs__dfxtp_4_1/a_437_503#
+ sky130_fd_sc_hs__dfxtp_4_1/a_27_74# sky130_fd_sc_hs__dfxtp_4_1/a_651_503# sky130_fd_sc_hs__dfxtp_4_1/a_696_458#
+ sky130_fd_sc_hs__dfxtp_4_1/a_544_485# sky130_fd_sc_hs__dfxtp_4_1/a_1178_124# sky130_fd_sc_hs__dfxtp_4_1/a_1034_424#
+ sky130_fd_sc_hs__dfxtp_4
Xsky130_fd_sc_hs__dfxtp_4_29 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__dfxtp_4_29/Q sky130_fd_sc_hs__a22o_1_17/X
+ sky130_fd_sc_hs__inv_4_19/A sky130_fd_sc_hs__dfxtp_4_29/a_1226_296# sky130_fd_sc_hs__dfxtp_4_29/a_735_102#
+ sky130_fd_sc_hs__dfxtp_4_29/a_1141_508# sky130_fd_sc_hs__dfxtp_4_29/a_206_368# sky130_fd_sc_hs__dfxtp_4_29/a_437_503#
+ sky130_fd_sc_hs__dfxtp_4_29/a_27_74# sky130_fd_sc_hs__dfxtp_4_29/a_651_503# sky130_fd_sc_hs__dfxtp_4_29/a_696_458#
+ sky130_fd_sc_hs__dfxtp_4_29/a_544_485# sky130_fd_sc_hs__dfxtp_4_29/a_1178_124# sky130_fd_sc_hs__dfxtp_4_29/a_1034_424#
+ sky130_fd_sc_hs__dfxtp_4
Xsky130_fd_sc_hs__dfxtp_4_18 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__dfxtp_4_18/Q sky130_fd_sc_hs__a22o_1_5/X
+ sky130_fd_sc_hs__inv_4_19/A sky130_fd_sc_hs__dfxtp_4_18/a_1226_296# sky130_fd_sc_hs__dfxtp_4_18/a_735_102#
+ sky130_fd_sc_hs__dfxtp_4_18/a_1141_508# sky130_fd_sc_hs__dfxtp_4_18/a_206_368# sky130_fd_sc_hs__dfxtp_4_18/a_437_503#
+ sky130_fd_sc_hs__dfxtp_4_18/a_27_74# sky130_fd_sc_hs__dfxtp_4_18/a_651_503# sky130_fd_sc_hs__dfxtp_4_18/a_696_458#
+ sky130_fd_sc_hs__dfxtp_4_18/a_544_485# sky130_fd_sc_hs__dfxtp_4_18/a_1178_124# sky130_fd_sc_hs__dfxtp_4_18/a_1034_424#
+ sky130_fd_sc_hs__dfxtp_4
Xsky130_fd_sc_hs__inv_4_6 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_7/Y rst sky130_fd_sc_hs__inv_4
Xsky130_fd_sc_hs__clkbuf_2_1 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__dfxtp_4_1/D din[14]
+ sky130_fd_sc_hs__clkbuf_2_1/a_43_192# sky130_fd_sc_hs__clkbuf_2
Xsky130_fd_sc_hs__clkbuf_2_12 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__dfxtp_4_24/D din[10]
+ sky130_fd_sc_hs__clkbuf_2_13/a_43_192# sky130_fd_sc_hs__clkbuf_2
Xsky130_fd_sc_hs__a22o_1_23 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__a22o_1_23/X sky130_fd_sc_hs__dfxtp_4_46/Q
+ sky130_fd_sc_hs__inv_4_21/Y sky130_fd_sc_hs__dfxtp_4_45/Q sky130_fd_sc_hs__buf_2_14/X
+ sky130_fd_sc_hs__a22o_1_23/a_222_392# sky130_fd_sc_hs__a22o_1_23/a_230_79# sky130_fd_sc_hs__a22o_1_23/a_52_123#
+ sky130_fd_sc_hs__a22o_1_23/a_132_392# sky130_fd_sc_hs__a22o_1
Xsky130_fd_sc_hs__clkbuf_2_23 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__dfxtp_4_39/D din[3]
+ sky130_fd_sc_hs__clkbuf_2_23/a_43_192# sky130_fd_sc_hs__clkbuf_2
Xsky130_fd_sc_hs__a22o_1_12 DVSS DVDD DVDD DVSS dout[2] sky130_fd_sc_hs__dfxtp_4_19/Q
+ sky130_fd_sc_hs__a22o_1_9/B1 sky130_fd_sc_hs__dfxtp_4_18/Q sky130_fd_sc_hs__inv_4_19/A
+ sky130_fd_sc_hs__a22o_1_14/a_222_392# sky130_fd_sc_hs__a22o_1_14/a_230_79# sky130_fd_sc_hs__a22o_1_14/a_52_123#
+ sky130_fd_sc_hs__a22o_1_14/a_132_392# sky130_fd_sc_hs__a22o_1
Xsky130_fd_sc_hs__buf_2_3 DVSS DVDD DVDD DVSS clk_prbs sky130_fd_sc_hs__buf_2_3/X
+ sky130_fd_sc_hs__buf_2_3/a_21_260# sky130_fd_sc_hs__buf_2
Xsky130_fd_sc_hs__clkinv_2_1 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__clkinv_2_1/Y rst
+ sky130_fd_sc_hs__clkinv_2
Xsky130_fd_sc_hs__dfxtp_4_2 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__dfxtp_4_3/Q sky130_fd_sc_hs__dfxtp_4_3/D
+ sky130_fd_sc_hs__clkbuf_4_1/X sky130_fd_sc_hs__dfxtp_4_3/a_1226_296# sky130_fd_sc_hs__dfxtp_4_3/a_735_102#
+ sky130_fd_sc_hs__dfxtp_4_3/a_1141_508# sky130_fd_sc_hs__dfxtp_4_3/a_206_368# sky130_fd_sc_hs__dfxtp_4_3/a_437_503#
+ sky130_fd_sc_hs__dfxtp_4_3/a_27_74# sky130_fd_sc_hs__dfxtp_4_3/a_651_503# sky130_fd_sc_hs__dfxtp_4_3/a_696_458#
+ sky130_fd_sc_hs__dfxtp_4_3/a_544_485# sky130_fd_sc_hs__dfxtp_4_3/a_1178_124# sky130_fd_sc_hs__dfxtp_4_3/a_1034_424#
+ sky130_fd_sc_hs__dfxtp_4
Xsky130_fd_sc_hs__dfxtp_4_19 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__dfxtp_4_19/Q sky130_fd_sc_hs__a22o_1_7/X
+ sky130_fd_sc_hs__inv_4_19/A sky130_fd_sc_hs__dfxtp_4_19/a_1226_296# sky130_fd_sc_hs__dfxtp_4_19/a_735_102#
+ sky130_fd_sc_hs__dfxtp_4_19/a_1141_508# sky130_fd_sc_hs__dfxtp_4_19/a_206_368# sky130_fd_sc_hs__dfxtp_4_19/a_437_503#
+ sky130_fd_sc_hs__dfxtp_4_19/a_27_74# sky130_fd_sc_hs__dfxtp_4_19/a_651_503# sky130_fd_sc_hs__dfxtp_4_19/a_696_458#
+ sky130_fd_sc_hs__dfxtp_4_19/a_544_485# sky130_fd_sc_hs__dfxtp_4_19/a_1178_124# sky130_fd_sc_hs__dfxtp_4_19/a_1034_424#
+ sky130_fd_sc_hs__dfxtp_4
Xsky130_fd_sc_hs__clkbuf_2_2 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__dfxtp_4_3/D din[15]
+ sky130_fd_sc_hs__clkbuf_2_3/a_43_192# sky130_fd_sc_hs__clkbuf_2
Xsky130_fd_sc_hs__clkbuf_2_13 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__dfxtp_4_24/D din[10]
+ sky130_fd_sc_hs__clkbuf_2_13/a_43_192# sky130_fd_sc_hs__clkbuf_2
Xsky130_fd_sc_hs__clkbuf_2_24 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__dfxtp_4_35/D din[4]
+ sky130_fd_sc_hs__clkbuf_2_25/a_43_192# sky130_fd_sc_hs__clkbuf_2
Xsky130_fd_sc_hs__a22o_1_13 DVSS DVDD DVDD DVSS dout[1] sky130_fd_sc_hs__dfxtp_4_37/Q
+ sky130_fd_sc_hs__a22o_1_9/B1 sky130_fd_sc_hs__dfxtp_4_29/Q sky130_fd_sc_hs__inv_4_19/A
+ sky130_fd_sc_hs__a22o_1_15/a_222_392# sky130_fd_sc_hs__a22o_1_15/a_230_79# sky130_fd_sc_hs__a22o_1_15/a_52_123#
+ sky130_fd_sc_hs__a22o_1_15/a_132_392# sky130_fd_sc_hs__a22o_1
Xsky130_fd_sc_hs__inv_4_7 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__inv_4_7/Y rst sky130_fd_sc_hs__inv_4
Xsky130_fd_sc_hs__dfxtp_4_3 DVSS DVDD DVDD DVSS sky130_fd_sc_hs__dfxtp_4_3/Q sky130_fd_sc_hs__dfxtp_4_3/D
+ sky130_fd_sc_hs__clkbuf_4_1/X sky130_fd_sc_hs__dfxtp_4_3/a_1226_296# sky130_fd_sc_hs__dfxtp_4_3/a_735_102#
+ sky130_fd_sc_hs__dfxtp_4_3/a_1141_508# sky130_fd_sc_hs__dfxtp_4_3/a_206_368# sky130_fd_sc_hs__dfxtp_4_3/a_437_503#
+ sky130_fd_sc_hs__dfxtp_4_3/a_27_74# sky130_fd_sc_hs__dfxtp_4_3/a_651_503# sky130_fd_sc_hs__dfxtp_4_3/a_696_458#
+ sky130_fd_sc_hs__dfxtp_4_3/a_544_485# sky130_fd_sc_hs__dfxtp_4_3/a_1178_124# sky130_fd_sc_hs__dfxtp_4_3/a_1034_424#
+ sky130_fd_sc_hs__dfxtp_4
Xsky130_fd_sc_hs__buf_2_4 DVSS DVDD DVDD DVSS clk_prbs sky130_fd_sc_hs__buf_2_5/X
+ sky130_fd_sc_hs__buf_2_5/a_21_260# sky130_fd_sc_hs__buf_2
.ends

.subckt sky130_fd_sc_hs__and2_4 VNB VPB VPWR VGND X A B a_83_269# a_504_119#
X0 a_83_269# A a_504_119# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X1 VPWR a_83_269# X VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X2 VGND a_83_269# X VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X3 X a_83_269# VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X4 X a_83_269# VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X5 VPWR a_83_269# X VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X6 VPWR B a_83_269# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X7 a_83_269# A VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X8 VGND a_83_269# X VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X9 VPWR A a_83_269# VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X10 VGND B a_504_119# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X11 a_504_119# A a_83_269# VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X12 X a_83_269# VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X13 a_504_119# B VGND VNB sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X14 X a_83_269# VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X15 a_83_269# B VPWR VPB sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
.ends

.subckt digital_top rst rst_prbs inj_error ref_clk_ext_p ref_clk_ext_n CTL_BUF_N[5]
+ CTL_BUF_N[4] CTL_BUF_N[3] CTL_BUF_N[2] CTL_BUF_N[1] CTL_BUF_N[0] CTL_BUF_P[5] CTL_BUF_P[4]
+ CTL_BUF_P[3] CTL_BUF_P[2] CTL_BUF_P[1] CTL_BUF_P[0] osc_en aux_osc_en inj_en fftl_en
+ con_perb[3] con_perb[2] con_perb[1] con_perb[0] div_ratio_half[5] div_ratio_half[4]
+ div_ratio_half[3] div_ratio_half[2] div_ratio_half[1] div_ratio_half[0] fine_control_avg_window_select[4]
+ fine_control_avg_window_select[3] fine_control_avg_window_select[2] fine_control_avg_window_select[1]
+ fine_control_avg_window_select[0] fine_con_step_size[3] fine_con_step_size[2] fine_con_step_size[1]
+ fine_con_step_size[0] manual_control_osc[12] manual_control_osc[11] manual_control_osc[10]
+ manual_control_osc[9] manual_control_osc[8] manual_control_osc[7] manual_control_osc[6]
+ manual_control_osc[5] manual_control_osc[4] manual_control_osc[3] manual_control_osc[2]
+ manual_control_osc[1] manual_control_osc[0] pi1_con[3] pi1_con[2] pi1_con[1] pi1_con[0]
+ pi2_con[3] pi2_con[2] pi2_con[1] pi2_con[0] pi3_con[3] pi3_con[2] pi3_con[1] pi3_con[0]
+ pi4_con[3] pi4_con[2] pi4_con[1] pi4_con[0] pi5_con[3] pi5_con[2] pi5_con[1] pi5_con[0]
+ test_mux_select[3] test_mux_select[2] test_mux_select[1] test_mux_select[0] test_mux_clk_I_select[1]
+ test_mux_clk_I_select[0] test_mux_clk_Q_select[1] test_mux_clk_Q_select[0] dout_p
+ dout_n test_mux_misc test_mux_clk_Q test_mux_clk_I DVSS: DVDD: AVDD
Xsky130_fd_sc_hs__or2b_4_1 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__or2b_4_1/A sky130_fd_sc_hs__nor4_2_1/A
+ sky130_fd_sc_hs__or2b_4_1/X sky130_fd_sc_hs__or2b_4_1/a_676_48# sky130_fd_sc_hs__or2b_4_1/a_489_392#
+ sky130_fd_sc_hs__or2b_4_1/a_81_296# sky130_fd_sc_hs__or2b_4
Xsky130_fd_sc_hs__buf_2_160 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__buf_2_161/A sky130_fd_sc_hs__buf_2_161/X
+ sky130_fd_sc_hs__buf_2_161/a_21_260# sky130_fd_sc_hs__buf_2
Xsky130_fd_sc_hs__clkbuf_4_6 DVSS: DVDD: DVDD: DVSS: pi2_con[0] sky130_fd_sc_hs__clkbuf_4_7/X
+ sky130_fd_sc_hs__clkbuf_4_7/a_83_270# sky130_fd_sc_hs__clkbuf_4
Xsky130_fd_sc_hs__einvp_2_50 DVSS: DVDD: DVDD: DVSS: dout_n sky130_fd_sc_hs__buf_8_1/X
+ sky130_fd_sc_hs__dlrtp_1_37/Q sky130_fd_sc_hs__einvp_2_51/a_263_323# sky130_fd_sc_hs__einvp_2_51/a_36_74#
+ sky130_fd_sc_hs__einvp_2_51/a_27_368# sky130_fd_sc_hs__einvp_2
Xsky130_fd_sc_hs__einvp_2_61 DVSS: DVDD: DVDD: DVSS: dout_p sky130_fd_sc_hs__einvp_2_97/A
+ sky130_fd_sc_hs__dlrtp_1_51/Q sky130_fd_sc_hs__einvp_2_61/a_263_323# sky130_fd_sc_hs__einvp_2_61/a_36_74#
+ sky130_fd_sc_hs__einvp_2_61/a_27_368# sky130_fd_sc_hs__einvp_2
Xsky130_fd_sc_hs__einvp_2_72 DVSS: DVDD: DVDD: DVSS: dout_p sky130_fd_sc_hs__einvp_2_97/A
+ sky130_fd_sc_hs__buf_2_35/X sky130_fd_sc_hs__einvp_2_73/a_263_323# sky130_fd_sc_hs__einvp_2_73/a_36_74#
+ sky130_fd_sc_hs__einvp_2_73/a_27_368# sky130_fd_sc_hs__einvp_2
Xsky130_fd_sc_hs__einvp_2_83 DVSS: DVDD: DVDD: DVSS: dout_p sky130_fd_sc_hs__einvp_2_99/A
+ sky130_fd_sc_hs__buf_2_31/X sky130_fd_sc_hs__einvp_2_83/a_263_323# sky130_fd_sc_hs__einvp_2_83/a_36_74#
+ sky130_fd_sc_hs__einvp_2_83/a_27_368# sky130_fd_sc_hs__einvp_2
Xsky130_fd_sc_hs__einvp_2_94 DVSS: DVDD: DVDD: DVSS: dout_p sky130_fd_sc_hs__einvp_2_97/A
+ sky130_fd_sc_hs__buf_2_71/X sky130_fd_sc_hs__einvp_2_95/a_263_323# sky130_fd_sc_hs__einvp_2_95/a_36_74#
+ sky130_fd_sc_hs__einvp_2_95/a_27_368# sky130_fd_sc_hs__einvp_2
Xsky130_fd_sc_hs__clkinv_4_6 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__clkinv_4_7/Y
+ sky130_fd_sc_hs__nor4_2_1/B sky130_fd_sc_hs__clkinv_4
Xsky130_fd_sc_hs__and2_2_0 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__and2_2_1/A sky130_fd_sc_hs__and2_2_1/B
+ sky130_fd_sc_hs__inv_4_9/A sky130_fd_sc_hs__and2_2_1/a_31_74# sky130_fd_sc_hs__and2_2_1/a_118_74#
+ sky130_fd_sc_hs__and2_2
Xsky130_fd_sc_hs__conb_1_60 DVSS: DVDD: DVDD: DVSS: prbs_generator_syn_7/eqn[8] prbs_generator_syn_7/eqn[1]
+ sky130_fd_sc_hs__conb_1_61/a_165_290# sky130_fd_sc_hs__conb_1_61/a_21_290# sky130_fd_sc_hs__conb_1
Xsky130_fd_sc_hs__conb_1_71 DVSS: DVDD: DVDD: DVSS: prbs_generator_syn_7/eqn[31] prbs_generator_syn_7/cke
+ sky130_fd_sc_hs__conb_1_71/a_165_290# sky130_fd_sc_hs__conb_1_71/a_21_290# sky130_fd_sc_hs__conb_1
Xsky130_fd_sc_hs__conb_1_82 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__conb_1_83/LO
+ sky130_fd_sc_hs__conb_1_83/HI sky130_fd_sc_hs__conb_1_83/a_165_290# sky130_fd_sc_hs__conb_1_83/a_21_290#
+ sky130_fd_sc_hs__conb_1
Xsky130_fd_sc_hs__conb_1_93 DVSS: DVDD: DVDD: DVSS: qr_4t1_mux_top_1/din_3_dummy sky130_fd_sc_hs__conb_1_93/HI
+ sky130_fd_sc_hs__conb_1_93/a_165_290# sky130_fd_sc_hs__conb_1_93/a_21_290# sky130_fd_sc_hs__conb_1
Xsky130_fd_sc_hs__dlrtp_1_105 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__dlrtp_1_105/Q
+ sky130_fd_sc_hs__dlrtp_1_9/GATE sky130_fd_sc_hs__conb_1_133/HI sky130_fd_sc_hs__o21bai_2_31/Y
+ sky130_fd_sc_hs__dlrtp_1_105/a_216_424# sky130_fd_sc_hs__dlrtp_1_105/a_759_508#
+ sky130_fd_sc_hs__dlrtp_1_105/a_565_74# sky130_fd_sc_hs__dlrtp_1_105/a_27_424# sky130_fd_sc_hs__dlrtp_1_105/a_1045_74#
+ sky130_fd_sc_hs__dlrtp_1_105/a_643_74# sky130_fd_sc_hs__dlrtp_1_105/a_817_48# sky130_fd_sc_hs__dlrtp_1_105/a_568_392#
+ sky130_fd_sc_hs__dlrtp_1_105/a_363_74# sky130_fd_sc_hs__dlrtp_1_105/a_769_74# sky130_fd_sc_hs__dlrtp_1
Xsky130_fd_sc_hs__dlrtp_1_116 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__buf_2_119/A
+ sky130_fd_sc_hs__dlrtp_1_9/GATE sky130_fd_sc_hs__conb_1_131/HI sky130_fd_sc_hs__buf_2_121/X
+ sky130_fd_sc_hs__dlrtp_1_117/a_216_424# sky130_fd_sc_hs__dlrtp_1_117/a_759_508#
+ sky130_fd_sc_hs__dlrtp_1_117/a_565_74# sky130_fd_sc_hs__dlrtp_1_117/a_27_424# sky130_fd_sc_hs__dlrtp_1_117/a_1045_74#
+ sky130_fd_sc_hs__dlrtp_1_117/a_643_74# sky130_fd_sc_hs__dlrtp_1_117/a_817_48# sky130_fd_sc_hs__dlrtp_1_117/a_568_392#
+ sky130_fd_sc_hs__dlrtp_1_117/a_363_74# sky130_fd_sc_hs__dlrtp_1_117/a_769_74# sky130_fd_sc_hs__dlrtp_1
Xsky130_fd_sc_hs__dlrtp_1_127 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__dlrtp_1_127/Q
+ sky130_fd_sc_hs__clkbuf_2_3/A sky130_fd_sc_hs__conb_1_135/HI sky130_fd_sc_hs__buf_2_139/X
+ sky130_fd_sc_hs__dlrtp_1_127/a_216_424# sky130_fd_sc_hs__dlrtp_1_127/a_759_508#
+ sky130_fd_sc_hs__dlrtp_1_127/a_565_74# sky130_fd_sc_hs__dlrtp_1_127/a_27_424# sky130_fd_sc_hs__dlrtp_1_127/a_1045_74#
+ sky130_fd_sc_hs__dlrtp_1_127/a_643_74# sky130_fd_sc_hs__dlrtp_1_127/a_817_48# sky130_fd_sc_hs__dlrtp_1_127/a_568_392#
+ sky130_fd_sc_hs__dlrtp_1_127/a_363_74# sky130_fd_sc_hs__dlrtp_1_127/a_769_74# sky130_fd_sc_hs__dlrtp_1
Xsky130_fd_sc_hs__dlrtp_1_138 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__dlrtp_1_139/Q
+ sky130_fd_sc_hs__clkbuf_16_53/X sky130_fd_sc_hs__conb_1_135/HI sky130_fd_sc_hs__dlrtp_1_139/D
+ sky130_fd_sc_hs__dlrtp_1_139/a_216_424# sky130_fd_sc_hs__dlrtp_1_139/a_759_508#
+ sky130_fd_sc_hs__dlrtp_1_139/a_565_74# sky130_fd_sc_hs__dlrtp_1_139/a_27_424# sky130_fd_sc_hs__dlrtp_1_139/a_1045_74#
+ sky130_fd_sc_hs__dlrtp_1_139/a_643_74# sky130_fd_sc_hs__dlrtp_1_139/a_817_48# sky130_fd_sc_hs__dlrtp_1_139/a_568_392#
+ sky130_fd_sc_hs__dlrtp_1_139/a_363_74# sky130_fd_sc_hs__dlrtp_1_139/a_769_74# sky130_fd_sc_hs__dlrtp_1
Xsky130_fd_sc_hs__dlrtp_1_149 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__dlrtp_1_149/Q
+ sky130_fd_sc_hs__clkbuf_16_53/X sky130_fd_sc_hs__conb_1_127/HI sky130_fd_sc_hs__buf_2_157/X
+ sky130_fd_sc_hs__dlrtp_1_149/a_216_424# sky130_fd_sc_hs__dlrtp_1_149/a_759_508#
+ sky130_fd_sc_hs__dlrtp_1_149/a_565_74# sky130_fd_sc_hs__dlrtp_1_149/a_27_424# sky130_fd_sc_hs__dlrtp_1_149/a_1045_74#
+ sky130_fd_sc_hs__dlrtp_1_149/a_643_74# sky130_fd_sc_hs__dlrtp_1_149/a_817_48# sky130_fd_sc_hs__dlrtp_1_149/a_568_392#
+ sky130_fd_sc_hs__dlrtp_1_149/a_363_74# sky130_fd_sc_hs__dlrtp_1_149/a_769_74# sky130_fd_sc_hs__dlrtp_1
Xsky130_fd_sc_hs__inv_4_8 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__inv_4_9/Y sky130_fd_sc_hs__inv_4_9/A
+ sky130_fd_sc_hs__inv_4
Xsky130_fd_sc_hs__dlrtp_1_40 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__dlrtp_1_41/Q
+ sky130_fd_sc_hs__clkbuf_16_53/A sky130_fd_sc_hs__conb_1_121/HI sky130_fd_sc_hs__buf_2_19/X
+ sky130_fd_sc_hs__dlrtp_1_41/a_216_424# sky130_fd_sc_hs__dlrtp_1_41/a_759_508# sky130_fd_sc_hs__dlrtp_1_41/a_565_74#
+ sky130_fd_sc_hs__dlrtp_1_41/a_27_424# sky130_fd_sc_hs__dlrtp_1_41/a_1045_74# sky130_fd_sc_hs__dlrtp_1_41/a_643_74#
+ sky130_fd_sc_hs__dlrtp_1_41/a_817_48# sky130_fd_sc_hs__dlrtp_1_41/a_568_392# sky130_fd_sc_hs__dlrtp_1_41/a_363_74#
+ sky130_fd_sc_hs__dlrtp_1_41/a_769_74# sky130_fd_sc_hs__dlrtp_1
Xsky130_fd_sc_hs__dlrtp_1_51 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__dlrtp_1_51/Q
+ sky130_fd_sc_hs__clkbuf_16_53/A sky130_fd_sc_hs__conb_1_123/HI sky130_fd_sc_hs__inv_4_11/A
+ sky130_fd_sc_hs__dlrtp_1_51/a_216_424# sky130_fd_sc_hs__dlrtp_1_51/a_759_508# sky130_fd_sc_hs__dlrtp_1_51/a_565_74#
+ sky130_fd_sc_hs__dlrtp_1_51/a_27_424# sky130_fd_sc_hs__dlrtp_1_51/a_1045_74# sky130_fd_sc_hs__dlrtp_1_51/a_643_74#
+ sky130_fd_sc_hs__dlrtp_1_51/a_817_48# sky130_fd_sc_hs__dlrtp_1_51/a_568_392# sky130_fd_sc_hs__dlrtp_1_51/a_363_74#
+ sky130_fd_sc_hs__dlrtp_1_51/a_769_74# sky130_fd_sc_hs__dlrtp_1
Xsky130_fd_sc_hs__dlrtp_1_62 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__dlrtp_1_63/Q
+ sky130_fd_sc_hs__clkbuf_16_53/A sky130_fd_sc_hs__conb_1_125/HI sky130_fd_sc_hs__buf_2_53/X
+ sky130_fd_sc_hs__dlrtp_1_63/a_216_424# sky130_fd_sc_hs__dlrtp_1_63/a_759_508# sky130_fd_sc_hs__dlrtp_1_63/a_565_74#
+ sky130_fd_sc_hs__dlrtp_1_63/a_27_424# sky130_fd_sc_hs__dlrtp_1_63/a_1045_74# sky130_fd_sc_hs__dlrtp_1_63/a_643_74#
+ sky130_fd_sc_hs__dlrtp_1_63/a_817_48# sky130_fd_sc_hs__dlrtp_1_63/a_568_392# sky130_fd_sc_hs__dlrtp_1_63/a_363_74#
+ sky130_fd_sc_hs__dlrtp_1_63/a_769_74# sky130_fd_sc_hs__dlrtp_1
Xsky130_fd_sc_hs__dlrtp_1_73 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__dlrtp_1_75/Q
+ sky130_fd_sc_hs__clkbuf_16_53/X sky130_fd_sc_hs__conb_1_129/HI sky130_fd_sc_hs__buf_2_47/X
+ sky130_fd_sc_hs__dlrtp_1_75/a_216_424# sky130_fd_sc_hs__dlrtp_1_75/a_759_508# sky130_fd_sc_hs__dlrtp_1_75/a_565_74#
+ sky130_fd_sc_hs__dlrtp_1_75/a_27_424# sky130_fd_sc_hs__dlrtp_1_75/a_1045_74# sky130_fd_sc_hs__dlrtp_1_75/a_643_74#
+ sky130_fd_sc_hs__dlrtp_1_75/a_817_48# sky130_fd_sc_hs__dlrtp_1_75/a_568_392# sky130_fd_sc_hs__dlrtp_1_75/a_363_74#
+ sky130_fd_sc_hs__dlrtp_1_75/a_769_74# sky130_fd_sc_hs__dlrtp_1
Xsky130_fd_sc_hs__dlrtp_1_84 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__dlrtp_1_85/Q
+ sky130_fd_sc_hs__clkbuf_16_53/X sky130_fd_sc_hs__conb_1_137/HI sky130_fd_sc_hs__inv_4_17/A
+ sky130_fd_sc_hs__dlrtp_1_85/a_216_424# sky130_fd_sc_hs__dlrtp_1_85/a_759_508# sky130_fd_sc_hs__dlrtp_1_85/a_565_74#
+ sky130_fd_sc_hs__dlrtp_1_85/a_27_424# sky130_fd_sc_hs__dlrtp_1_85/a_1045_74# sky130_fd_sc_hs__dlrtp_1_85/a_643_74#
+ sky130_fd_sc_hs__dlrtp_1_85/a_817_48# sky130_fd_sc_hs__dlrtp_1_85/a_568_392# sky130_fd_sc_hs__dlrtp_1_85/a_363_74#
+ sky130_fd_sc_hs__dlrtp_1_85/a_769_74# sky130_fd_sc_hs__dlrtp_1
Xsky130_fd_sc_hs__dlrtp_1_95 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__dlrtp_1_95/Q
+ sky130_fd_sc_hs__dlrtp_1_9/GATE sky130_fd_sc_hs__conb_1_133/HI sky130_fd_sc_hs__buf_2_101/X
+ sky130_fd_sc_hs__dlrtp_1_95/a_216_424# sky130_fd_sc_hs__dlrtp_1_95/a_759_508# sky130_fd_sc_hs__dlrtp_1_95/a_565_74#
+ sky130_fd_sc_hs__dlrtp_1_95/a_27_424# sky130_fd_sc_hs__dlrtp_1_95/a_1045_74# sky130_fd_sc_hs__dlrtp_1_95/a_643_74#
+ sky130_fd_sc_hs__dlrtp_1_95/a_817_48# sky130_fd_sc_hs__dlrtp_1_95/a_568_392# sky130_fd_sc_hs__dlrtp_1_95/a_363_74#
+ sky130_fd_sc_hs__dlrtp_1_95/a_769_74# sky130_fd_sc_hs__dlrtp_1
Xsky130_fd_sc_hs__einvp_2_0 DVSS: DVDD: DVDD: DVSS: dout_n sky130_fd_sc_hs__einvp_2_9/A
+ sky130_fd_sc_hs__buf_2_99/X sky130_fd_sc_hs__einvp_2_1/a_263_323# sky130_fd_sc_hs__einvp_2_1/a_36_74#
+ sky130_fd_sc_hs__einvp_2_1/a_27_368# sky130_fd_sc_hs__einvp_2
Xsky130_fd_sc_hs__clkbuf_2_3 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__clkbuf_2_3/X
+ sky130_fd_sc_hs__clkbuf_2_3/A sky130_fd_sc_hs__clkbuf_2_3/a_43_192# sky130_fd_sc_hs__clkbuf_2
Xsky130_fd_sc_hs__clkbuf_2_14 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__einvp_2_89/TE
+ sky130_fd_sc_hs__dlrtp_1_85/Q sky130_fd_sc_hs__clkbuf_2_15/a_43_192# sky130_fd_sc_hs__clkbuf_2
Xsky130_fd_sc_hs__clkbuf_2_25 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__dlrtp_1_89/D
+ sky130_fd_sc_hs__o21ai_2_21/Y sky130_fd_sc_hs__clkbuf_2_25/a_43_192# sky130_fd_sc_hs__clkbuf_2
Xsky130_fd_sc_hs__clkbuf_2_36 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__dlrtp_1_98/D
+ sky130_fd_sc_hs__o21bai_2_35/Y sky130_fd_sc_hs__clkbuf_2_37/a_43_192# sky130_fd_sc_hs__clkbuf_2
Xsky130_fd_sc_hs__clkbuf_2_47 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__dlrtp_1_17/D
+ sky130_fd_sc_hs__o21bai_2_41/Y sky130_fd_sc_hs__clkbuf_2_47/a_43_192# sky130_fd_sc_hs__clkbuf_2
Xsky130_fd_sc_hs__clkbuf_2_58 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__dlrtp_1_35/D
+ sky130_fd_sc_hs__o21ai_2_45/Y sky130_fd_sc_hs__clkbuf_2_59/a_43_192# sky130_fd_sc_hs__clkbuf_2
Xsky130_fd_sc_hs__clkbuf_2_69 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__dlrtp_1_153/D
+ sky130_fd_sc_hs__o21bai_2_67/Y sky130_fd_sc_hs__clkbuf_2_69/a_43_192# sky130_fd_sc_hs__clkbuf_2
Xsky130_fd_sc_hs__clkinv_2_3 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__clkinv_2_3/Y
+ sky130_fd_sc_hs__inv_4_7/Y sky130_fd_sc_hs__clkinv_2
Xsky130_fd_sc_hs__buf_2_5 DVSS: DVDD: DVDD: DVSS: manual_control_osc[8] sky130_fd_sc_hs__buf_2_5/X
+ sky130_fd_sc_hs__buf_2_5/a_21_260# sky130_fd_sc_hs__buf_2
Xsky130_fd_sc_hs__dlrtp_1_7 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__dlrtp_1_7/Q sky130_fd_sc_hs__dlrtp_1_9/GATE
+ sky130_fd_sc_hs__conb_1_117/HI sky130_fd_sc_hs__inv_4_21/A sky130_fd_sc_hs__dlrtp_1_7/a_216_424#
+ sky130_fd_sc_hs__dlrtp_1_7/a_759_508# sky130_fd_sc_hs__dlrtp_1_7/a_565_74# sky130_fd_sc_hs__dlrtp_1_7/a_27_424#
+ sky130_fd_sc_hs__dlrtp_1_7/a_1045_74# sky130_fd_sc_hs__dlrtp_1_7/a_643_74# sky130_fd_sc_hs__dlrtp_1_7/a_817_48#
+ sky130_fd_sc_hs__dlrtp_1_7/a_568_392# sky130_fd_sc_hs__dlrtp_1_7/a_363_74# sky130_fd_sc_hs__dlrtp_1_7/a_769_74#
+ sky130_fd_sc_hs__dlrtp_1
Xsky130_fd_sc_hs__buf_2_10 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__buf_2_7/X sky130_fd_sc_hs__buf_2_11/X
+ sky130_fd_sc_hs__buf_2_11/a_21_260# sky130_fd_sc_hs__buf_2
Xsky130_fd_sc_hs__buf_2_21 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__buf_2_25/X sky130_fd_sc_hs__buf_2_21/X
+ sky130_fd_sc_hs__buf_2_21/a_21_260# sky130_fd_sc_hs__buf_2
Xsky130_fd_sc_hs__buf_2_32 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__buf_2_33/A sky130_fd_sc_hs__inv_4_13/A
+ sky130_fd_sc_hs__buf_2_33/a_21_260# sky130_fd_sc_hs__buf_2
Xsky130_fd_sc_hs__buf_2_43 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__buf_2_43/A sky130_fd_sc_hs__buf_2_55/A
+ sky130_fd_sc_hs__buf_2_43/a_21_260# sky130_fd_sc_hs__buf_2
Xsky130_fd_sc_hs__buf_2_54 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__buf_2_55/A sky130_fd_sc_hs__buf_2_55/X
+ sky130_fd_sc_hs__buf_2_55/a_21_260# sky130_fd_sc_hs__buf_2
Xsky130_fd_sc_hs__buf_2_65 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__inv_4_11/Y sky130_fd_sc_hs__buf_2_65/X
+ sky130_fd_sc_hs__buf_2_65/a_21_260# sky130_fd_sc_hs__buf_2
Xsky130_fd_sc_hs__buf_2_76 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__buf_2_77/A sky130_fd_sc_hs__buf_2_77/X
+ sky130_fd_sc_hs__buf_2_77/a_21_260# sky130_fd_sc_hs__buf_2
Xsky130_fd_sc_hs__buf_2_87 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__buf_2_87/A sky130_fd_sc_hs__inv_4_19/A
+ sky130_fd_sc_hs__buf_2_87/a_21_260# sky130_fd_sc_hs__buf_2
Xsky130_fd_sc_hs__buf_2_98 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__buf_2_98/A sky130_fd_sc_hs__buf_2_98/X
+ sky130_fd_sc_hs__buf_2_98/a_21_260# sky130_fd_sc_hs__buf_2
Xsky130_fd_sc_hs__o21bai_2_12 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__nand2_2_7/A
+ sky130_fd_sc_hs__o21bai_2_5/A1 sky130_fd_sc_hs__dlrtp_1_65/D sky130_fd_sc_hs__o21bai_2_13/Y
+ sky130_fd_sc_hs__o21bai_2_13/a_27_74# sky130_fd_sc_hs__o21bai_2_13/a_225_74# sky130_fd_sc_hs__o21bai_2_13/a_507_368#
+ sky130_fd_sc_hs__o21bai_2
Xsky130_fd_sc_hs__o21bai_2_23 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__clkinv_4_3/Y
+ sky130_fd_sc_hs__buf_8_3/X sky130_fd_sc_hs__buf_2_101/X sky130_fd_sc_hs__buf_2_103/A
+ sky130_fd_sc_hs__o21bai_2_23/a_27_74# sky130_fd_sc_hs__o21bai_2_23/a_225_74# sky130_fd_sc_hs__o21bai_2_23/a_507_368#
+ sky130_fd_sc_hs__o21bai_2
Xsky130_fd_sc_hs__o21bai_2_34 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__clkinv_4_5/Y
+ sky130_fd_sc_hs__or2b_2_3/A sky130_fd_sc_hs__buf_2_107/X sky130_fd_sc_hs__o21bai_2_35/Y
+ sky130_fd_sc_hs__o21bai_2_35/a_27_74# sky130_fd_sc_hs__o21bai_2_35/a_225_74# sky130_fd_sc_hs__o21bai_2_35/a_507_368#
+ sky130_fd_sc_hs__o21bai_2
Xsky130_fd_sc_hs__o21bai_2_45 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__clkinv_4_5/Y
+ sky130_fd_sc_hs__nand2_2_15/B sky130_fd_sc_hs__buf_2_121/X sky130_fd_sc_hs__buf_2_117/A
+ sky130_fd_sc_hs__o21bai_2_45/a_27_74# sky130_fd_sc_hs__o21bai_2_45/a_225_74# sky130_fd_sc_hs__o21bai_2_45/a_507_368#
+ sky130_fd_sc_hs__o21bai_2
Xsky130_fd_sc_hs__o21bai_2_56 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__o21ai_2_51/A1
+ sky130_fd_sc_hs__o21bai_4_3/A2 sky130_fd_sc_hs__dlrtp_1_133/D sky130_fd_sc_hs__buf_2_139/A
+ sky130_fd_sc_hs__o21bai_2_57/a_27_74# sky130_fd_sc_hs__o21bai_2_57/a_225_74# sky130_fd_sc_hs__o21bai_2_57/a_507_368#
+ sky130_fd_sc_hs__o21bai_2
Xsky130_fd_sc_hs__o21bai_2_67 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__o21bai_2_5/A1
+ sky130_fd_sc_hs__nand2_2_9/B sky130_fd_sc_hs__buf_2_47/X sky130_fd_sc_hs__o21bai_2_67/Y
+ sky130_fd_sc_hs__o21bai_2_67/a_27_74# sky130_fd_sc_hs__o21bai_2_67/a_225_74# sky130_fd_sc_hs__o21bai_2_67/a_507_368#
+ sky130_fd_sc_hs__o21bai_2
Xsky130_fd_sc_hs__o21bai_4_1 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__buf_2_30/A sky130_fd_sc_hs__inv_8_1/Y
+ sky130_fd_sc_hs__nand2_2_3/B sky130_fd_sc_hs__buf_2_49/X sky130_fd_sc_hs__o21bai_4_1/a_28_368#
+ sky130_fd_sc_hs__o21bai_4_1/a_27_74# sky130_fd_sc_hs__o21bai_4_1/a_828_48# sky130_fd_sc_hs__o21bai_4
Xsky130_fd_sc_hs__conb_1_210 DVSS: DVDD: DVDD: DVSS: prbs_generator_syn_21/eqn[30]
+ sky130_fd_sc_hs__conb_1_211/HI sky130_fd_sc_hs__conb_1_211/a_165_290# sky130_fd_sc_hs__conb_1_211/a_21_290#
+ sky130_fd_sc_hs__conb_1
Xsky130_fd_sc_hs__conb_1_221 DVSS: DVDD: DVDD: DVSS: prbs_generator_syn_25/eqn[31]
+ prbs_generator_syn_25/cke sky130_fd_sc_hs__conb_1_221/a_165_290# sky130_fd_sc_hs__conb_1_221/a_21_290#
+ sky130_fd_sc_hs__conb_1
Xsky130_fd_sc_hs__conb_1_232 DVSS: DVDD: DVDD: DVSS: prbs_generator_syn_27/eqn[9]
+ sky130_fd_sc_hs__conb_1_233/HI sky130_fd_sc_hs__conb_1_233/a_165_290# sky130_fd_sc_hs__conb_1_233/a_21_290#
+ sky130_fd_sc_hs__conb_1
Xsky130_fd_sc_hs__conb_1_243 DVSS: DVDD: DVDD: DVSS: prbs_generator_syn_31/eqn[9]
+ sky130_fd_sc_hs__conb_1_243/HI sky130_fd_sc_hs__conb_1_243/a_165_290# sky130_fd_sc_hs__conb_1_243/a_21_290#
+ sky130_fd_sc_hs__conb_1
Xsky130_fd_sc_hs__conb_1_254 DVSS: DVDD: DVDD: DVSS: prbs_generator_syn_27/eqn[31]
+ prbs_generator_syn_27/cke sky130_fd_sc_hs__conb_1_255/a_165_290# sky130_fd_sc_hs__conb_1_255/a_21_290#
+ sky130_fd_sc_hs__conb_1
Xsky130_fd_sc_hs__conb_1_265 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__conb_1_265/LO
+ sky130_fd_sc_hs__conb_1_265/HI sky130_fd_sc_hs__conb_1_265/a_165_290# sky130_fd_sc_hs__conb_1_265/a_21_290#
+ sky130_fd_sc_hs__conb_1
Xsky130_fd_sc_hs__clkbuf_8_13 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__clkbuf_8_13/X
+ sky130_fd_sc_hs__clkbuf_8_13/A sky130_fd_sc_hs__clkbuf_8_13/a_125_368# sky130_fd_sc_hs__clkbuf_8
Xsky130_fd_sc_hs__clkbuf_8_24 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__clkbuf_8_25/X
+ sky130_fd_sc_hs__clkbuf_8_25/A sky130_fd_sc_hs__clkbuf_8_25/a_125_368# sky130_fd_sc_hs__clkbuf_8
Xsky130_fd_sc_hs__clkbuf_8_35 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__clkbuf_8_35/X
+ sky130_fd_sc_hs__clkbuf_8_35/A sky130_fd_sc_hs__clkbuf_8_35/a_125_368# sky130_fd_sc_hs__clkbuf_8
Xsky130_fd_sc_hs__clkbuf_8_46 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__or2b_2_3/A
+ sky130_fd_sc_hs__nand2_2_29/Y sky130_fd_sc_hs__clkbuf_8_47/a_125_368# sky130_fd_sc_hs__clkbuf_8
Xsky130_fd_sc_hs__clkbuf_8_57 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__o21bai_2_3/A2
+ sky130_fd_sc_hs__nand2_2_33/Y sky130_fd_sc_hs__clkbuf_8_57/a_125_368# sky130_fd_sc_hs__clkbuf_8
Xsky130_fd_sc_hs__clkbuf_8_68 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__or4_2_1/C sky130_fd_sc_hs__clkbuf_8_69/A
+ sky130_fd_sc_hs__clkbuf_8_69/a_125_368# sky130_fd_sc_hs__clkbuf_8
Xsky130_fd_sc_hs__clkbuf_8_79 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__clkbuf_8_79/X
+ sky130_fd_sc_hs__clkbuf_8_79/A sky130_fd_sc_hs__clkbuf_8_79/a_125_368# sky130_fd_sc_hs__clkbuf_8
Xsky130_fd_sc_hs__nand2_2_6 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__nand2_2_7/Y sky130_fd_sc_hs__buf_2_65/X
+ sky130_fd_sc_hs__nand2_2_7/A sky130_fd_sc_hs__nand2_2_7/a_27_74# sky130_fd_sc_hs__nand2_2
Xsky130_fd_sc_hs__or2b_4_2 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__or2b_4_3/A sky130_fd_sc_hs__nor2_4_3/Y
+ sky130_fd_sc_hs__or2b_4_3/X sky130_fd_sc_hs__or2b_4_3/a_676_48# sky130_fd_sc_hs__or2b_4_3/a_489_392#
+ sky130_fd_sc_hs__or2b_4_3/a_81_296# sky130_fd_sc_hs__or2b_4
Xprbs_generator_syn_30 prbs_generator_syn_31/clk prbs_generator_syn_31/rst prbs_generator_syn_31/cke
+ sky130_fd_sc_hs__conb_1_273/LO sky130_fd_sc_hs__conb_1_273/LO sky130_fd_sc_hs__conb_1_273/HI
+ sky130_fd_sc_hs__conb_1_273/HI sky130_fd_sc_hs__conb_1_273/HI sky130_fd_sc_hs__conb_1_273/HI
+ sky130_fd_sc_hs__conb_1_273/HI sky130_fd_sc_hs__conb_1_273/HI sky130_fd_sc_hs__conb_1_273/HI
+ sky130_fd_sc_hs__conb_1_273/LO sky130_fd_sc_hs__conb_1_273/LO prbs_generator_syn_31/eqn[31]
+ prbs_generator_syn_31/cke prbs_generator_syn_31/eqn[31] prbs_generator_syn_31/cke
+ prbs_generator_syn_31/eqn[31] prbs_generator_syn_31/cke prbs_generator_syn_31/cke
+ prbs_generator_syn_31/eqn[1] prbs_generator_syn_31/eqn[1] prbs_generator_syn_31/eqn[1]
+ prbs_generator_syn_31/eqn[1] prbs_generator_syn_31/eqn[1] prbs_generator_syn_31/eqn[2]
+ sky130_fd_sc_hs__conb_1_271/LO sky130_fd_sc_hs__conb_1_271/HI sky130_fd_sc_hs__conb_1_271/HI
+ sky130_fd_sc_hs__conb_1_271/LO sky130_fd_sc_hs__conb_1_271/LO sky130_fd_sc_hs__conb_1_271/HI
+ sky130_fd_sc_hs__conb_1_271/LO sky130_fd_sc_hs__conb_1_271/HI prbs_generator_syn_31/eqn[31]
+ prbs_generator_syn_31/eqn[30] prbs_generator_syn_31/eqn[30] prbs_generator_syn_31/eqn[28]
+ prbs_generator_syn_31/eqn[28] prbs_generator_syn_31/eqn[28] prbs_generator_syn_31/eqn[28]
+ prbs_generator_syn_31/eqn[28] prbs_generator_syn_31/eqn[28] prbs_generator_syn_31/eqn[28]
+ prbs_generator_syn_31/eqn[21] prbs_generator_syn_31/eqn[20] prbs_generator_syn_31/eqn[21]
+ prbs_generator_syn_31/eqn[21] prbs_generator_syn_31/eqn[21] prbs_generator_syn_31/eqn[21]
+ prbs_generator_syn_31/eqn[21] prbs_generator_syn_31/eqn[9] prbs_generator_syn_31/eqn[9]
+ prbs_generator_syn_31/eqn[9] prbs_generator_syn_31/eqn[9] prbs_generator_syn_31/eqn[9]
+ prbs_generator_syn_31/eqn[9] prbs_generator_syn_31/eqn[8] prbs_generator_syn_31/eqn[8]
+ prbs_generator_syn_31/eqn[8] prbs_generator_syn_31/eqn[8] prbs_generator_syn_31/eqn[8]
+ prbs_generator_syn_31/eqn[8] prbs_generator_syn_31/eqn[2] prbs_generator_syn_31/eqn[1]
+ prbs_generator_syn_31/eqn[2] prbs_generator_syn_31/inj_err prbs_generator_syn_31/eqn[31]
+ prbs_generator_syn_31/eqn[31] hr_16t4_mux_top_1/din[8] DVSS: DVDD: prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_1/a_293_74#
+ prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_15/X prbs_generator_syn_31/sky130_fd_sc_hs__nand2_1_35/B
+ prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_51/Y prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_9/A
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_9/CLK prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_47/a_27_74#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_37/a_1226_296# prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_3/B
+ prbs_generator_syn_31/sky130_fd_sc_hs__nor2b_1_7/a_27_112# prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_29/B
+ prbs_generator_syn_31/sky130_fd_sc_hs__sdlclkp_2_1/a_580_74# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_1/a_1141_508#
+ prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_5/Y prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_41/a_230_79#
+ prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_61/a_138_385# prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_43/a_132_392#
+ prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_3/a_222_392# prbs_generator_syn_31/sky130_fd_sc_hs__nor2b_1_9/a_27_112#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_61/a_27_74# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_35/a_206_368#
+ prbs_generator_syn_31/sky130_fd_sc_hs__nand2_2_3/Y prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_25/B
+ prbs_generator_syn_31/sky130_fd_sc_hs__nand2_1_11/a_117_74# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_67/a_651_503#
+ prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_45/X prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_39/a_696_458#
+ prbs_generator_syn_31/sky130_fd_sc_hs__sdlclkp_2_1/a_1198_74# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_45/a_1034_424#
+ prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_17/a_222_392# prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_55/a_222_392#
+ prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_53/Y prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_35/A
+ prbs_generator_syn_31/m3_13600_1651# prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_59/a_52_123#
+ prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_5/a_293_74# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_35/a_1226_296#
+ prbs_generator_syn_31/sky130_fd_sc_hs__nand2_1_51/B prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_5/a_651_503#
+ prbs_generator_syn_31/sky130_fd_sc_hs__nand2_1_21/B prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_8/a_27_74#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_15/a_27_74# prbs_generator_syn_31/sky130_fd_sc_hs__and2b_2_1/X
+ prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_13/X prbs_generator_syn_31/sky130_fd_sc_hs__nand2_2_3/a_27_74#
+ prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_50/a_138_385# prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_33/a_132_392#
+ prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_1/a_376_368# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_25/a_206_368#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_35/a_437_503# prbs_generator_syn_31/sky130_fd_sc_hs__sdlclkp_2_1/a_708_451#
+ prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_45/a_230_79# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_29/a_696_458#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_32/a_27_74# prbs_generator_syn_31/sky130_fd_sc_hs__nor2b_1_4/Y
+ prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_59/a_293_74# prbs_generator_syn_31/sky130_fd_sc_hs__nand2_1_47/a_117_74#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_73/a_735_102# prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_21/a_112_119#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_23/a_1141_508# prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_25/a_293_74#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_7/Q prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_3/a_112_119#
+ prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_35/B prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_51/X
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_53/a_1178_124# prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_23/a_132_392#
+ prbs_generator_syn_31/sky130_fd_sc_hs__nand2_1_3/B prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_15/a_206_368#
+ prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_63/a_132_392# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_55/a_27_74#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_25/a_437_503# prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_41/a_52_123#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_47/a_651_503# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_73/a_1141_508#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_19/a_696_458# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_57/a_696_458#
+ prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_7/X prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_43/a_1034_424#
+ prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_55/A prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_11/a_112_119#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_21/a_1141_508# prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_35/a_222_392#
+ prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_49/a_230_79# prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_67/Y
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_71/a_27_74# prbs_generator_syn_31/sky130_fd_sc_hs__nand2_1_33/B
+ prbs_generator_syn_31/sky130_fd_sc_hs__conb_1_1/LO prbs_generator_syn_31/sky130_fd_sc_hs__nand2_1_19/a_117_74#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_51/a_1178_124# prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_33/X
+ prbs_generator_syn_31/sky130_fd_sc_hs__nand2_1_29/B prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_41/Y
+ prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_53/a_132_392# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_45/a_206_368#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_15/a_437_503# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_37/a_651_503#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_39/a_544_485# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_53/a_735_102#
+ prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_45/a_52_123# prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_1/B
+ prbs_generator_syn_31/sky130_fd_sc_hs__nand2_2_3/B prbs_generator_syn_31/sky130_fd_sc_hs__clkbuf_16_1/A
+ prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_21/X prbs_generator_syn_31/sky130_fd_sc_hs__nand2_1_25/B
+ prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_39/a_376_368# prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_63/X
+ prbs_generator_syn_31/m3_13600_3481# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_69/a_1178_124#
+ prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_21/a_138_385# prbs_generator_syn_31/sky130_fd_sc_hs__nor2b_1_8/Y
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_19/a_1178_124# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_49/a_27_74#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_45/a_437_503# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_27/a_651_503#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_71/a_1141_508# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_65/a_651_503#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_29/a_544_485# prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_3/a_138_385#
+ prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_55/X prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_43/a_735_102#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_41/a_1034_424# prbs_generator_syn_31/sky130_fd_sc_hs__nand2_1_9/B
+ prbs_generator_syn_31/sky130_fd_sc_hs__nor2b_1_9/Y prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_59/a_1034_424#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_39/a_1141_508# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_33/a_1226_296#
+ prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_49/a_52_123# prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_47/Y
+ prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_43/Y prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_4/a_651_503#
+ prbs_generator_syn_31/sky130_fd_sc_hs__nand2_1_49/B prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_19/A
+ prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_11/a_138_385# prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_5/X
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_63/a_206_368# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_17/a_651_503#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_19/a_544_485# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_55/a_651_503#
+ prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_9/Y prbs_generator_syn_31/sky130_fd_sc_hs__nand2_1_17/B
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_57/a_544_485# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_67/a_696_458#
+ prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_35/X prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_19/a_27_74#
+ prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_45/a_222_392# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_32/a_1226_296#
+ prbs_generator_syn_31/sky130_fd_sc_hs__nand2_1_43/B prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_25/A
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_1/a_206_368# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_49/a_1226_296#
+ prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_1/a_112_119# prbs_generator_syn_31/sky130_fd_sc_hs__or2_1_1/X
+ prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_59/a_376_368# prbs_generator_syn_31/sky130_fd_sc_hs__nand2_1_19/B
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_5/a_696_458# prbs_generator_syn_31/sky130_fd_sc_hs__nor2b_1_1/Y
+ prbs_generator_syn_31/sky130_fd_sc_hs__nor2b_1_5/a_278_368# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_17/a_1178_124#
+ prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_39/X prbs_generator_syn_31/m3_13600_5433#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_63/a_437_503# prbs_generator_syn_31/sky130_fd_sc_hs__nand2_2_5/B
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_23/a_735_102# prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_53/A
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_61/a_735_102# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_57/a_1034_424#
+ prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_63/B prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_37/a_1141_508#
+ prbs_generator_syn_31/sky130_fd_sc_hs__nand2_1_47/B prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_29/X
+ prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_65/Y prbs_generator_syn_31/m3_13600_4701#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_1/a_437_503# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_67/a_1178_124#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_9/a_735_102# prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_13/a_132_392#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_15/a_1178_124# prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_15/A
+ prbs_generator_syn_31/sky130_fd_sc_hs__nand2_1_1/B prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_43/B
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_35/a_651_503# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_8/D
+ prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_29/A prbs_generator_syn_31/sky130_fd_sc_hs__nand2_1_7/B
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_13/a_735_102# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_47/a_696_458#
+ prbs_generator_syn_31/sky130_fd_sc_hs__nand2_1_31/B prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_51/a_735_102#
+ prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_59/X prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_35/a_1141_508#
+ prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_25/a_222_392# prbs_generator_syn_31/sky130_fd_sc_hs__sdlclkp_2_1/a_288_48#
+ prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_55/B prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_17/B
+ prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_43/A prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_7/A
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_65/a_1178_124# prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_59/Y
+ prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_41/X prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_21/a_230_79#
+ prbs_generator_syn_31/sky130_fd_sc_hs__nand2_1_57/a_117_74# prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_1/a_222_392#
+ prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_19/B prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_35/a_293_74#
+ prbs_generator_syn_31/sky130_fd_sc_hs__nand2_1_23/a_117_74# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_73/a_206_368#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_25/a_651_503# prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_1/a_138_385#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_37/a_696_458# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_67/a_544_485#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_43/a_27_74# prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_9/X
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_55/a_1034_424# prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_39/a_112_119#
+ prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_15/a_222_392# prbs_generator_syn_31/sky130_fd_sc_hs__conb_1_1/HI
+ prbs_generator_syn_31/sky130_fd_sc_hs__nand2_1_23/B prbs_generator_syn_31/sky130_fd_sc_hs__nand2_1_53/B
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_9/a_1178_124# prbs_generator_syn_31/sky130_fd_sc_hs__nor2b_1_4/A
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_47/a_1226_296# prbs_generator_syn_31/m3_13600_11045#
+ prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_17/X prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_29/a_376_368#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_5/a_544_485# prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_3/X
+ prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_31/a_132_392# prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_61/A
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_15/a_651_503# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_73/a_437_503#
+ prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_25/a_230_79# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_27/a_696_458#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_65/a_696_458# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_33/a_735_102#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_71/a_735_102# prbs_generator_syn_31/m3_13600_7263#
+ prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_43/a_222_392# prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_50/Y
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_8/a_1178_124# prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_53/B
+ prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_19/a_376_368# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_63/a_1178_124#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_4/a_696_458# prbs_generator_syn_31/sky130_fd_sc_hs__nor2b_1_4/a_278_368#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_13/a_1178_124# prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_61/a_132_392#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_53/a_206_368# prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_21/a_52_123#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_45/a_651_503# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_17/a_696_458#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_47/a_544_485# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_55/a_696_458#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_21/a_735_102# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_37/a_27_74#
+ prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_61/B prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_61/X
+ prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_59/a_112_119# prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_31/A
+ prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_33/a_222_392# prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_29/a_230_79#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_45/a_1226_296# prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_9/a_132_392#
+ prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_5/A prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_57/Y
+ prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_31/X prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_51/a_27_74#
+ prbs_generator_syn_31/sky130_fd_sc_hs__nor2b_1_8/a_27_112# prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_47/a_376_368#
+ prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_53/a_293_74# prbs_generator_syn_31/sky130_fd_sc_hs__nand2_1_43/a_117_74#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_8/a_735_102# prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_21/a_293_74#
+ prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_39/a_138_385# prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_63/Y
+ prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_51/a_132_392# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_43/a_206_368#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_53/a_437_503# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_37/a_544_485#
+ prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_57/X prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_53/a_1034_424#
+ prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_25/a_52_123# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_33/a_1141_508#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_63/Q prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_23/a_222_392#
+ prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_63/a_222_392# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_7/a_1178_124#
+ prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_53/X prbs_generator_syn_31/sky130_fd_sc_hs__nand2_2_5/Y
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_61/a_1178_124# prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_1/a_230_79#
+ prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_43/a_230_79# prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_11/a_230_79#
+ prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_41/a_132_392# prbs_generator_syn_31/sky130_fd_sc_hs__nand2_1_13/a_117_74#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_43/a_437_503# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_27/a_544_485#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_63/a_651_503# prbs_generator_syn_31/sky130_fd_sc_hs__nand2_1_7/a_117_74#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_35/a_696_458# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_65/a_544_485#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_51/a_1034_424# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_41/a_735_102#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_32/a_1141_508# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_49/a_1141_508#
+ prbs_generator_syn_31/sky130_fd_sc_hs__nand2_1_55/B prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_53/a_222_392#
+ prbs_generator_syn_31/sky130_fd_sc_hs__sdlclkp_2_1/a_114_112# prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_9/a_293_74#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_43/a_1226_296# prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_29/a_52_123#
+ prbs_generator_syn_31/sky130_fd_sc_hs__nand2_1_37/B prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_1/a_651_503#
+ prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_27/a_376_368# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_4/a_544_485#
+ prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_67/a_376_368# prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_27/X
+ prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_1/X prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_59/a_138_385#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_29/a_1178_124# prbs_generator_syn_31/m3_13600_2871#
+ prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_5/a_230_79# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_23/a_206_368#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_61/a_206_368# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_17/a_544_485#
+ prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_15/a_230_79# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_25/a_696_458#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_55/a_544_485# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_32/a_735_102#
+ prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_29/a_293_74# prbs_generator_syn_31/sky130_fd_sc_hs__nand2_1_17/a_117_74#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_69/a_1034_424# prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_29/a_112_119#
+ prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_37/X prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_31/B
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_19/a_1034_424# prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_33/A
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_9/a_206_368# prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_57/a_376_368#
+ prbs_generator_syn_31/sky130_fd_sc_hs__sdlclkp_2_1/a_706_317# prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_11/B
+ prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_1/a_52_123# prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_39/B
+ prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_21/a_132_392# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_13/a_206_368#
+ prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_43/a_52_123# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_51/a_206_368#
+ prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_47/X prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_23/a_437_503#
+ prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_11/a_52_123# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_61/a_437_503#
+ prbs_generator_syn_31/sky130_fd_sc_hs__nor2b_1_7/Y prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_51/A
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_15/a_696_458# prbs_generator_syn_31/sky130_fd_sc_hs__nor2b_1_5/Y
+ prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_9/a_230_79# prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_25/X
+ prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_19/a_112_119# prbs_generator_syn_31/sky130_fd_sc_hs__nand2_1_45/B
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_5/a_1178_124# prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_19/a_230_79#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_41/a_1226_296# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_59/a_1226_296#
+ prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_63/a_230_79# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_51/Q
+ prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_7/a_132_392# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_9/a_437_503#
+ prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_46/a_376_368# prbs_generator_syn_31/sky130_fd_sc_hs__nand2_1_33/a_117_74#
+ prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_11/a_293_74# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_27/a_1178_124#
+ prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_11/a_132_392# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_13/a_437_503#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_51/a_437_503# prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_5/a_52_123#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_35/a_544_485# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_73/a_651_503#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_45/a_696_458# prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_15/a_52_123#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_47/a_1141_508# prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_47/a_112_119#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_4/a_1178_124# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_17/a_1034_424#
+ prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_23/B prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_37/a_376_368#
+ prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_15/B prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_7/Y
+ prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_29/a_138_385# prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_33/a_230_79#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_25/a_1178_124# prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_47/a_293_74#
+ prbs_generator_syn_31/sky130_fd_sc_hs__nand2_1_37/a_117_74# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_33/a_206_368#
+ prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_15/a_293_74# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_71/a_206_368#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_25/a_544_485# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_67/a_1034_424#
+ prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_13/a_222_392# prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_9/a_52_123#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_15/a_1034_424# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_57/a_1226_296#
+ prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_19/a_52_123# prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_23/X
+ prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_63/a_52_123# prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_19/a_138_385#
+ prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_9/a_376_368# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_21/a_206_368#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_33/a_437_503# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_71/a_437_503#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_53/a_651_503# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_15/a_544_485#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_63/a_696_458# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_65/a_1034_424#
+ prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_19/a_293_74# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_45/a_1141_508#
+ prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_27/a_112_119# prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_67/a_112_119#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_1/a_1178_124# prbs_generator_syn_31/sky130_fd_sc_hs__conb_1_1/a_21_290#
+ prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_63/a_293_74# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_8/a_206_368#
+ prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_17/a_376_368# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_63/a_27_74#
+ prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_21/A prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_55/a_376_368#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_1/a_696_458# prbs_generator_syn_31/sky130_fd_sc_hs__nor2b_1_1/a_278_368#
+ prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_47/a_138_385# prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_33/a_52_123#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_9/a_1034_424# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_21/a_437_503#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_1/a_27_74# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_43/a_651_503#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_1/Q prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_45/a_544_485#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_69/a_735_102# prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_57/a_112_119#
+ prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_31/a_222_392# prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_13/A
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_55/a_1226_296# prbs_generator_syn_31/sky130_fd_sc_hs__nand2_2_5/a_27_74#
+ prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_53/a_230_79# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_8/a_437_503#
+ prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_67/a_293_74# prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_33/a_293_74#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_7/a_735_102# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_23/a_1178_124#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_41/a_206_368# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_8/a_1034_424#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_63/a_1034_424# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_59/a_735_102#
+ prbs_generator_syn_31/sky130_fd_sc_hs__nand2_1_5/B prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_43/a_1141_508#
+ prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_46/a_112_119# prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_61/a_222_392#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_13/a_1034_424# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_73/a_1178_124#
+ prbs_generator_syn_31/sky130_fd_sc_hs__nand2_1_27/B prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_13/B
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_57/a_27_74# prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_57/a_230_79#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_21/a_1178_124# prbs_generator_syn_31/sky130_fd_sc_hs__nor2b_1_1/a_27_112#
+ prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_27/a_138_385# prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_23/a_230_79#
+ prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_67/a_138_385# prbs_generator_syn_31/sky130_fd_sc_hs__nand2_1_41/B
+ prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_9/a_222_392# prbs_generator_syn_31/sky130_fd_sc_hs__nand2_1_27/a_117_74#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_32/a_206_368# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_23/a_651_503#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_41/a_437_503# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_73/a_27_74#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_61/a_651_503# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_63/a_544_485#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_49/a_735_102# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_73/a_696_458#
+ prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_37/a_112_119# prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_51/a_222_392#
+ prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_43/X prbs_generator_syn_31/sky130_fd_sc_hs__nand2_2_1/B
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_9/a_651_503# prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_53/a_52_123#
+ prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_49/X prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_25/a_376_368#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_1/a_544_485# prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_65/a_376_368#
+ prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_57/a_138_385# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_27/a_27_74#
+ prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_39/a_132_392# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_7/a_1034_424#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_13/a_651_503# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_32/a_437_503#
+ prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_27/a_230_79# prbs_generator_syn_31/m3_13600_12265#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_51/a_651_503# prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_59/B
+ prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_47/A prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_61/a_1034_424#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_41/a_1141_508# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_59/a_1141_508#
+ prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_41/a_222_392# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_53/a_1226_296#
+ prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_3/A prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_71/a_1178_124#
+ prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_9/a_112_119# prbs_generator_syn_31/sky130_fd_sc_hs__nand2_1_3/a_117_74#
+ prbs_generator_syn_31/m3_13600_8483# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_39/a_1178_124#
+ prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_57/a_52_123# prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_46/a_138_385#
+ prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_23/a_52_123# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_67/a_27_74#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_53/a_696_458# prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_17/a_112_119#
+ prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_11/A prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_55/a_112_119#
+ prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_1/A prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_51/a_1226_296#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_29/a_1034_424# prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_59/A
+ prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_23/A prbs_generator_syn_31/sky130_fd_sc_hs__nand2_1_39/B
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_5/a_27_74# prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_57/a_293_74#
+ prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_37/a_138_385# prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_59/a_132_392#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_33/a_651_503# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_71/a_651_503#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_43/a_696_458# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_73/a_544_485#
+ prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_27/a_52_123# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_57/a_1141_508#
+ prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_21/a_222_392# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_35/a_27_74#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_69/a_1226_296# prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_37/B
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_19/a_1226_296# prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_35/a_376_368#
+ prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_47/a_230_79# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_37/a_1178_124#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_5/a_1034_424# prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_49/a_132_392#
+ prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_7/a_222_392# prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_27/a_293_74#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_21/a_651_503# prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_9/a_138_385#
+ prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_11/a_222_392# prbs_generator_syn_31/m3_13600_14095#
+ prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_50/A prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_27/a_1034_424#
+ prbs_generator_syn_31/sky130_fd_sc_hs__nand2_1_13/B prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_8/a_651_503#
+ prbs_generator_syn_31/m3_13600_9703# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_35/a_1178_124#
+ prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_17/a_138_385# prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_55/a_138_385#
+ prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_7/a_230_79# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_4/a_1034_424#
+ prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_7/a_376_368# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_69/a_206_368#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_23/a_696_458# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_53/a_544_485#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_39/a_735_102# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_61/a_696_458#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_55/a_1141_508# prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_25/a_112_119#
+ prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_65/a_112_119# prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_43/a_293_74#
+ prbs_generator_syn_31/sky130_fd_sc_hs__nand2_1_57/B prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_25/a_1034_424#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_7/a_206_368# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_17/a_1226_296#
+ prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_15/a_376_368# prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_53/a_376_368#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_9/a_696_458# prbs_generator_syn_31/m3_13600_431#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_45/a_27_74# prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_47/a_52_123#
+ prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_29/a_132_392# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_59/a_206_368#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_69/a_437_503# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_41/a_651_503#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_43/a_544_485# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_13/a_696_458#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_29/a_735_102# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_51/a_696_458#
+ prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_61/Y prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_67/a_1226_296#
+ prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_5/a_132_392# prbs_generator_syn_31/sky130_fd_sc_hs__and2b_2_1/a_198_48#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_7/a_437_503# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_15/a_1226_296#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_69/a_27_74# prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_46/a_293_74#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_1/a_1034_424# prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_19/a_132_392#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_49/a_206_368# prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_7/a_52_123#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_59/a_437_503# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_32/a_651_503#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_7/a_27_74# prbs_generator_syn_31/sky130_fd_sc_hs__nand2_2_1/a_27_74#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_19/a_735_102# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_57/a_735_102#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_65/a_1226_296# prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_37/A
+ prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_33/a_376_368# prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_37/a_230_79#
+ prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_25/a_138_385# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_39/a_27_74#
+ prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_65/a_138_385# prbs_generator_syn_31/sky130_fd_sc_hs__nor2b_1_9/a_278_368#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_49/a_437_503# prbs_generator_syn_31/sky130_fd_sc_hs__and2b_2_1/a_505_74#
+ prbs_generator_syn_31/sky130_fd_sc_hs__nand2_1_51/a_117_74# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_23/a_544_485#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_33/a_696_458# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_61/a_544_485#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_9/a_1226_296# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_53/a_1141_508#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_71/a_696_458# prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_35/a_112_119#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_23/a_1034_424# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_9/a_544_485#
+ prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_63/a_376_368# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_33/a_1178_124#
+ prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_5/a_376_368# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_13/a_544_485#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_73/a_1034_424# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_21/a_696_458#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_51/a_544_485# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_8/a_1226_296#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_51/a_1141_508# prbs_generator_syn_31/sky130_fd_sc_hs__nand2_1_55/a_117_74#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_21/a_1034_424# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_63/a_1226_296#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_23/a_27_74# prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_7/a_112_119#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_13/a_1226_296# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_8/a_696_458#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_32/a_1178_124# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_49/a_1178_124#
+ prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_37/a_52_123# prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_27/a_132_392#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_71/Q prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_67/a_735_102#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_69/a_1141_508# prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_15/a_112_119#
+ prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_53/a_112_119# prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_39/a_222_392#
+ prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_55/a_230_79# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_19/a_1141_508#
+ prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_37/a_293_74# prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_43/a_376_368#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_5/a_735_102# prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_35/a_138_385#
+ prbs_generator_syn_31/sky130_fd_sc_hs__sdlclkp_2_1/a_114_424# prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_57/a_132_392#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_71/a_1034_424# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_7/a_1226_296#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_33/a_544_485# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_41/a_696_458#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_71/a_544_485# prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_21/B
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_61/a_1226_296# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_39/a_1034_424#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_17/a_27_74# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_9/a_27_74#
+ prbs_generator_syn_31/sky130_fd_sc_hs__nor2b_1_5/a_27_112# prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_47/a_132_392#
+ prbs_generator_syn_31/sky130_fd_sc_hs__nor2b_1_8/a_278_368# prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_9/B
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_39/a_206_368# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_33/a_27_74#
+ prbs_generator_syn_31/sky130_fd_sc_hs__nand2_1_41/a_117_74# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_69/a_651_503#
+ prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_51/a_293_74# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_21/a_544_485#
+ prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_7/a_138_385# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_32/a_696_458#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_47/a_735_102# prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_33/a_112_119#
+ prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_59/a_222_392# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_17/a_1141_508#
+ prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_55/a_52_123# prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_3/a_293_74#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_7/a_651_503# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_29/a_1226_296#
+ prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_23/a_376_368# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_8/a_544_485#
+ prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_47/B prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_47/a_1178_124#
+ prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_15/a_138_385# prbs_generator_syn_31/sky130_fd_sc_hs__sdlclkp_2_1/a_1195_374#
+ prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_53/a_138_385# prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_37/a_132_392#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_29/a_206_368# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_39/a_437_503#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_59/a_651_503# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_37/a_735_102#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_67/a_1141_508# prbs_generator_syn_31/sky130_fd_sc_hs__and2b_2_1/a_27_74#
+ prbs_generator_syn_31/sky130_fd_sc_hs__conb_1_1/a_165_290# prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_55/a_293_74#
+ prbs_generator_syn_31/sky130_fd_sc_hs__nand2_1_45/a_117_74# prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_63/a_112_119#
+ prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_49/a_222_392# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_37/a_1034_424#
+ prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_23/a_293_74# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_15/a_1141_508#
+ prbs_generator_syn_31/sky130_fd_sc_hs__nand2_1_5/a_117_74# prbs_generator_syn_31/m3_13600_13485#
+ prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_5/a_112_119# prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_13/a_376_368#
+ prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_51/a_376_368# prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_7/a_293_74#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_19/a_206_368# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_57/a_206_368#
+ prbs_generator_syn_31/sky130_fd_sc_hs__sdlclkp_2_1/a_318_74# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_29/a_437_503#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_49/a_651_503# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_25/a_27_74#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_5/a_1226_296# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_41/a_544_485#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_27/a_735_102# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_65/a_1141_508#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_65/a_735_102# prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_3/a_230_79#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_35/a_1034_424# prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_13/a_230_79#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_41/a_27_74# prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_3/a_132_392#
+ prbs_generator_syn_31/sky130_fd_sc_hs__nand2_1_49/a_117_74# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_27/a_1226_296#
+ prbs_generator_syn_31/sky130_fd_sc_hs__nand2_1_15/a_117_74# prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_41/a_376_368#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_45/a_1178_124# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_4/a_735_102#
+ prbs_generator_syn_31/sky130_fd_sc_hs__nand2_1_9/a_117_74# prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_33/a_138_385#
+ prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_17/a_132_392# prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_55/a_132_392#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_9/a_1141_508# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_19/a_437_503#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_57/a_437_503# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_4/a_1226_296#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_32/a_544_485# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_17/a_735_102#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_55/a_735_102# prbs_generator_syn_31/m3_13600_2261#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_65/a_27_74# prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_29/a_222_392#
+ prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_43/a_112_119# prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_19/X
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_25/a_1226_296# prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_31/a_376_368#
+ prbs_generator_syn_31/sky130_fd_sc_hs__or2_1_1/a_63_368# prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_17/a_230_79#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_4/a_27_74# prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_61/a_230_79#
+ prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_63/a_138_385# prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_5/a_222_392#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_8/a_1141_508# prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_41/a_293_74#
+ prbs_generator_syn_31/sky130_fd_sc_hs__nand2_1_31/a_117_74# prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_5/a_138_385#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_63/a_1141_508# prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_19/a_222_392#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_13/a_1141_508# prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_3/a_52_123#
+ prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_13/a_52_123# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_43/a_1178_124#
+ prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_61/a_376_368# prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_35/a_132_392#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_67/a_206_368# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_1/a_1226_296#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_69/a_696_458# prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_31/a_230_79#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_35/a_735_102# prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_23/a_112_119#
+ prbs_generator_syn_31/sky130_fd_sc_hs__nand2_1_35/a_117_74# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_59/a_27_74#
+ prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_13/a_293_74# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_5/a_206_368#
+ prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_50/a_376_368# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_7/a_696_458#
+ prbs_generator_syn_31/sky130_fd_sc_hs__nor2b_1_7/a_278_368# prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_17/a_52_123#
+ prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_43/a_138_385# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_7/a_1141_508#
+ prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_61/a_52_123# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_67/a_437_503#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_61/a_1141_508# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_25/a_735_102#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_59/a_696_458# prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_13/a_112_119#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_33/a_1034_424# prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_51/a_112_119#
+ prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_35/a_230_79# prbs_generator_syn_31/m3_13600_4091#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_23/a_1226_296# prbs_generator_syn_31/sky130_fd_sc_hs__nand2_1_39/a_117_74#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_29/a_27_74# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_5/a_437_503#
+ prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_17/a_293_74# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_41/a_1178_124#
+ prbs_generator_syn_31/sky130_fd_sc_hs__or2_1_1/a_152_368# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_59/a_1178_124#
+ prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_61/a_293_74# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_47/a_206_368#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_39/a_651_503# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_49/a_696_458#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_15/a_735_102# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_32/a_1034_424#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_73/a_1226_296# prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_27/a_222_392#
+ prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_41/a_112_119# prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_31/a_52_123#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_49/a_1034_424# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_29/a_1141_508#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_21/a_1226_296# prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_39/a_230_79#
+ prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_23/a_138_385# prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_51/a_230_79#
+ prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_45/a_132_392# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_37/a_206_368#
+ prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_65/a_293_74# prbs_generator_syn_31/sky130_fd_sc_hs__nand2_1_53/a_117_74#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_47/a_437_503# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_29/a_651_503#
+ prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_31/a_293_74# prbs_generator_syn_31/sky130_fd_sc_hs__nand2_1_21/a_117_74#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_69/a_544_485# prbs_generator_syn_31/sky130_fd_sc_hs__clkbuf_16_1/a_114_74#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_45/a_735_102# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_13/a_27_74#
+ prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_31/a_112_119# prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_57/a_222_392#
+ prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_35/a_52_123# prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_21/a_376_368#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_7/a_544_485# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_57/a_1178_124#
+ prbs_generator_syn_31/m3_13600_6043# prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_13/a_138_385#
+ prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_51/a_138_385# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_5/a_1141_508#
+ prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_3/a_376_368# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_27/a_206_368#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_65/a_206_368# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_37/a_437_503#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_19/a_651_503# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_57/a_651_503#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_59/a_544_485# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_71/a_1226_296#
+ prbs_generator_syn_31/sky130_fd_sc_hs__nand2_1_25/a_117_74# prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_61/a_112_119#
+ prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_47/a_222_392# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_27/a_1141_508#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_53/a_27_74# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_4/a_206_368#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_39/a_1226_296# prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_11/a_376_368#
+ prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_39/a_52_123# prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_41/a_138_385#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_4/a_1141_508# prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_25/a_132_392#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_17/a_206_368# prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_41/A
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_55/a_206_368# prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_51/a_52_123#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_27/a_437_503# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_65/a_437_503#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_49/a_544_485# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_63/a_735_102#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_47/a_1034_424# prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_50/a_112_119#
+ prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_37/a_222_392# prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_59/a_230_79#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_25/a_1141_508# prbs_generator_syn_31/sky130_fd_sc_hs__nor2b_1_4/a_27_112#
+ prbs_generator_syn_31/sky130_fd_sc_hs__sdlclkp_2_1/a_685_81# prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_1/a_132_392#
+ prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_39/a_293_74# prbs_generator_syn_31/sky130_fd_sc_hs__nand2_1_29/a_117_74#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_4/a_437_503# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_55/a_1178_124#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_21/a_27_74# prbs_generator_syn_31/m3_13600_12875#
+ prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_50/a_293_74# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_1/a_735_102#
+ prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_31/a_138_385# prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_15/a_132_392#
+ prbs_generator_syn_31/sky130_fd_sc_hs__nand2_1_1/a_117_74# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_17/a_437_503#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_55/a_437_503# prbs_generator_syn
Xsky130_fd_sc_hs__buf_2_150 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__buf_2_151/A sky130_fd_sc_hs__buf_2_151/X
+ sky130_fd_sc_hs__buf_2_151/a_21_260# sky130_fd_sc_hs__buf_2
Xsky130_fd_sc_hs__buf_2_161 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__buf_2_161/A sky130_fd_sc_hs__buf_2_161/X
+ sky130_fd_sc_hs__buf_2_161/a_21_260# sky130_fd_sc_hs__buf_2
Xsky130_fd_sc_hs__einvp_2_40 DVSS: DVDD: DVDD: DVSS: dout_n sky130_fd_sc_hs__buf_8_1/A
+ sky130_fd_sc_hs__dlrtp_1_35/Q sky130_fd_sc_hs__einvp_2_41/a_263_323# sky130_fd_sc_hs__einvp_2_41/a_36_74#
+ sky130_fd_sc_hs__einvp_2_41/a_27_368# sky130_fd_sc_hs__einvp_2
Xsky130_fd_sc_hs__einvp_2_51 DVSS: DVDD: DVDD: DVSS: dout_n sky130_fd_sc_hs__buf_8_1/X
+ sky130_fd_sc_hs__dlrtp_1_37/Q sky130_fd_sc_hs__einvp_2_51/a_263_323# sky130_fd_sc_hs__einvp_2_51/a_36_74#
+ sky130_fd_sc_hs__einvp_2_51/a_27_368# sky130_fd_sc_hs__einvp_2
Xsky130_fd_sc_hs__clkbuf_4_7 DVSS: DVDD: DVDD: DVSS: pi2_con[0] sky130_fd_sc_hs__clkbuf_4_7/X
+ sky130_fd_sc_hs__clkbuf_4_7/a_83_270# sky130_fd_sc_hs__clkbuf_4
Xsky130_fd_sc_hs__einvp_2_62 DVSS: DVDD: DVDD: DVSS: dout_p sky130_fd_sc_hs__einvp_2_65/A
+ sky130_fd_sc_hs__dlrtp_1_49/Q sky130_fd_sc_hs__einvp_2_63/a_263_323# sky130_fd_sc_hs__einvp_2_63/a_36_74#
+ sky130_fd_sc_hs__einvp_2_63/a_27_368# sky130_fd_sc_hs__einvp_2
Xsky130_fd_sc_hs__einvp_2_73 DVSS: DVDD: DVDD: DVSS: dout_p sky130_fd_sc_hs__einvp_2_97/A
+ sky130_fd_sc_hs__buf_2_35/X sky130_fd_sc_hs__einvp_2_73/a_263_323# sky130_fd_sc_hs__einvp_2_73/a_36_74#
+ sky130_fd_sc_hs__einvp_2_73/a_27_368# sky130_fd_sc_hs__einvp_2
Xsky130_fd_sc_hs__einvp_2_84 DVSS: DVDD: DVDD: DVSS: dout_p sky130_fd_sc_hs__einvp_2_97/A
+ sky130_fd_sc_hs__dlrtp_1_69/Q sky130_fd_sc_hs__einvp_2_85/a_263_323# sky130_fd_sc_hs__einvp_2_85/a_36_74#
+ sky130_fd_sc_hs__einvp_2_85/a_27_368# sky130_fd_sc_hs__einvp_2
Xsky130_fd_sc_hs__einvp_2_95 DVSS: DVDD: DVDD: DVSS: dout_p sky130_fd_sc_hs__einvp_2_97/A
+ sky130_fd_sc_hs__buf_2_71/X sky130_fd_sc_hs__einvp_2_95/a_263_323# sky130_fd_sc_hs__einvp_2_95/a_36_74#
+ sky130_fd_sc_hs__einvp_2_95/a_27_368# sky130_fd_sc_hs__einvp_2
Xsky130_fd_sc_hs__clkinv_4_7 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__clkinv_4_7/Y
+ sky130_fd_sc_hs__nor4_2_1/B sky130_fd_sc_hs__clkinv_4
Xsky130_fd_sc_hs__and2_2_1 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__and2_2_1/A sky130_fd_sc_hs__and2_2_1/B
+ sky130_fd_sc_hs__inv_4_9/A sky130_fd_sc_hs__and2_2_1/a_31_74# sky130_fd_sc_hs__and2_2_1/a_118_74#
+ sky130_fd_sc_hs__and2_2
Xsky130_fd_sc_hs__conb_1_50 DVSS: DVDD: DVDD: DVSS: prbs_generator_syn_7/eqn[9] sky130_fd_sc_hs__conb_1_51/HI
+ sky130_fd_sc_hs__conb_1_51/a_165_290# sky130_fd_sc_hs__conb_1_51/a_21_290# sky130_fd_sc_hs__conb_1
Xsky130_fd_sc_hs__conb_1_61 DVSS: DVDD: DVDD: DVSS: prbs_generator_syn_7/eqn[8] prbs_generator_syn_7/eqn[1]
+ sky130_fd_sc_hs__conb_1_61/a_165_290# sky130_fd_sc_hs__conb_1_61/a_21_290# sky130_fd_sc_hs__conb_1
Xsky130_fd_sc_hs__conb_1_72 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__conb_1_73/LO
+ sky130_fd_sc_hs__conb_1_73/HI sky130_fd_sc_hs__conb_1_73/a_165_290# sky130_fd_sc_hs__conb_1_73/a_21_290#
+ sky130_fd_sc_hs__conb_1
Xsky130_fd_sc_hs__conb_1_83 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__conb_1_83/LO
+ sky130_fd_sc_hs__conb_1_83/HI sky130_fd_sc_hs__conb_1_83/a_165_290# sky130_fd_sc_hs__conb_1_83/a_21_290#
+ sky130_fd_sc_hs__conb_1
Xsky130_fd_sc_hs__conb_1_94 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__conb_1_95/LO
+ sky130_fd_sc_hs__conb_1_95/HI sky130_fd_sc_hs__conb_1_95/a_165_290# sky130_fd_sc_hs__conb_1_95/a_21_290#
+ sky130_fd_sc_hs__conb_1
Xsky130_fd_sc_hs__dlrtp_1_106 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__einvp_2_27/TE
+ sky130_fd_sc_hs__dlrtp_1_9/GATE sky130_fd_sc_hs__conb_1_133/HI sky130_fd_sc_hs__dlrtp_1_107/D
+ sky130_fd_sc_hs__dlrtp_1_107/a_216_424# sky130_fd_sc_hs__dlrtp_1_107/a_759_508#
+ sky130_fd_sc_hs__dlrtp_1_107/a_565_74# sky130_fd_sc_hs__dlrtp_1_107/a_27_424# sky130_fd_sc_hs__dlrtp_1_107/a_1045_74#
+ sky130_fd_sc_hs__dlrtp_1_107/a_643_74# sky130_fd_sc_hs__dlrtp_1_107/a_817_48# sky130_fd_sc_hs__dlrtp_1_107/a_568_392#
+ sky130_fd_sc_hs__dlrtp_1_107/a_363_74# sky130_fd_sc_hs__dlrtp_1_107/a_769_74# sky130_fd_sc_hs__dlrtp_1
Xsky130_fd_sc_hs__dlrtp_1_117 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__buf_2_119/A
+ sky130_fd_sc_hs__dlrtp_1_9/GATE sky130_fd_sc_hs__conb_1_131/HI sky130_fd_sc_hs__buf_2_121/X
+ sky130_fd_sc_hs__dlrtp_1_117/a_216_424# sky130_fd_sc_hs__dlrtp_1_117/a_759_508#
+ sky130_fd_sc_hs__dlrtp_1_117/a_565_74# sky130_fd_sc_hs__dlrtp_1_117/a_27_424# sky130_fd_sc_hs__dlrtp_1_117/a_1045_74#
+ sky130_fd_sc_hs__dlrtp_1_117/a_643_74# sky130_fd_sc_hs__dlrtp_1_117/a_817_48# sky130_fd_sc_hs__dlrtp_1_117/a_568_392#
+ sky130_fd_sc_hs__dlrtp_1_117/a_363_74# sky130_fd_sc_hs__dlrtp_1_117/a_769_74# sky130_fd_sc_hs__dlrtp_1
Xsky130_fd_sc_hs__dlrtp_1_128 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__buf_2_17/A
+ sky130_fd_sc_hs__clkbuf_2_3/A sky130_fd_sc_hs__conb_1_121/HI sky130_fd_sc_hs__buf_2_137/X
+ sky130_fd_sc_hs__dlrtp_1_129/a_216_424# sky130_fd_sc_hs__dlrtp_1_129/a_759_508#
+ sky130_fd_sc_hs__dlrtp_1_129/a_565_74# sky130_fd_sc_hs__dlrtp_1_129/a_27_424# sky130_fd_sc_hs__dlrtp_1_129/a_1045_74#
+ sky130_fd_sc_hs__dlrtp_1_129/a_643_74# sky130_fd_sc_hs__dlrtp_1_129/a_817_48# sky130_fd_sc_hs__dlrtp_1_129/a_568_392#
+ sky130_fd_sc_hs__dlrtp_1_129/a_363_74# sky130_fd_sc_hs__dlrtp_1_129/a_769_74# sky130_fd_sc_hs__dlrtp_1
Xsky130_fd_sc_hs__dlrtp_1_139 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__dlrtp_1_139/Q
+ sky130_fd_sc_hs__clkbuf_16_53/X sky130_fd_sc_hs__conb_1_135/HI sky130_fd_sc_hs__dlrtp_1_139/D
+ sky130_fd_sc_hs__dlrtp_1_139/a_216_424# sky130_fd_sc_hs__dlrtp_1_139/a_759_508#
+ sky130_fd_sc_hs__dlrtp_1_139/a_565_74# sky130_fd_sc_hs__dlrtp_1_139/a_27_424# sky130_fd_sc_hs__dlrtp_1_139/a_1045_74#
+ sky130_fd_sc_hs__dlrtp_1_139/a_643_74# sky130_fd_sc_hs__dlrtp_1_139/a_817_48# sky130_fd_sc_hs__dlrtp_1_139/a_568_392#
+ sky130_fd_sc_hs__dlrtp_1_139/a_363_74# sky130_fd_sc_hs__dlrtp_1_139/a_769_74# sky130_fd_sc_hs__dlrtp_1
Xsky130_fd_sc_hs__inv_4_9 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__inv_4_9/Y sky130_fd_sc_hs__inv_4_9/A
+ sky130_fd_sc_hs__inv_4
Xsky130_fd_sc_hs__dlrtp_1_30 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__dlrtp_1_31/Q
+ sky130_fd_sc_hs__clkbuf_2_3/A sky130_fd_sc_hs__conb_1_121/HI sky130_fd_sc_hs__buf_2_133/X
+ sky130_fd_sc_hs__dlrtp_1_31/a_216_424# sky130_fd_sc_hs__dlrtp_1_31/a_759_508# sky130_fd_sc_hs__dlrtp_1_31/a_565_74#
+ sky130_fd_sc_hs__dlrtp_1_31/a_27_424# sky130_fd_sc_hs__dlrtp_1_31/a_1045_74# sky130_fd_sc_hs__dlrtp_1_31/a_643_74#
+ sky130_fd_sc_hs__dlrtp_1_31/a_817_48# sky130_fd_sc_hs__dlrtp_1_31/a_568_392# sky130_fd_sc_hs__dlrtp_1_31/a_363_74#
+ sky130_fd_sc_hs__dlrtp_1_31/a_769_74# sky130_fd_sc_hs__dlrtp_1
Xsky130_fd_sc_hs__dlrtp_1_41 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__dlrtp_1_41/Q
+ sky130_fd_sc_hs__clkbuf_16_53/A sky130_fd_sc_hs__conb_1_121/HI sky130_fd_sc_hs__buf_2_19/X
+ sky130_fd_sc_hs__dlrtp_1_41/a_216_424# sky130_fd_sc_hs__dlrtp_1_41/a_759_508# sky130_fd_sc_hs__dlrtp_1_41/a_565_74#
+ sky130_fd_sc_hs__dlrtp_1_41/a_27_424# sky130_fd_sc_hs__dlrtp_1_41/a_1045_74# sky130_fd_sc_hs__dlrtp_1_41/a_643_74#
+ sky130_fd_sc_hs__dlrtp_1_41/a_817_48# sky130_fd_sc_hs__dlrtp_1_41/a_568_392# sky130_fd_sc_hs__dlrtp_1_41/a_363_74#
+ sky130_fd_sc_hs__dlrtp_1_41/a_769_74# sky130_fd_sc_hs__dlrtp_1
Xsky130_fd_sc_hs__dlrtp_1_52 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__dlrtp_1_53/Q
+ sky130_fd_sc_hs__clkbuf_16_53/A sky130_fd_sc_hs__conb_1_123/HI sky130_fd_sc_hs__dlrtp_1_53/D
+ sky130_fd_sc_hs__dlrtp_1_53/a_216_424# sky130_fd_sc_hs__dlrtp_1_53/a_759_508# sky130_fd_sc_hs__dlrtp_1_53/a_565_74#
+ sky130_fd_sc_hs__dlrtp_1_53/a_27_424# sky130_fd_sc_hs__dlrtp_1_53/a_1045_74# sky130_fd_sc_hs__dlrtp_1_53/a_643_74#
+ sky130_fd_sc_hs__dlrtp_1_53/a_817_48# sky130_fd_sc_hs__dlrtp_1_53/a_568_392# sky130_fd_sc_hs__dlrtp_1_53/a_363_74#
+ sky130_fd_sc_hs__dlrtp_1_53/a_769_74# sky130_fd_sc_hs__dlrtp_1
Xsky130_fd_sc_hs__dlrtp_1_63 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__dlrtp_1_63/Q
+ sky130_fd_sc_hs__clkbuf_16_53/A sky130_fd_sc_hs__conb_1_125/HI sky130_fd_sc_hs__buf_2_53/X
+ sky130_fd_sc_hs__dlrtp_1_63/a_216_424# sky130_fd_sc_hs__dlrtp_1_63/a_759_508# sky130_fd_sc_hs__dlrtp_1_63/a_565_74#
+ sky130_fd_sc_hs__dlrtp_1_63/a_27_424# sky130_fd_sc_hs__dlrtp_1_63/a_1045_74# sky130_fd_sc_hs__dlrtp_1_63/a_643_74#
+ sky130_fd_sc_hs__dlrtp_1_63/a_817_48# sky130_fd_sc_hs__dlrtp_1_63/a_568_392# sky130_fd_sc_hs__dlrtp_1_63/a_363_74#
+ sky130_fd_sc_hs__dlrtp_1_63/a_769_74# sky130_fd_sc_hs__dlrtp_1
Xsky130_fd_sc_hs__dlrtp_1_74 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__dlrtp_1_74/Q
+ sky130_fd_sc_hs__clkbuf_16_53/X sky130_fd_sc_hs__conb_1_129/HI sky130_fd_sc_hs__dlrtp_1_74/D
+ sky130_fd_sc_hs__dlrtp_1_74/a_216_424# sky130_fd_sc_hs__dlrtp_1_74/a_759_508# sky130_fd_sc_hs__dlrtp_1_74/a_565_74#
+ sky130_fd_sc_hs__dlrtp_1_74/a_27_424# sky130_fd_sc_hs__dlrtp_1_74/a_1045_74# sky130_fd_sc_hs__dlrtp_1_74/a_643_74#
+ sky130_fd_sc_hs__dlrtp_1_74/a_817_48# sky130_fd_sc_hs__dlrtp_1_74/a_568_392# sky130_fd_sc_hs__dlrtp_1_74/a_363_74#
+ sky130_fd_sc_hs__dlrtp_1_74/a_769_74# sky130_fd_sc_hs__dlrtp_1
Xsky130_fd_sc_hs__dlrtp_1_85 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__dlrtp_1_85/Q
+ sky130_fd_sc_hs__clkbuf_16_53/X sky130_fd_sc_hs__conb_1_137/HI sky130_fd_sc_hs__inv_4_17/A
+ sky130_fd_sc_hs__dlrtp_1_85/a_216_424# sky130_fd_sc_hs__dlrtp_1_85/a_759_508# sky130_fd_sc_hs__dlrtp_1_85/a_565_74#
+ sky130_fd_sc_hs__dlrtp_1_85/a_27_424# sky130_fd_sc_hs__dlrtp_1_85/a_1045_74# sky130_fd_sc_hs__dlrtp_1_85/a_643_74#
+ sky130_fd_sc_hs__dlrtp_1_85/a_817_48# sky130_fd_sc_hs__dlrtp_1_85/a_568_392# sky130_fd_sc_hs__dlrtp_1_85/a_363_74#
+ sky130_fd_sc_hs__dlrtp_1_85/a_769_74# sky130_fd_sc_hs__dlrtp_1
Xsky130_fd_sc_hs__dlrtp_1_96 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__dlrtp_1_97/Q
+ sky130_fd_sc_hs__dlrtp_1_9/GATE sky130_fd_sc_hs__conb_1_133/HI sky130_fd_sc_hs__buf_2_98/X
+ sky130_fd_sc_hs__dlrtp_1_97/a_216_424# sky130_fd_sc_hs__dlrtp_1_97/a_759_508# sky130_fd_sc_hs__dlrtp_1_97/a_565_74#
+ sky130_fd_sc_hs__dlrtp_1_97/a_27_424# sky130_fd_sc_hs__dlrtp_1_97/a_1045_74# sky130_fd_sc_hs__dlrtp_1_97/a_643_74#
+ sky130_fd_sc_hs__dlrtp_1_97/a_817_48# sky130_fd_sc_hs__dlrtp_1_97/a_568_392# sky130_fd_sc_hs__dlrtp_1_97/a_363_74#
+ sky130_fd_sc_hs__dlrtp_1_97/a_769_74# sky130_fd_sc_hs__dlrtp_1
Xsky130_fd_sc_hs__einvp_2_1 DVSS: DVDD: DVDD: DVSS: dout_n sky130_fd_sc_hs__einvp_2_9/A
+ sky130_fd_sc_hs__buf_2_99/X sky130_fd_sc_hs__einvp_2_1/a_263_323# sky130_fd_sc_hs__einvp_2_1/a_36_74#
+ sky130_fd_sc_hs__einvp_2_1/a_27_368# sky130_fd_sc_hs__einvp_2
Xsky130_fd_sc_hs__clkbuf_2_4 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__dlrtp_1_53/D
+ sky130_fd_sc_hs__buf_2_45/X sky130_fd_sc_hs__clkbuf_2_5/a_43_192# sky130_fd_sc_hs__clkbuf_2
Xsky130_fd_sc_hs__clkbuf_2_15 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__einvp_2_89/TE
+ sky130_fd_sc_hs__dlrtp_1_85/Q sky130_fd_sc_hs__clkbuf_2_15/a_43_192# sky130_fd_sc_hs__clkbuf_2
Xsky130_fd_sc_hs__clkbuf_2_26 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__dlrtp_1_79/D
+ sky130_fd_sc_hs__o21ai_2_23/Y sky130_fd_sc_hs__clkbuf_2_28/a_43_192# sky130_fd_sc_hs__clkbuf_2
Xsky130_fd_sc_hs__clkbuf_2_37 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__dlrtp_1_98/D
+ sky130_fd_sc_hs__o21bai_2_35/Y sky130_fd_sc_hs__clkbuf_2_37/a_43_192# sky130_fd_sc_hs__clkbuf_2
Xsky130_fd_sc_hs__clkbuf_2_48 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__dlrtp_1_25/D
+ sky130_fd_sc_hs__o21ai_2_37/Y sky130_fd_sc_hs__clkbuf_2_49/a_43_192# sky130_fd_sc_hs__clkbuf_2
Xsky130_fd_sc_hs__clkbuf_2_59 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__dlrtp_1_35/D
+ sky130_fd_sc_hs__o21ai_2_45/Y sky130_fd_sc_hs__clkbuf_2_59/a_43_192# sky130_fd_sc_hs__clkbuf_2
Xsky130_fd_sc_hs__buf_2_6 DVSS: DVDD: DVDD: DVSS: manual_control_osc[3] sky130_fd_sc_hs__buf_2_7/X
+ sky130_fd_sc_hs__buf_2_7/a_21_260# sky130_fd_sc_hs__buf_2
Xsky130_fd_sc_hs__dlrtp_1_8 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__dlrtp_1_8/Q sky130_fd_sc_hs__dlrtp_1_9/GATE
+ sky130_fd_sc_hs__conb_1_117/HI sky130_fd_sc_hs__dlrtp_1_8/D sky130_fd_sc_hs__dlrtp_1_8/a_216_424#
+ sky130_fd_sc_hs__dlrtp_1_8/a_759_508# sky130_fd_sc_hs__dlrtp_1_8/a_565_74# sky130_fd_sc_hs__dlrtp_1_8/a_27_424#
+ sky130_fd_sc_hs__dlrtp_1_8/a_1045_74# sky130_fd_sc_hs__dlrtp_1_8/a_643_74# sky130_fd_sc_hs__dlrtp_1_8/a_817_48#
+ sky130_fd_sc_hs__dlrtp_1_8/a_568_392# sky130_fd_sc_hs__dlrtp_1_8/a_363_74# sky130_fd_sc_hs__dlrtp_1_8/a_769_74#
+ sky130_fd_sc_hs__dlrtp_1
Xsky130_fd_sc_hs__buf_2_11 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__buf_2_7/X sky130_fd_sc_hs__buf_2_11/X
+ sky130_fd_sc_hs__buf_2_11/a_21_260# sky130_fd_sc_hs__buf_2
Xsky130_fd_sc_hs__buf_2_22 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__buf_2_41/X sky130_fd_sc_hs__buf_2_23/X
+ sky130_fd_sc_hs__buf_2_23/a_21_260# sky130_fd_sc_hs__buf_2
Xsky130_fd_sc_hs__buf_2_33 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__buf_2_33/A sky130_fd_sc_hs__inv_4_13/A
+ sky130_fd_sc_hs__buf_2_33/a_21_260# sky130_fd_sc_hs__buf_2
Xsky130_fd_sc_hs__buf_2_44 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__buf_2_45/A sky130_fd_sc_hs__buf_2_45/X
+ sky130_fd_sc_hs__buf_2_45/a_21_260# sky130_fd_sc_hs__buf_2
Xsky130_fd_sc_hs__buf_2_55 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__buf_2_55/A sky130_fd_sc_hs__buf_2_55/X
+ sky130_fd_sc_hs__buf_2_55/a_21_260# sky130_fd_sc_hs__buf_2
Xsky130_fd_sc_hs__buf_2_66 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__buf_2_67/A sky130_fd_sc_hs__buf_2_67/X
+ sky130_fd_sc_hs__buf_2_67/a_21_260# sky130_fd_sc_hs__buf_2
Xsky130_fd_sc_hs__buf_2_77 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__buf_2_77/A sky130_fd_sc_hs__buf_2_77/X
+ sky130_fd_sc_hs__buf_2_77/a_21_260# sky130_fd_sc_hs__buf_2
Xsky130_fd_sc_hs__buf_2_88 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__buf_2_89/A sky130_fd_sc_hs__buf_2_89/X
+ sky130_fd_sc_hs__buf_2_89/a_21_260# sky130_fd_sc_hs__buf_2
Xsky130_fd_sc_hs__buf_2_99 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__buf_2_99/A sky130_fd_sc_hs__buf_2_99/X
+ sky130_fd_sc_hs__buf_2_99/a_21_260# sky130_fd_sc_hs__buf_2
Xsky130_fd_sc_hs__o21bai_2_13 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__nand2_2_7/A
+ sky130_fd_sc_hs__o21bai_2_5/A1 sky130_fd_sc_hs__dlrtp_1_65/D sky130_fd_sc_hs__o21bai_2_13/Y
+ sky130_fd_sc_hs__o21bai_2_13/a_27_74# sky130_fd_sc_hs__o21bai_2_13/a_225_74# sky130_fd_sc_hs__o21bai_2_13/a_507_368#
+ sky130_fd_sc_hs__o21bai_2
Xsky130_fd_sc_hs__o21bai_2_24 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__buf_8_3/X sky130_fd_sc_hs__clkbuf_4_81/X
+ sky130_fd_sc_hs__buf_2_101/X sky130_fd_sc_hs__buf_2_98/A sky130_fd_sc_hs__o21bai_2_25/a_27_74#
+ sky130_fd_sc_hs__o21bai_2_25/a_225_74# sky130_fd_sc_hs__o21bai_2_25/a_507_368# sky130_fd_sc_hs__o21bai_2
Xsky130_fd_sc_hs__o21bai_2_35 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__clkinv_4_5/Y
+ sky130_fd_sc_hs__or2b_2_3/A sky130_fd_sc_hs__buf_2_107/X sky130_fd_sc_hs__o21bai_2_35/Y
+ sky130_fd_sc_hs__o21bai_2_35/a_27_74# sky130_fd_sc_hs__o21bai_2_35/a_225_74# sky130_fd_sc_hs__o21bai_2_35/a_507_368#
+ sky130_fd_sc_hs__o21bai_2
Xsky130_fd_sc_hs__o21bai_2_46 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__clkinv_4_3/Y
+ sky130_fd_sc_hs__or2b_2_1/X sky130_fd_sc_hs__dlrtp_1_115/D sky130_fd_sc_hs__buf_2_121/A
+ sky130_fd_sc_hs__o21bai_2_47/a_27_74# sky130_fd_sc_hs__o21bai_2_47/a_225_74# sky130_fd_sc_hs__o21bai_2_47/a_507_368#
+ sky130_fd_sc_hs__o21bai_2
Xsky130_fd_sc_hs__o21bai_2_57 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__o21ai_2_51/A1
+ sky130_fd_sc_hs__o21bai_4_3/A2 sky130_fd_sc_hs__dlrtp_1_133/D sky130_fd_sc_hs__buf_2_139/A
+ sky130_fd_sc_hs__o21bai_2_57/a_27_74# sky130_fd_sc_hs__o21bai_2_57/a_225_74# sky130_fd_sc_hs__o21bai_2_57/a_507_368#
+ sky130_fd_sc_hs__o21bai_2
Xsky130_fd_sc_hs__o21bai_2_68 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__inv_8_1/Y sky130_fd_sc_hs__nand2_2_9/B
+ sky130_fd_sc_hs__dlrtp_1_153/D sky130_fd_sc_hs__o21bai_2_69/Y sky130_fd_sc_hs__o21bai_2_69/a_27_74#
+ sky130_fd_sc_hs__o21bai_2_69/a_225_74# sky130_fd_sc_hs__o21bai_2_69/a_507_368# sky130_fd_sc_hs__o21bai_2
Xsky130_fd_sc_hs__o21bai_4_2 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__o21bai_4_3/Y
+ sky130_fd_sc_hs__nand2_2_15/B sky130_fd_sc_hs__o21bai_4_3/A2 sky130_fd_sc_hs__dlrtp_1_25/D
+ sky130_fd_sc_hs__o21bai_4_3/a_28_368# sky130_fd_sc_hs__o21bai_4_3/a_27_74# sky130_fd_sc_hs__o21bai_4_3/a_828_48#
+ sky130_fd_sc_hs__o21bai_4
Xsky130_fd_sc_hs__conb_1_200 DVSS: DVDD: DVDD: DVSS: prbs_generator_syn_19/eqn[30]
+ sky130_fd_sc_hs__conb_1_201/HI sky130_fd_sc_hs__conb_1_201/a_165_290# sky130_fd_sc_hs__conb_1_201/a_21_290#
+ sky130_fd_sc_hs__conb_1
Xsky130_fd_sc_hs__conb_1_211 DVSS: DVDD: DVDD: DVSS: prbs_generator_syn_21/eqn[30]
+ sky130_fd_sc_hs__conb_1_211/HI sky130_fd_sc_hs__conb_1_211/a_165_290# sky130_fd_sc_hs__conb_1_211/a_21_290#
+ sky130_fd_sc_hs__conb_1
Xsky130_fd_sc_hs__conb_1_222 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__conb_1_223/LO
+ sky130_fd_sc_hs__conb_1_223/HI sky130_fd_sc_hs__conb_1_223/a_165_290# sky130_fd_sc_hs__conb_1_223/a_21_290#
+ sky130_fd_sc_hs__conb_1
Xsky130_fd_sc_hs__conb_1_233 DVSS: DVDD: DVDD: DVSS: prbs_generator_syn_27/eqn[9]
+ sky130_fd_sc_hs__conb_1_233/HI sky130_fd_sc_hs__conb_1_233/a_165_290# sky130_fd_sc_hs__conb_1_233/a_21_290#
+ sky130_fd_sc_hs__conb_1
Xsky130_fd_sc_hs__conb_1_244 DVSS: DVDD: DVDD: DVSS: prbs_generator_syn_31/eqn[21]
+ prbs_generator_syn_31/eqn[20] sky130_fd_sc_hs__conb_1_245/a_165_290# sky130_fd_sc_hs__conb_1_245/a_21_290#
+ sky130_fd_sc_hs__conb_1
Xsky130_fd_sc_hs__conb_1_255 DVSS: DVDD: DVDD: DVSS: prbs_generator_syn_27/eqn[31]
+ prbs_generator_syn_27/cke sky130_fd_sc_hs__conb_1_255/a_165_290# sky130_fd_sc_hs__conb_1_255/a_21_290#
+ sky130_fd_sc_hs__conb_1
Xsky130_fd_sc_hs__conb_1_266 DVSS: DVDD: DVDD: DVSS: prbs_generator_syn_31/eqn[8]
+ sky130_fd_sc_hs__conb_1_267/HI sky130_fd_sc_hs__conb_1_267/a_165_290# sky130_fd_sc_hs__conb_1_267/a_21_290#
+ sky130_fd_sc_hs__conb_1
Xsky130_fd_sc_hs__clkbuf_8_14 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__clkbuf_8_15/X
+ sky130_fd_sc_hs__clkbuf_8_15/A sky130_fd_sc_hs__clkbuf_8_15/a_125_368# sky130_fd_sc_hs__clkbuf_8
Xsky130_fd_sc_hs__clkbuf_8_25 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__clkbuf_8_25/X
+ sky130_fd_sc_hs__clkbuf_8_25/A sky130_fd_sc_hs__clkbuf_8_25/a_125_368# sky130_fd_sc_hs__clkbuf_8
Xsky130_fd_sc_hs__clkbuf_8_36 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__nand2_2_15/B
+ sky130_fd_sc_hs__or2b_2_1/X sky130_fd_sc_hs__clkbuf_8_37/a_125_368# sky130_fd_sc_hs__clkbuf_8
Xsky130_fd_sc_hs__clkbuf_8_47 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__or2b_2_3/A
+ sky130_fd_sc_hs__nand2_2_29/Y sky130_fd_sc_hs__clkbuf_8_47/a_125_368# sky130_fd_sc_hs__clkbuf_8
Xsky130_fd_sc_hs__clkbuf_8_58 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__or4_2_1/A sky130_fd_sc_hs__clkbuf_8_59/A
+ sky130_fd_sc_hs__clkbuf_8_59/a_125_368# sky130_fd_sc_hs__clkbuf_8
Xsky130_fd_sc_hs__clkbuf_8_69 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__or4_2_1/C sky130_fd_sc_hs__clkbuf_8_69/A
+ sky130_fd_sc_hs__clkbuf_8_69/a_125_368# sky130_fd_sc_hs__clkbuf_8
Xsky130_fd_sc_hs__nand2_2_7 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__nand2_2_7/Y sky130_fd_sc_hs__buf_2_65/X
+ sky130_fd_sc_hs__nand2_2_7/A sky130_fd_sc_hs__nand2_2_7/a_27_74# sky130_fd_sc_hs__nand2_2
Xsky130_fd_sc_hs__or2b_4_3 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__or2b_4_3/A sky130_fd_sc_hs__nor2_4_3/Y
+ sky130_fd_sc_hs__or2b_4_3/X sky130_fd_sc_hs__or2b_4_3/a_676_48# sky130_fd_sc_hs__or2b_4_3/a_489_392#
+ sky130_fd_sc_hs__or2b_4_3/a_81_296# sky130_fd_sc_hs__or2b_4
Xprbs_generator_syn_20 prbs_generator_syn_31/clk prbs_generator_syn_31/rst prbs_generator_syn_21/cke
+ sky130_fd_sc_hs__conb_1_223/LO sky130_fd_sc_hs__conb_1_223/LO sky130_fd_sc_hs__conb_1_223/LO
+ prbs_generator_syn_25/eqn[1] prbs_generator_syn_25/eqn[1] prbs_generator_syn_25/eqn[1]
+ prbs_generator_syn_25/eqn[1] prbs_generator_syn_25/eqn[1] sky130_fd_sc_hs__conb_1_223/LO
+ sky130_fd_sc_hs__conb_1_223/LO sky130_fd_sc_hs__conb_1_223/LO prbs_generator_syn_21/eqn[31]
+ prbs_generator_syn_25/eqn[9] sky130_fd_sc_hs__conb_1_215/HI prbs_generator_syn_25/eqn[9]
+ sky130_fd_sc_hs__conb_1_215/HI prbs_generator_syn_25/eqn[9] prbs_generator_syn_21/cke
+ prbs_generator_syn_21/eqn[0] prbs_generator_syn_23/eqn[20] prbs_generator_syn_23/eqn[22]
+ prbs_generator_syn_23/eqn[20] prbs_generator_syn_23/eqn[22] sky130_fd_sc_hs__conb_1_181/HI
+ sky130_fd_sc_hs__conb_1_181/HI prbs_generator_syn_23/eqn[28] prbs_generator_syn_23/eqn[28]
+ sky130_fd_sc_hs__conb_1_227/HI sky130_fd_sc_hs__conb_1_227/HI sky130_fd_sc_hs__conb_1_227/HI
+ sky130_fd_sc_hs__conb_1_227/HI sky130_fd_sc_hs__conb_1_227/HI prbs_generator_syn_21/eqn[31]
+ prbs_generator_syn_21/eqn[30] prbs_generator_syn_21/eqn[30] prbs_generator_syn_21/eqn[30]
+ prbs_generator_syn_21/eqn[30] prbs_generator_syn_21/eqn[30] prbs_generator_syn_21/eqn[30]
+ prbs_generator_syn_21/eqn[30] prbs_generator_syn_21/eqn[30] prbs_generator_syn_21/eqn[22]
+ prbs_generator_syn_21/eqn[22] prbs_generator_syn_21/eqn[20] prbs_generator_syn_21/eqn[22]
+ prbs_generator_syn_21/eqn[22] prbs_generator_syn_21/eqn[22] prbs_generator_syn_21/eqn[22]
+ prbs_generator_syn_21/eqn[22] prbs_generator_syn_21/eqn[22] prbs_generator_syn_21/eqn[9]
+ prbs_generator_syn_21/eqn[9] prbs_generator_syn_21/eqn[9] prbs_generator_syn_21/eqn[9]
+ prbs_generator_syn_21/eqn[9] prbs_generator_syn_21/eqn[8] prbs_generator_syn_21/eqn[8]
+ prbs_generator_syn_21/eqn[8] prbs_generator_syn_21/eqn[8] prbs_generator_syn_21/eqn[8]
+ prbs_generator_syn_21/eqn[8] prbs_generator_syn_21/eqn[8] prbs_generator_syn_21/eqn[1]
+ prbs_generator_syn_21/eqn[0] prbs_generator_syn_31/inj_err prbs_generator_syn_21/eqn[31]
+ prbs_generator_syn_21/eqn[31] prbs_generator_syn_21/out DVSS: DVDD: prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_1/a_293_74#
+ prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_15/X prbs_generator_syn_21/sky130_fd_sc_hs__nand2_1_35/B
+ prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_51/Y prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_9/A
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_9/CLK prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_47/a_27_74#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_37/a_1226_296# prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_3/B
+ prbs_generator_syn_21/sky130_fd_sc_hs__nor2b_1_7/a_27_112# prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_29/B
+ prbs_generator_syn_21/sky130_fd_sc_hs__sdlclkp_2_1/a_580_74# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_1/a_1141_508#
+ prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_5/Y prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_41/a_230_79#
+ prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_61/a_138_385# prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_43/a_132_392#
+ prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_3/a_222_392# prbs_generator_syn_21/sky130_fd_sc_hs__nor2b_1_9/a_27_112#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_61/a_27_74# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_35/a_206_368#
+ prbs_generator_syn_21/sky130_fd_sc_hs__nand2_2_3/Y prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_25/B
+ prbs_generator_syn_21/sky130_fd_sc_hs__nand2_1_11/a_117_74# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_67/a_651_503#
+ prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_45/X prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_39/a_696_458#
+ prbs_generator_syn_21/sky130_fd_sc_hs__sdlclkp_2_1/a_1198_74# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_45/a_1034_424#
+ prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_17/a_222_392# prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_55/a_222_392#
+ prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_53/Y prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_35/A
+ prbs_generator_syn_21/m3_13600_1651# prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_59/a_52_123#
+ prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_5/a_293_74# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_35/a_1226_296#
+ prbs_generator_syn_21/sky130_fd_sc_hs__nand2_1_51/B prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_5/a_651_503#
+ prbs_generator_syn_21/sky130_fd_sc_hs__nand2_1_21/B prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_8/a_27_74#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_15/a_27_74# prbs_generator_syn_21/sky130_fd_sc_hs__and2b_2_1/X
+ prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_13/X prbs_generator_syn_21/sky130_fd_sc_hs__nand2_2_3/a_27_74#
+ prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_50/a_138_385# prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_33/a_132_392#
+ prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_1/a_376_368# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_25/a_206_368#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_35/a_437_503# prbs_generator_syn_21/sky130_fd_sc_hs__sdlclkp_2_1/a_708_451#
+ prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_45/a_230_79# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_29/a_696_458#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_32/a_27_74# prbs_generator_syn_21/sky130_fd_sc_hs__nor2b_1_4/Y
+ prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_59/a_293_74# prbs_generator_syn_21/sky130_fd_sc_hs__nand2_1_47/a_117_74#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_73/a_735_102# prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_21/a_112_119#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_23/a_1141_508# prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_25/a_293_74#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_7/Q prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_3/a_112_119#
+ prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_35/B prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_51/X
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_53/a_1178_124# prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_23/a_132_392#
+ prbs_generator_syn_21/sky130_fd_sc_hs__nand2_1_3/B prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_15/a_206_368#
+ prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_63/a_132_392# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_55/a_27_74#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_25/a_437_503# prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_41/a_52_123#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_47/a_651_503# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_73/a_1141_508#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_19/a_696_458# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_57/a_696_458#
+ prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_7/X prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_43/a_1034_424#
+ prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_55/A prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_11/a_112_119#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_21/a_1141_508# prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_35/a_222_392#
+ prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_49/a_230_79# prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_67/Y
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_71/a_27_74# prbs_generator_syn_21/sky130_fd_sc_hs__nand2_1_33/B
+ prbs_generator_syn_21/sky130_fd_sc_hs__conb_1_1/LO prbs_generator_syn_21/sky130_fd_sc_hs__nand2_1_19/a_117_74#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_51/a_1178_124# prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_33/X
+ prbs_generator_syn_21/sky130_fd_sc_hs__nand2_1_29/B prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_41/Y
+ prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_53/a_132_392# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_45/a_206_368#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_15/a_437_503# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_37/a_651_503#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_39/a_544_485# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_53/a_735_102#
+ prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_45/a_52_123# prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_1/B
+ prbs_generator_syn_21/sky130_fd_sc_hs__nand2_2_3/B prbs_generator_syn_21/sky130_fd_sc_hs__clkbuf_16_1/A
+ prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_21/X prbs_generator_syn_21/sky130_fd_sc_hs__nand2_1_25/B
+ prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_39/a_376_368# prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_63/X
+ prbs_generator_syn_21/m3_13600_3481# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_69/a_1178_124#
+ prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_21/a_138_385# prbs_generator_syn_21/sky130_fd_sc_hs__nor2b_1_8/Y
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_19/a_1178_124# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_49/a_27_74#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_45/a_437_503# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_27/a_651_503#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_71/a_1141_508# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_65/a_651_503#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_29/a_544_485# prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_3/a_138_385#
+ prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_55/X prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_43/a_735_102#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_41/a_1034_424# prbs_generator_syn_21/sky130_fd_sc_hs__nand2_1_9/B
+ prbs_generator_syn_21/sky130_fd_sc_hs__nor2b_1_9/Y prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_59/a_1034_424#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_39/a_1141_508# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_33/a_1226_296#
+ prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_49/a_52_123# prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_47/Y
+ prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_43/Y prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_4/a_651_503#
+ prbs_generator_syn_21/sky130_fd_sc_hs__nand2_1_49/B prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_19/A
+ prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_11/a_138_385# prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_5/X
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_63/a_206_368# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_17/a_651_503#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_19/a_544_485# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_55/a_651_503#
+ prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_9/Y prbs_generator_syn_21/sky130_fd_sc_hs__nand2_1_17/B
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_57/a_544_485# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_67/a_696_458#
+ prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_35/X prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_19/a_27_74#
+ prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_45/a_222_392# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_32/a_1226_296#
+ prbs_generator_syn_21/sky130_fd_sc_hs__nand2_1_43/B prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_25/A
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_1/a_206_368# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_49/a_1226_296#
+ prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_1/a_112_119# prbs_generator_syn_21/sky130_fd_sc_hs__or2_1_1/X
+ prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_59/a_376_368# prbs_generator_syn_21/sky130_fd_sc_hs__nand2_1_19/B
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_5/a_696_458# prbs_generator_syn_21/sky130_fd_sc_hs__nor2b_1_1/Y
+ prbs_generator_syn_21/sky130_fd_sc_hs__nor2b_1_5/a_278_368# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_17/a_1178_124#
+ prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_39/X prbs_generator_syn_21/m3_13600_5433#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_63/a_437_503# prbs_generator_syn_21/sky130_fd_sc_hs__nand2_2_5/B
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_23/a_735_102# prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_53/A
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_61/a_735_102# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_57/a_1034_424#
+ prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_63/B prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_37/a_1141_508#
+ prbs_generator_syn_21/sky130_fd_sc_hs__nand2_1_47/B prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_29/X
+ prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_65/Y prbs_generator_syn_21/m3_13600_4701#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_1/a_437_503# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_67/a_1178_124#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_9/a_735_102# prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_13/a_132_392#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_15/a_1178_124# prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_15/A
+ prbs_generator_syn_21/sky130_fd_sc_hs__nand2_1_1/B prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_43/B
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_35/a_651_503# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_8/D
+ prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_29/A prbs_generator_syn_21/sky130_fd_sc_hs__nand2_1_7/B
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_13/a_735_102# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_47/a_696_458#
+ prbs_generator_syn_21/sky130_fd_sc_hs__nand2_1_31/B prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_51/a_735_102#
+ prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_59/X prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_35/a_1141_508#
+ prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_25/a_222_392# prbs_generator_syn_21/sky130_fd_sc_hs__sdlclkp_2_1/a_288_48#
+ prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_55/B prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_17/B
+ prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_43/A prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_7/A
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_65/a_1178_124# prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_59/Y
+ prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_41/X prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_21/a_230_79#
+ prbs_generator_syn_21/sky130_fd_sc_hs__nand2_1_57/a_117_74# prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_1/a_222_392#
+ prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_19/B prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_35/a_293_74#
+ prbs_generator_syn_21/sky130_fd_sc_hs__nand2_1_23/a_117_74# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_73/a_206_368#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_25/a_651_503# prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_1/a_138_385#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_37/a_696_458# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_67/a_544_485#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_43/a_27_74# prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_9/X
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_55/a_1034_424# prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_39/a_112_119#
+ prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_15/a_222_392# prbs_generator_syn_21/sky130_fd_sc_hs__conb_1_1/HI
+ prbs_generator_syn_21/sky130_fd_sc_hs__nand2_1_23/B prbs_generator_syn_21/sky130_fd_sc_hs__nand2_1_53/B
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_9/a_1178_124# prbs_generator_syn_21/sky130_fd_sc_hs__nor2b_1_4/A
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_47/a_1226_296# prbs_generator_syn_21/m3_13600_11045#
+ prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_17/X prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_29/a_376_368#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_5/a_544_485# prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_3/X
+ prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_31/a_132_392# prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_61/A
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_15/a_651_503# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_73/a_437_503#
+ prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_25/a_230_79# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_27/a_696_458#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_65/a_696_458# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_33/a_735_102#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_71/a_735_102# prbs_generator_syn_21/m3_13600_7263#
+ prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_43/a_222_392# prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_50/Y
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_8/a_1178_124# prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_53/B
+ prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_19/a_376_368# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_63/a_1178_124#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_4/a_696_458# prbs_generator_syn_21/sky130_fd_sc_hs__nor2b_1_4/a_278_368#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_13/a_1178_124# prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_61/a_132_392#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_53/a_206_368# prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_21/a_52_123#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_45/a_651_503# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_17/a_696_458#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_47/a_544_485# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_55/a_696_458#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_21/a_735_102# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_37/a_27_74#
+ prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_61/B prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_61/X
+ prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_59/a_112_119# prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_31/A
+ prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_33/a_222_392# prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_29/a_230_79#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_45/a_1226_296# prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_9/a_132_392#
+ prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_5/A prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_57/Y
+ prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_31/X prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_51/a_27_74#
+ prbs_generator_syn_21/sky130_fd_sc_hs__nor2b_1_8/a_27_112# prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_47/a_376_368#
+ prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_53/a_293_74# prbs_generator_syn_21/sky130_fd_sc_hs__nand2_1_43/a_117_74#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_8/a_735_102# prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_21/a_293_74#
+ prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_39/a_138_385# prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_63/Y
+ prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_51/a_132_392# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_43/a_206_368#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_53/a_437_503# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_37/a_544_485#
+ prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_57/X prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_53/a_1034_424#
+ prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_25/a_52_123# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_33/a_1141_508#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_63/Q prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_23/a_222_392#
+ prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_63/a_222_392# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_7/a_1178_124#
+ prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_53/X prbs_generator_syn_21/sky130_fd_sc_hs__nand2_2_5/Y
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_61/a_1178_124# prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_1/a_230_79#
+ prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_43/a_230_79# prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_11/a_230_79#
+ prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_41/a_132_392# prbs_generator_syn_21/sky130_fd_sc_hs__nand2_1_13/a_117_74#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_43/a_437_503# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_27/a_544_485#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_63/a_651_503# prbs_generator_syn_21/sky130_fd_sc_hs__nand2_1_7/a_117_74#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_35/a_696_458# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_65/a_544_485#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_51/a_1034_424# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_41/a_735_102#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_32/a_1141_508# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_49/a_1141_508#
+ prbs_generator_syn_21/sky130_fd_sc_hs__nand2_1_55/B prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_53/a_222_392#
+ prbs_generator_syn_21/sky130_fd_sc_hs__sdlclkp_2_1/a_114_112# prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_9/a_293_74#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_43/a_1226_296# prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_29/a_52_123#
+ prbs_generator_syn_21/sky130_fd_sc_hs__nand2_1_37/B prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_1/a_651_503#
+ prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_27/a_376_368# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_4/a_544_485#
+ prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_67/a_376_368# prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_27/X
+ prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_1/X prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_59/a_138_385#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_29/a_1178_124# prbs_generator_syn_21/m3_13600_2871#
+ prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_5/a_230_79# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_23/a_206_368#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_61/a_206_368# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_17/a_544_485#
+ prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_15/a_230_79# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_25/a_696_458#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_55/a_544_485# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_32/a_735_102#
+ prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_29/a_293_74# prbs_generator_syn_21/sky130_fd_sc_hs__nand2_1_17/a_117_74#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_69/a_1034_424# prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_29/a_112_119#
+ prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_37/X prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_31/B
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_19/a_1034_424# prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_33/A
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_9/a_206_368# prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_57/a_376_368#
+ prbs_generator_syn_21/sky130_fd_sc_hs__sdlclkp_2_1/a_706_317# prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_11/B
+ prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_1/a_52_123# prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_39/B
+ prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_21/a_132_392# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_13/a_206_368#
+ prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_43/a_52_123# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_51/a_206_368#
+ prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_47/X prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_23/a_437_503#
+ prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_11/a_52_123# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_61/a_437_503#
+ prbs_generator_syn_21/sky130_fd_sc_hs__nor2b_1_7/Y prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_51/A
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_15/a_696_458# prbs_generator_syn_21/sky130_fd_sc_hs__nor2b_1_5/Y
+ prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_9/a_230_79# prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_25/X
+ prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_19/a_112_119# prbs_generator_syn_21/sky130_fd_sc_hs__nand2_1_45/B
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_5/a_1178_124# prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_19/a_230_79#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_41/a_1226_296# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_59/a_1226_296#
+ prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_63/a_230_79# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_51/Q
+ prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_7/a_132_392# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_9/a_437_503#
+ prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_46/a_376_368# prbs_generator_syn_21/sky130_fd_sc_hs__nand2_1_33/a_117_74#
+ prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_11/a_293_74# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_27/a_1178_124#
+ prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_11/a_132_392# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_13/a_437_503#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_51/a_437_503# prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_5/a_52_123#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_35/a_544_485# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_73/a_651_503#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_45/a_696_458# prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_15/a_52_123#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_47/a_1141_508# prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_47/a_112_119#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_4/a_1178_124# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_17/a_1034_424#
+ prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_23/B prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_37/a_376_368#
+ prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_15/B prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_7/Y
+ prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_29/a_138_385# prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_33/a_230_79#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_25/a_1178_124# prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_47/a_293_74#
+ prbs_generator_syn_21/sky130_fd_sc_hs__nand2_1_37/a_117_74# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_33/a_206_368#
+ prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_15/a_293_74# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_71/a_206_368#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_25/a_544_485# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_67/a_1034_424#
+ prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_13/a_222_392# prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_9/a_52_123#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_15/a_1034_424# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_57/a_1226_296#
+ prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_19/a_52_123# prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_23/X
+ prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_63/a_52_123# prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_19/a_138_385#
+ prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_9/a_376_368# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_21/a_206_368#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_33/a_437_503# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_71/a_437_503#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_53/a_651_503# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_15/a_544_485#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_63/a_696_458# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_65/a_1034_424#
+ prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_19/a_293_74# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_45/a_1141_508#
+ prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_27/a_112_119# prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_67/a_112_119#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_1/a_1178_124# prbs_generator_syn_21/sky130_fd_sc_hs__conb_1_1/a_21_290#
+ prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_63/a_293_74# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_8/a_206_368#
+ prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_17/a_376_368# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_63/a_27_74#
+ prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_21/A prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_55/a_376_368#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_1/a_696_458# prbs_generator_syn_21/sky130_fd_sc_hs__nor2b_1_1/a_278_368#
+ prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_47/a_138_385# prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_33/a_52_123#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_9/a_1034_424# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_21/a_437_503#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_1/a_27_74# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_43/a_651_503#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_1/Q prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_45/a_544_485#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_69/a_735_102# prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_57/a_112_119#
+ prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_31/a_222_392# prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_13/A
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_55/a_1226_296# prbs_generator_syn_21/sky130_fd_sc_hs__nand2_2_5/a_27_74#
+ prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_53/a_230_79# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_8/a_437_503#
+ prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_67/a_293_74# prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_33/a_293_74#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_7/a_735_102# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_23/a_1178_124#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_41/a_206_368# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_8/a_1034_424#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_63/a_1034_424# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_59/a_735_102#
+ prbs_generator_syn_21/sky130_fd_sc_hs__nand2_1_5/B prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_43/a_1141_508#
+ prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_46/a_112_119# prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_61/a_222_392#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_13/a_1034_424# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_73/a_1178_124#
+ prbs_generator_syn_21/sky130_fd_sc_hs__nand2_1_27/B prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_13/B
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_57/a_27_74# prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_57/a_230_79#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_21/a_1178_124# prbs_generator_syn_21/sky130_fd_sc_hs__nor2b_1_1/a_27_112#
+ prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_27/a_138_385# prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_23/a_230_79#
+ prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_67/a_138_385# prbs_generator_syn_21/sky130_fd_sc_hs__nand2_1_41/B
+ prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_9/a_222_392# prbs_generator_syn_21/sky130_fd_sc_hs__nand2_1_27/a_117_74#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_32/a_206_368# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_23/a_651_503#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_41/a_437_503# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_73/a_27_74#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_61/a_651_503# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_63/a_544_485#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_49/a_735_102# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_73/a_696_458#
+ prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_37/a_112_119# prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_51/a_222_392#
+ prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_43/X prbs_generator_syn_21/sky130_fd_sc_hs__nand2_2_1/B
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_9/a_651_503# prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_53/a_52_123#
+ prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_49/X prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_25/a_376_368#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_1/a_544_485# prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_65/a_376_368#
+ prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_57/a_138_385# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_27/a_27_74#
+ prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_39/a_132_392# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_7/a_1034_424#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_13/a_651_503# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_32/a_437_503#
+ prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_27/a_230_79# prbs_generator_syn_21/m3_13600_12265#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_51/a_651_503# prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_59/B
+ prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_47/A prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_61/a_1034_424#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_41/a_1141_508# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_59/a_1141_508#
+ prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_41/a_222_392# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_53/a_1226_296#
+ prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_3/A prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_71/a_1178_124#
+ prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_9/a_112_119# prbs_generator_syn_21/sky130_fd_sc_hs__nand2_1_3/a_117_74#
+ prbs_generator_syn_21/m3_13600_8483# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_39/a_1178_124#
+ prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_57/a_52_123# prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_46/a_138_385#
+ prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_23/a_52_123# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_67/a_27_74#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_53/a_696_458# prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_17/a_112_119#
+ prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_11/A prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_55/a_112_119#
+ prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_1/A prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_51/a_1226_296#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_29/a_1034_424# prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_59/A
+ prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_23/A prbs_generator_syn_21/sky130_fd_sc_hs__nand2_1_39/B
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_5/a_27_74# prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_57/a_293_74#
+ prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_37/a_138_385# prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_59/a_132_392#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_33/a_651_503# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_71/a_651_503#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_43/a_696_458# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_73/a_544_485#
+ prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_27/a_52_123# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_57/a_1141_508#
+ prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_21/a_222_392# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_35/a_27_74#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_69/a_1226_296# prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_37/B
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_19/a_1226_296# prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_35/a_376_368#
+ prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_47/a_230_79# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_37/a_1178_124#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_5/a_1034_424# prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_49/a_132_392#
+ prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_7/a_222_392# prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_27/a_293_74#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_21/a_651_503# prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_9/a_138_385#
+ prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_11/a_222_392# prbs_generator_syn_21/m3_13600_14095#
+ prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_50/A prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_27/a_1034_424#
+ prbs_generator_syn_21/sky130_fd_sc_hs__nand2_1_13/B prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_8/a_651_503#
+ prbs_generator_syn_21/m3_13600_9703# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_35/a_1178_124#
+ prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_17/a_138_385# prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_55/a_138_385#
+ prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_7/a_230_79# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_4/a_1034_424#
+ prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_7/a_376_368# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_69/a_206_368#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_23/a_696_458# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_53/a_544_485#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_39/a_735_102# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_61/a_696_458#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_55/a_1141_508# prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_25/a_112_119#
+ prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_65/a_112_119# prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_43/a_293_74#
+ prbs_generator_syn_21/sky130_fd_sc_hs__nand2_1_57/B prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_25/a_1034_424#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_7/a_206_368# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_17/a_1226_296#
+ prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_15/a_376_368# prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_53/a_376_368#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_9/a_696_458# prbs_generator_syn_21/m3_13600_431#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_45/a_27_74# prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_47/a_52_123#
+ prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_29/a_132_392# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_59/a_206_368#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_69/a_437_503# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_41/a_651_503#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_43/a_544_485# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_13/a_696_458#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_29/a_735_102# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_51/a_696_458#
+ prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_61/Y prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_67/a_1226_296#
+ prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_5/a_132_392# prbs_generator_syn_21/sky130_fd_sc_hs__and2b_2_1/a_198_48#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_7/a_437_503# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_15/a_1226_296#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_69/a_27_74# prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_46/a_293_74#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_1/a_1034_424# prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_19/a_132_392#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_49/a_206_368# prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_7/a_52_123#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_59/a_437_503# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_32/a_651_503#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_7/a_27_74# prbs_generator_syn_21/sky130_fd_sc_hs__nand2_2_1/a_27_74#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_19/a_735_102# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_57/a_735_102#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_65/a_1226_296# prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_37/A
+ prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_33/a_376_368# prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_37/a_230_79#
+ prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_25/a_138_385# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_39/a_27_74#
+ prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_65/a_138_385# prbs_generator_syn_21/sky130_fd_sc_hs__nor2b_1_9/a_278_368#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_49/a_437_503# prbs_generator_syn_21/sky130_fd_sc_hs__and2b_2_1/a_505_74#
+ prbs_generator_syn_21/sky130_fd_sc_hs__nand2_1_51/a_117_74# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_23/a_544_485#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_33/a_696_458# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_61/a_544_485#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_9/a_1226_296# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_53/a_1141_508#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_71/a_696_458# prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_35/a_112_119#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_23/a_1034_424# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_9/a_544_485#
+ prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_63/a_376_368# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_33/a_1178_124#
+ prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_5/a_376_368# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_13/a_544_485#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_73/a_1034_424# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_21/a_696_458#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_51/a_544_485# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_8/a_1226_296#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_51/a_1141_508# prbs_generator_syn_21/sky130_fd_sc_hs__nand2_1_55/a_117_74#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_21/a_1034_424# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_63/a_1226_296#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_23/a_27_74# prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_7/a_112_119#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_13/a_1226_296# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_8/a_696_458#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_32/a_1178_124# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_49/a_1178_124#
+ prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_37/a_52_123# prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_27/a_132_392#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_71/Q prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_67/a_735_102#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_69/a_1141_508# prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_15/a_112_119#
+ prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_53/a_112_119# prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_39/a_222_392#
+ prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_55/a_230_79# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_19/a_1141_508#
+ prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_37/a_293_74# prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_43/a_376_368#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_5/a_735_102# prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_35/a_138_385#
+ prbs_generator_syn_21/sky130_fd_sc_hs__sdlclkp_2_1/a_114_424# prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_57/a_132_392#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_71/a_1034_424# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_7/a_1226_296#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_33/a_544_485# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_41/a_696_458#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_71/a_544_485# prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_21/B
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_61/a_1226_296# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_39/a_1034_424#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_17/a_27_74# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_9/a_27_74#
+ prbs_generator_syn_21/sky130_fd_sc_hs__nor2b_1_5/a_27_112# prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_47/a_132_392#
+ prbs_generator_syn_21/sky130_fd_sc_hs__nor2b_1_8/a_278_368# prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_9/B
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_39/a_206_368# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_33/a_27_74#
+ prbs_generator_syn_21/sky130_fd_sc_hs__nand2_1_41/a_117_74# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_69/a_651_503#
+ prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_51/a_293_74# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_21/a_544_485#
+ prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_7/a_138_385# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_32/a_696_458#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_47/a_735_102# prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_33/a_112_119#
+ prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_59/a_222_392# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_17/a_1141_508#
+ prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_55/a_52_123# prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_3/a_293_74#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_7/a_651_503# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_29/a_1226_296#
+ prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_23/a_376_368# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_8/a_544_485#
+ prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_47/B prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_47/a_1178_124#
+ prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_15/a_138_385# prbs_generator_syn_21/sky130_fd_sc_hs__sdlclkp_2_1/a_1195_374#
+ prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_53/a_138_385# prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_37/a_132_392#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_29/a_206_368# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_39/a_437_503#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_59/a_651_503# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_37/a_735_102#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_67/a_1141_508# prbs_generator_syn_21/sky130_fd_sc_hs__and2b_2_1/a_27_74#
+ prbs_generator_syn_21/sky130_fd_sc_hs__conb_1_1/a_165_290# prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_55/a_293_74#
+ prbs_generator_syn_21/sky130_fd_sc_hs__nand2_1_45/a_117_74# prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_63/a_112_119#
+ prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_49/a_222_392# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_37/a_1034_424#
+ prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_23/a_293_74# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_15/a_1141_508#
+ prbs_generator_syn_21/sky130_fd_sc_hs__nand2_1_5/a_117_74# prbs_generator_syn_21/m3_13600_13485#
+ prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_5/a_112_119# prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_13/a_376_368#
+ prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_51/a_376_368# prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_7/a_293_74#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_19/a_206_368# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_57/a_206_368#
+ prbs_generator_syn_21/sky130_fd_sc_hs__sdlclkp_2_1/a_318_74# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_29/a_437_503#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_49/a_651_503# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_25/a_27_74#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_5/a_1226_296# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_41/a_544_485#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_27/a_735_102# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_65/a_1141_508#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_65/a_735_102# prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_3/a_230_79#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_35/a_1034_424# prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_13/a_230_79#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_41/a_27_74# prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_3/a_132_392#
+ prbs_generator_syn_21/sky130_fd_sc_hs__nand2_1_49/a_117_74# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_27/a_1226_296#
+ prbs_generator_syn_21/sky130_fd_sc_hs__nand2_1_15/a_117_74# prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_41/a_376_368#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_45/a_1178_124# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_4/a_735_102#
+ prbs_generator_syn_21/sky130_fd_sc_hs__nand2_1_9/a_117_74# prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_33/a_138_385#
+ prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_17/a_132_392# prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_55/a_132_392#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_9/a_1141_508# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_19/a_437_503#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_57/a_437_503# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_4/a_1226_296#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_32/a_544_485# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_17/a_735_102#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_55/a_735_102# prbs_generator_syn_21/m3_13600_2261#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_65/a_27_74# prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_29/a_222_392#
+ prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_43/a_112_119# prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_19/X
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_25/a_1226_296# prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_31/a_376_368#
+ prbs_generator_syn_21/sky130_fd_sc_hs__or2_1_1/a_63_368# prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_17/a_230_79#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_4/a_27_74# prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_61/a_230_79#
+ prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_63/a_138_385# prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_5/a_222_392#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_8/a_1141_508# prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_41/a_293_74#
+ prbs_generator_syn_21/sky130_fd_sc_hs__nand2_1_31/a_117_74# prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_5/a_138_385#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_63/a_1141_508# prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_19/a_222_392#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_13/a_1141_508# prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_3/a_52_123#
+ prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_13/a_52_123# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_43/a_1178_124#
+ prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_61/a_376_368# prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_35/a_132_392#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_67/a_206_368# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_1/a_1226_296#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_69/a_696_458# prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_31/a_230_79#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_35/a_735_102# prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_23/a_112_119#
+ prbs_generator_syn_21/sky130_fd_sc_hs__nand2_1_35/a_117_74# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_59/a_27_74#
+ prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_13/a_293_74# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_5/a_206_368#
+ prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_50/a_376_368# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_7/a_696_458#
+ prbs_generator_syn_21/sky130_fd_sc_hs__nor2b_1_7/a_278_368# prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_17/a_52_123#
+ prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_43/a_138_385# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_7/a_1141_508#
+ prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_61/a_52_123# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_67/a_437_503#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_61/a_1141_508# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_25/a_735_102#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_59/a_696_458# prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_13/a_112_119#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_33/a_1034_424# prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_51/a_112_119#
+ prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_35/a_230_79# prbs_generator_syn_21/m3_13600_4091#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_23/a_1226_296# prbs_generator_syn_21/sky130_fd_sc_hs__nand2_1_39/a_117_74#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_29/a_27_74# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_5/a_437_503#
+ prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_17/a_293_74# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_41/a_1178_124#
+ prbs_generator_syn_21/sky130_fd_sc_hs__or2_1_1/a_152_368# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_59/a_1178_124#
+ prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_61/a_293_74# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_47/a_206_368#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_39/a_651_503# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_49/a_696_458#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_15/a_735_102# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_32/a_1034_424#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_73/a_1226_296# prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_27/a_222_392#
+ prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_41/a_112_119# prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_31/a_52_123#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_49/a_1034_424# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_29/a_1141_508#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_21/a_1226_296# prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_39/a_230_79#
+ prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_23/a_138_385# prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_51/a_230_79#
+ prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_45/a_132_392# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_37/a_206_368#
+ prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_65/a_293_74# prbs_generator_syn_21/sky130_fd_sc_hs__nand2_1_53/a_117_74#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_47/a_437_503# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_29/a_651_503#
+ prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_31/a_293_74# prbs_generator_syn_21/sky130_fd_sc_hs__nand2_1_21/a_117_74#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_69/a_544_485# prbs_generator_syn_21/sky130_fd_sc_hs__clkbuf_16_1/a_114_74#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_45/a_735_102# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_13/a_27_74#
+ prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_31/a_112_119# prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_57/a_222_392#
+ prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_35/a_52_123# prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_21/a_376_368#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_7/a_544_485# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_57/a_1178_124#
+ prbs_generator_syn_21/m3_13600_6043# prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_13/a_138_385#
+ prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_51/a_138_385# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_5/a_1141_508#
+ prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_3/a_376_368# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_27/a_206_368#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_65/a_206_368# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_37/a_437_503#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_19/a_651_503# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_57/a_651_503#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_59/a_544_485# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_71/a_1226_296#
+ prbs_generator_syn_21/sky130_fd_sc_hs__nand2_1_25/a_117_74# prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_61/a_112_119#
+ prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_47/a_222_392# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_27/a_1141_508#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_53/a_27_74# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_4/a_206_368#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_39/a_1226_296# prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_11/a_376_368#
+ prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_39/a_52_123# prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_41/a_138_385#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_4/a_1141_508# prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_25/a_132_392#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_17/a_206_368# prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_41/A
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_55/a_206_368# prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_51/a_52_123#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_27/a_437_503# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_65/a_437_503#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_49/a_544_485# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_63/a_735_102#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_47/a_1034_424# prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_50/a_112_119#
+ prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_37/a_222_392# prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_59/a_230_79#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_25/a_1141_508# prbs_generator_syn_21/sky130_fd_sc_hs__nor2b_1_4/a_27_112#
+ prbs_generator_syn_21/sky130_fd_sc_hs__sdlclkp_2_1/a_685_81# prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_1/a_132_392#
+ prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_39/a_293_74# prbs_generator_syn_21/sky130_fd_sc_hs__nand2_1_29/a_117_74#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_4/a_437_503# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_55/a_1178_124#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_21/a_27_74# prbs_generator_syn_21/m3_13600_12875#
+ prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_50/a_293_74# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_1/a_735_102#
+ prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_31/a_138_385# prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_15/a_132_392#
+ prbs_generator_syn_21/sky130_fd_sc_hs__nand2_1_1/a_117_74# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_17/a_437_503#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_55/a_437_503# prbs_generator_syn
Xsky130_fd_sc_hs__conb_1_0 DVSS: DVDD: DVDD: DVSS: prbs_generator_syn_1/eqn[9] sky130_fd_sc_hs__conb_1_1/HI
+ sky130_fd_sc_hs__conb_1_1/a_165_290# sky130_fd_sc_hs__conb_1_1/a_21_290# sky130_fd_sc_hs__conb_1
Xprbs_generator_syn_31 prbs_generator_syn_31/clk prbs_generator_syn_31/rst prbs_generator_syn_31/cke
+ sky130_fd_sc_hs__conb_1_273/LO sky130_fd_sc_hs__conb_1_273/LO sky130_fd_sc_hs__conb_1_273/HI
+ sky130_fd_sc_hs__conb_1_273/HI sky130_fd_sc_hs__conb_1_273/HI sky130_fd_sc_hs__conb_1_273/HI
+ sky130_fd_sc_hs__conb_1_273/HI sky130_fd_sc_hs__conb_1_273/HI sky130_fd_sc_hs__conb_1_273/HI
+ sky130_fd_sc_hs__conb_1_273/LO sky130_fd_sc_hs__conb_1_273/LO prbs_generator_syn_31/eqn[31]
+ prbs_generator_syn_31/cke prbs_generator_syn_31/eqn[31] prbs_generator_syn_31/cke
+ prbs_generator_syn_31/eqn[31] prbs_generator_syn_31/cke prbs_generator_syn_31/cke
+ prbs_generator_syn_31/eqn[1] prbs_generator_syn_31/eqn[1] prbs_generator_syn_31/eqn[1]
+ prbs_generator_syn_31/eqn[1] prbs_generator_syn_31/eqn[1] prbs_generator_syn_31/eqn[2]
+ sky130_fd_sc_hs__conb_1_271/LO sky130_fd_sc_hs__conb_1_271/HI sky130_fd_sc_hs__conb_1_271/HI
+ sky130_fd_sc_hs__conb_1_271/LO sky130_fd_sc_hs__conb_1_271/LO sky130_fd_sc_hs__conb_1_271/HI
+ sky130_fd_sc_hs__conb_1_271/LO sky130_fd_sc_hs__conb_1_271/HI prbs_generator_syn_31/eqn[31]
+ prbs_generator_syn_31/eqn[30] prbs_generator_syn_31/eqn[30] prbs_generator_syn_31/eqn[28]
+ prbs_generator_syn_31/eqn[28] prbs_generator_syn_31/eqn[28] prbs_generator_syn_31/eqn[28]
+ prbs_generator_syn_31/eqn[28] prbs_generator_syn_31/eqn[28] prbs_generator_syn_31/eqn[28]
+ prbs_generator_syn_31/eqn[21] prbs_generator_syn_31/eqn[20] prbs_generator_syn_31/eqn[21]
+ prbs_generator_syn_31/eqn[21] prbs_generator_syn_31/eqn[21] prbs_generator_syn_31/eqn[21]
+ prbs_generator_syn_31/eqn[21] prbs_generator_syn_31/eqn[9] prbs_generator_syn_31/eqn[9]
+ prbs_generator_syn_31/eqn[9] prbs_generator_syn_31/eqn[9] prbs_generator_syn_31/eqn[9]
+ prbs_generator_syn_31/eqn[9] prbs_generator_syn_31/eqn[8] prbs_generator_syn_31/eqn[8]
+ prbs_generator_syn_31/eqn[8] prbs_generator_syn_31/eqn[8] prbs_generator_syn_31/eqn[8]
+ prbs_generator_syn_31/eqn[8] prbs_generator_syn_31/eqn[2] prbs_generator_syn_31/eqn[1]
+ prbs_generator_syn_31/eqn[2] prbs_generator_syn_31/inj_err prbs_generator_syn_31/eqn[31]
+ prbs_generator_syn_31/eqn[31] hr_16t4_mux_top_1/din[8] DVSS: DVDD: prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_1/a_293_74#
+ prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_15/X prbs_generator_syn_31/sky130_fd_sc_hs__nand2_1_35/B
+ prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_51/Y prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_9/A
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_9/CLK prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_47/a_27_74#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_37/a_1226_296# prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_3/B
+ prbs_generator_syn_31/sky130_fd_sc_hs__nor2b_1_7/a_27_112# prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_29/B
+ prbs_generator_syn_31/sky130_fd_sc_hs__sdlclkp_2_1/a_580_74# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_1/a_1141_508#
+ prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_5/Y prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_41/a_230_79#
+ prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_61/a_138_385# prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_43/a_132_392#
+ prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_3/a_222_392# prbs_generator_syn_31/sky130_fd_sc_hs__nor2b_1_9/a_27_112#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_61/a_27_74# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_35/a_206_368#
+ prbs_generator_syn_31/sky130_fd_sc_hs__nand2_2_3/Y prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_25/B
+ prbs_generator_syn_31/sky130_fd_sc_hs__nand2_1_11/a_117_74# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_67/a_651_503#
+ prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_45/X prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_39/a_696_458#
+ prbs_generator_syn_31/sky130_fd_sc_hs__sdlclkp_2_1/a_1198_74# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_45/a_1034_424#
+ prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_17/a_222_392# prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_55/a_222_392#
+ prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_53/Y prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_35/A
+ prbs_generator_syn_31/m3_13600_1651# prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_59/a_52_123#
+ prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_5/a_293_74# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_35/a_1226_296#
+ prbs_generator_syn_31/sky130_fd_sc_hs__nand2_1_51/B prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_5/a_651_503#
+ prbs_generator_syn_31/sky130_fd_sc_hs__nand2_1_21/B prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_8/a_27_74#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_15/a_27_74# prbs_generator_syn_31/sky130_fd_sc_hs__and2b_2_1/X
+ prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_13/X prbs_generator_syn_31/sky130_fd_sc_hs__nand2_2_3/a_27_74#
+ prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_50/a_138_385# prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_33/a_132_392#
+ prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_1/a_376_368# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_25/a_206_368#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_35/a_437_503# prbs_generator_syn_31/sky130_fd_sc_hs__sdlclkp_2_1/a_708_451#
+ prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_45/a_230_79# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_29/a_696_458#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_32/a_27_74# prbs_generator_syn_31/sky130_fd_sc_hs__nor2b_1_4/Y
+ prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_59/a_293_74# prbs_generator_syn_31/sky130_fd_sc_hs__nand2_1_47/a_117_74#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_73/a_735_102# prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_21/a_112_119#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_23/a_1141_508# prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_25/a_293_74#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_7/Q prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_3/a_112_119#
+ prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_35/B prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_51/X
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_53/a_1178_124# prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_23/a_132_392#
+ prbs_generator_syn_31/sky130_fd_sc_hs__nand2_1_3/B prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_15/a_206_368#
+ prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_63/a_132_392# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_55/a_27_74#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_25/a_437_503# prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_41/a_52_123#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_47/a_651_503# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_73/a_1141_508#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_19/a_696_458# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_57/a_696_458#
+ prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_7/X prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_43/a_1034_424#
+ prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_55/A prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_11/a_112_119#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_21/a_1141_508# prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_35/a_222_392#
+ prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_49/a_230_79# prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_67/Y
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_71/a_27_74# prbs_generator_syn_31/sky130_fd_sc_hs__nand2_1_33/B
+ prbs_generator_syn_31/sky130_fd_sc_hs__conb_1_1/LO prbs_generator_syn_31/sky130_fd_sc_hs__nand2_1_19/a_117_74#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_51/a_1178_124# prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_33/X
+ prbs_generator_syn_31/sky130_fd_sc_hs__nand2_1_29/B prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_41/Y
+ prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_53/a_132_392# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_45/a_206_368#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_15/a_437_503# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_37/a_651_503#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_39/a_544_485# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_53/a_735_102#
+ prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_45/a_52_123# prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_1/B
+ prbs_generator_syn_31/sky130_fd_sc_hs__nand2_2_3/B prbs_generator_syn_31/sky130_fd_sc_hs__clkbuf_16_1/A
+ prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_21/X prbs_generator_syn_31/sky130_fd_sc_hs__nand2_1_25/B
+ prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_39/a_376_368# prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_63/X
+ prbs_generator_syn_31/m3_13600_3481# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_69/a_1178_124#
+ prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_21/a_138_385# prbs_generator_syn_31/sky130_fd_sc_hs__nor2b_1_8/Y
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_19/a_1178_124# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_49/a_27_74#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_45/a_437_503# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_27/a_651_503#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_71/a_1141_508# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_65/a_651_503#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_29/a_544_485# prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_3/a_138_385#
+ prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_55/X prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_43/a_735_102#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_41/a_1034_424# prbs_generator_syn_31/sky130_fd_sc_hs__nand2_1_9/B
+ prbs_generator_syn_31/sky130_fd_sc_hs__nor2b_1_9/Y prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_59/a_1034_424#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_39/a_1141_508# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_33/a_1226_296#
+ prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_49/a_52_123# prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_47/Y
+ prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_43/Y prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_4/a_651_503#
+ prbs_generator_syn_31/sky130_fd_sc_hs__nand2_1_49/B prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_19/A
+ prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_11/a_138_385# prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_5/X
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_63/a_206_368# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_17/a_651_503#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_19/a_544_485# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_55/a_651_503#
+ prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_9/Y prbs_generator_syn_31/sky130_fd_sc_hs__nand2_1_17/B
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_57/a_544_485# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_67/a_696_458#
+ prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_35/X prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_19/a_27_74#
+ prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_45/a_222_392# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_32/a_1226_296#
+ prbs_generator_syn_31/sky130_fd_sc_hs__nand2_1_43/B prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_25/A
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_1/a_206_368# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_49/a_1226_296#
+ prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_1/a_112_119# prbs_generator_syn_31/sky130_fd_sc_hs__or2_1_1/X
+ prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_59/a_376_368# prbs_generator_syn_31/sky130_fd_sc_hs__nand2_1_19/B
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_5/a_696_458# prbs_generator_syn_31/sky130_fd_sc_hs__nor2b_1_1/Y
+ prbs_generator_syn_31/sky130_fd_sc_hs__nor2b_1_5/a_278_368# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_17/a_1178_124#
+ prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_39/X prbs_generator_syn_31/m3_13600_5433#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_63/a_437_503# prbs_generator_syn_31/sky130_fd_sc_hs__nand2_2_5/B
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_23/a_735_102# prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_53/A
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_61/a_735_102# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_57/a_1034_424#
+ prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_63/B prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_37/a_1141_508#
+ prbs_generator_syn_31/sky130_fd_sc_hs__nand2_1_47/B prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_29/X
+ prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_65/Y prbs_generator_syn_31/m3_13600_4701#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_1/a_437_503# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_67/a_1178_124#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_9/a_735_102# prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_13/a_132_392#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_15/a_1178_124# prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_15/A
+ prbs_generator_syn_31/sky130_fd_sc_hs__nand2_1_1/B prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_43/B
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_35/a_651_503# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_8/D
+ prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_29/A prbs_generator_syn_31/sky130_fd_sc_hs__nand2_1_7/B
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_13/a_735_102# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_47/a_696_458#
+ prbs_generator_syn_31/sky130_fd_sc_hs__nand2_1_31/B prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_51/a_735_102#
+ prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_59/X prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_35/a_1141_508#
+ prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_25/a_222_392# prbs_generator_syn_31/sky130_fd_sc_hs__sdlclkp_2_1/a_288_48#
+ prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_55/B prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_17/B
+ prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_43/A prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_7/A
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_65/a_1178_124# prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_59/Y
+ prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_41/X prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_21/a_230_79#
+ prbs_generator_syn_31/sky130_fd_sc_hs__nand2_1_57/a_117_74# prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_1/a_222_392#
+ prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_19/B prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_35/a_293_74#
+ prbs_generator_syn_31/sky130_fd_sc_hs__nand2_1_23/a_117_74# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_73/a_206_368#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_25/a_651_503# prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_1/a_138_385#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_37/a_696_458# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_67/a_544_485#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_43/a_27_74# prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_9/X
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_55/a_1034_424# prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_39/a_112_119#
+ prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_15/a_222_392# prbs_generator_syn_31/sky130_fd_sc_hs__conb_1_1/HI
+ prbs_generator_syn_31/sky130_fd_sc_hs__nand2_1_23/B prbs_generator_syn_31/sky130_fd_sc_hs__nand2_1_53/B
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_9/a_1178_124# prbs_generator_syn_31/sky130_fd_sc_hs__nor2b_1_4/A
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_47/a_1226_296# prbs_generator_syn_31/m3_13600_11045#
+ prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_17/X prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_29/a_376_368#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_5/a_544_485# prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_3/X
+ prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_31/a_132_392# prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_61/A
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_15/a_651_503# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_73/a_437_503#
+ prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_25/a_230_79# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_27/a_696_458#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_65/a_696_458# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_33/a_735_102#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_71/a_735_102# prbs_generator_syn_31/m3_13600_7263#
+ prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_43/a_222_392# prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_50/Y
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_8/a_1178_124# prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_53/B
+ prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_19/a_376_368# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_63/a_1178_124#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_4/a_696_458# prbs_generator_syn_31/sky130_fd_sc_hs__nor2b_1_4/a_278_368#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_13/a_1178_124# prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_61/a_132_392#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_53/a_206_368# prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_21/a_52_123#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_45/a_651_503# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_17/a_696_458#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_47/a_544_485# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_55/a_696_458#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_21/a_735_102# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_37/a_27_74#
+ prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_61/B prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_61/X
+ prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_59/a_112_119# prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_31/A
+ prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_33/a_222_392# prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_29/a_230_79#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_45/a_1226_296# prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_9/a_132_392#
+ prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_5/A prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_57/Y
+ prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_31/X prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_51/a_27_74#
+ prbs_generator_syn_31/sky130_fd_sc_hs__nor2b_1_8/a_27_112# prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_47/a_376_368#
+ prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_53/a_293_74# prbs_generator_syn_31/sky130_fd_sc_hs__nand2_1_43/a_117_74#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_8/a_735_102# prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_21/a_293_74#
+ prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_39/a_138_385# prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_63/Y
+ prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_51/a_132_392# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_43/a_206_368#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_53/a_437_503# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_37/a_544_485#
+ prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_57/X prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_53/a_1034_424#
+ prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_25/a_52_123# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_33/a_1141_508#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_63/Q prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_23/a_222_392#
+ prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_63/a_222_392# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_7/a_1178_124#
+ prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_53/X prbs_generator_syn_31/sky130_fd_sc_hs__nand2_2_5/Y
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_61/a_1178_124# prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_1/a_230_79#
+ prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_43/a_230_79# prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_11/a_230_79#
+ prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_41/a_132_392# prbs_generator_syn_31/sky130_fd_sc_hs__nand2_1_13/a_117_74#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_43/a_437_503# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_27/a_544_485#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_63/a_651_503# prbs_generator_syn_31/sky130_fd_sc_hs__nand2_1_7/a_117_74#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_35/a_696_458# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_65/a_544_485#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_51/a_1034_424# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_41/a_735_102#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_32/a_1141_508# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_49/a_1141_508#
+ prbs_generator_syn_31/sky130_fd_sc_hs__nand2_1_55/B prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_53/a_222_392#
+ prbs_generator_syn_31/sky130_fd_sc_hs__sdlclkp_2_1/a_114_112# prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_9/a_293_74#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_43/a_1226_296# prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_29/a_52_123#
+ prbs_generator_syn_31/sky130_fd_sc_hs__nand2_1_37/B prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_1/a_651_503#
+ prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_27/a_376_368# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_4/a_544_485#
+ prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_67/a_376_368# prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_27/X
+ prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_1/X prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_59/a_138_385#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_29/a_1178_124# prbs_generator_syn_31/m3_13600_2871#
+ prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_5/a_230_79# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_23/a_206_368#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_61/a_206_368# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_17/a_544_485#
+ prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_15/a_230_79# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_25/a_696_458#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_55/a_544_485# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_32/a_735_102#
+ prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_29/a_293_74# prbs_generator_syn_31/sky130_fd_sc_hs__nand2_1_17/a_117_74#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_69/a_1034_424# prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_29/a_112_119#
+ prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_37/X prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_31/B
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_19/a_1034_424# prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_33/A
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_9/a_206_368# prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_57/a_376_368#
+ prbs_generator_syn_31/sky130_fd_sc_hs__sdlclkp_2_1/a_706_317# prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_11/B
+ prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_1/a_52_123# prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_39/B
+ prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_21/a_132_392# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_13/a_206_368#
+ prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_43/a_52_123# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_51/a_206_368#
+ prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_47/X prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_23/a_437_503#
+ prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_11/a_52_123# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_61/a_437_503#
+ prbs_generator_syn_31/sky130_fd_sc_hs__nor2b_1_7/Y prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_51/A
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_15/a_696_458# prbs_generator_syn_31/sky130_fd_sc_hs__nor2b_1_5/Y
+ prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_9/a_230_79# prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_25/X
+ prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_19/a_112_119# prbs_generator_syn_31/sky130_fd_sc_hs__nand2_1_45/B
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_5/a_1178_124# prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_19/a_230_79#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_41/a_1226_296# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_59/a_1226_296#
+ prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_63/a_230_79# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_51/Q
+ prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_7/a_132_392# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_9/a_437_503#
+ prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_46/a_376_368# prbs_generator_syn_31/sky130_fd_sc_hs__nand2_1_33/a_117_74#
+ prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_11/a_293_74# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_27/a_1178_124#
+ prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_11/a_132_392# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_13/a_437_503#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_51/a_437_503# prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_5/a_52_123#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_35/a_544_485# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_73/a_651_503#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_45/a_696_458# prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_15/a_52_123#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_47/a_1141_508# prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_47/a_112_119#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_4/a_1178_124# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_17/a_1034_424#
+ prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_23/B prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_37/a_376_368#
+ prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_15/B prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_7/Y
+ prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_29/a_138_385# prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_33/a_230_79#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_25/a_1178_124# prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_47/a_293_74#
+ prbs_generator_syn_31/sky130_fd_sc_hs__nand2_1_37/a_117_74# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_33/a_206_368#
+ prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_15/a_293_74# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_71/a_206_368#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_25/a_544_485# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_67/a_1034_424#
+ prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_13/a_222_392# prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_9/a_52_123#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_15/a_1034_424# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_57/a_1226_296#
+ prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_19/a_52_123# prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_23/X
+ prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_63/a_52_123# prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_19/a_138_385#
+ prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_9/a_376_368# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_21/a_206_368#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_33/a_437_503# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_71/a_437_503#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_53/a_651_503# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_15/a_544_485#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_63/a_696_458# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_65/a_1034_424#
+ prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_19/a_293_74# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_45/a_1141_508#
+ prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_27/a_112_119# prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_67/a_112_119#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_1/a_1178_124# prbs_generator_syn_31/sky130_fd_sc_hs__conb_1_1/a_21_290#
+ prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_63/a_293_74# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_8/a_206_368#
+ prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_17/a_376_368# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_63/a_27_74#
+ prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_21/A prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_55/a_376_368#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_1/a_696_458# prbs_generator_syn_31/sky130_fd_sc_hs__nor2b_1_1/a_278_368#
+ prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_47/a_138_385# prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_33/a_52_123#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_9/a_1034_424# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_21/a_437_503#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_1/a_27_74# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_43/a_651_503#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_1/Q prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_45/a_544_485#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_69/a_735_102# prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_57/a_112_119#
+ prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_31/a_222_392# prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_13/A
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_55/a_1226_296# prbs_generator_syn_31/sky130_fd_sc_hs__nand2_2_5/a_27_74#
+ prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_53/a_230_79# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_8/a_437_503#
+ prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_67/a_293_74# prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_33/a_293_74#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_7/a_735_102# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_23/a_1178_124#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_41/a_206_368# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_8/a_1034_424#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_63/a_1034_424# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_59/a_735_102#
+ prbs_generator_syn_31/sky130_fd_sc_hs__nand2_1_5/B prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_43/a_1141_508#
+ prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_46/a_112_119# prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_61/a_222_392#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_13/a_1034_424# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_73/a_1178_124#
+ prbs_generator_syn_31/sky130_fd_sc_hs__nand2_1_27/B prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_13/B
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_57/a_27_74# prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_57/a_230_79#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_21/a_1178_124# prbs_generator_syn_31/sky130_fd_sc_hs__nor2b_1_1/a_27_112#
+ prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_27/a_138_385# prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_23/a_230_79#
+ prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_67/a_138_385# prbs_generator_syn_31/sky130_fd_sc_hs__nand2_1_41/B
+ prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_9/a_222_392# prbs_generator_syn_31/sky130_fd_sc_hs__nand2_1_27/a_117_74#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_32/a_206_368# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_23/a_651_503#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_41/a_437_503# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_73/a_27_74#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_61/a_651_503# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_63/a_544_485#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_49/a_735_102# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_73/a_696_458#
+ prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_37/a_112_119# prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_51/a_222_392#
+ prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_43/X prbs_generator_syn_31/sky130_fd_sc_hs__nand2_2_1/B
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_9/a_651_503# prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_53/a_52_123#
+ prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_49/X prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_25/a_376_368#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_1/a_544_485# prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_65/a_376_368#
+ prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_57/a_138_385# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_27/a_27_74#
+ prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_39/a_132_392# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_7/a_1034_424#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_13/a_651_503# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_32/a_437_503#
+ prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_27/a_230_79# prbs_generator_syn_31/m3_13600_12265#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_51/a_651_503# prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_59/B
+ prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_47/A prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_61/a_1034_424#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_41/a_1141_508# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_59/a_1141_508#
+ prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_41/a_222_392# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_53/a_1226_296#
+ prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_3/A prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_71/a_1178_124#
+ prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_9/a_112_119# prbs_generator_syn_31/sky130_fd_sc_hs__nand2_1_3/a_117_74#
+ prbs_generator_syn_31/m3_13600_8483# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_39/a_1178_124#
+ prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_57/a_52_123# prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_46/a_138_385#
+ prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_23/a_52_123# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_67/a_27_74#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_53/a_696_458# prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_17/a_112_119#
+ prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_11/A prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_55/a_112_119#
+ prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_1/A prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_51/a_1226_296#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_29/a_1034_424# prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_59/A
+ prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_23/A prbs_generator_syn_31/sky130_fd_sc_hs__nand2_1_39/B
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_5/a_27_74# prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_57/a_293_74#
+ prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_37/a_138_385# prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_59/a_132_392#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_33/a_651_503# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_71/a_651_503#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_43/a_696_458# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_73/a_544_485#
+ prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_27/a_52_123# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_57/a_1141_508#
+ prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_21/a_222_392# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_35/a_27_74#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_69/a_1226_296# prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_37/B
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_19/a_1226_296# prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_35/a_376_368#
+ prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_47/a_230_79# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_37/a_1178_124#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_5/a_1034_424# prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_49/a_132_392#
+ prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_7/a_222_392# prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_27/a_293_74#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_21/a_651_503# prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_9/a_138_385#
+ prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_11/a_222_392# prbs_generator_syn_31/m3_13600_14095#
+ prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_50/A prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_27/a_1034_424#
+ prbs_generator_syn_31/sky130_fd_sc_hs__nand2_1_13/B prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_8/a_651_503#
+ prbs_generator_syn_31/m3_13600_9703# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_35/a_1178_124#
+ prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_17/a_138_385# prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_55/a_138_385#
+ prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_7/a_230_79# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_4/a_1034_424#
+ prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_7/a_376_368# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_69/a_206_368#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_23/a_696_458# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_53/a_544_485#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_39/a_735_102# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_61/a_696_458#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_55/a_1141_508# prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_25/a_112_119#
+ prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_65/a_112_119# prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_43/a_293_74#
+ prbs_generator_syn_31/sky130_fd_sc_hs__nand2_1_57/B prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_25/a_1034_424#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_7/a_206_368# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_17/a_1226_296#
+ prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_15/a_376_368# prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_53/a_376_368#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_9/a_696_458# prbs_generator_syn_31/m3_13600_431#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_45/a_27_74# prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_47/a_52_123#
+ prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_29/a_132_392# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_59/a_206_368#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_69/a_437_503# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_41/a_651_503#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_43/a_544_485# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_13/a_696_458#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_29/a_735_102# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_51/a_696_458#
+ prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_61/Y prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_67/a_1226_296#
+ prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_5/a_132_392# prbs_generator_syn_31/sky130_fd_sc_hs__and2b_2_1/a_198_48#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_7/a_437_503# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_15/a_1226_296#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_69/a_27_74# prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_46/a_293_74#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_1/a_1034_424# prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_19/a_132_392#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_49/a_206_368# prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_7/a_52_123#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_59/a_437_503# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_32/a_651_503#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_7/a_27_74# prbs_generator_syn_31/sky130_fd_sc_hs__nand2_2_1/a_27_74#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_19/a_735_102# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_57/a_735_102#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_65/a_1226_296# prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_37/A
+ prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_33/a_376_368# prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_37/a_230_79#
+ prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_25/a_138_385# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_39/a_27_74#
+ prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_65/a_138_385# prbs_generator_syn_31/sky130_fd_sc_hs__nor2b_1_9/a_278_368#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_49/a_437_503# prbs_generator_syn_31/sky130_fd_sc_hs__and2b_2_1/a_505_74#
+ prbs_generator_syn_31/sky130_fd_sc_hs__nand2_1_51/a_117_74# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_23/a_544_485#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_33/a_696_458# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_61/a_544_485#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_9/a_1226_296# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_53/a_1141_508#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_71/a_696_458# prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_35/a_112_119#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_23/a_1034_424# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_9/a_544_485#
+ prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_63/a_376_368# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_33/a_1178_124#
+ prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_5/a_376_368# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_13/a_544_485#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_73/a_1034_424# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_21/a_696_458#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_51/a_544_485# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_8/a_1226_296#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_51/a_1141_508# prbs_generator_syn_31/sky130_fd_sc_hs__nand2_1_55/a_117_74#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_21/a_1034_424# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_63/a_1226_296#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_23/a_27_74# prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_7/a_112_119#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_13/a_1226_296# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_8/a_696_458#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_32/a_1178_124# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_49/a_1178_124#
+ prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_37/a_52_123# prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_27/a_132_392#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_71/Q prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_67/a_735_102#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_69/a_1141_508# prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_15/a_112_119#
+ prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_53/a_112_119# prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_39/a_222_392#
+ prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_55/a_230_79# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_19/a_1141_508#
+ prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_37/a_293_74# prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_43/a_376_368#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_5/a_735_102# prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_35/a_138_385#
+ prbs_generator_syn_31/sky130_fd_sc_hs__sdlclkp_2_1/a_114_424# prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_57/a_132_392#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_71/a_1034_424# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_7/a_1226_296#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_33/a_544_485# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_41/a_696_458#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_71/a_544_485# prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_21/B
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_61/a_1226_296# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_39/a_1034_424#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_17/a_27_74# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_9/a_27_74#
+ prbs_generator_syn_31/sky130_fd_sc_hs__nor2b_1_5/a_27_112# prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_47/a_132_392#
+ prbs_generator_syn_31/sky130_fd_sc_hs__nor2b_1_8/a_278_368# prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_9/B
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_39/a_206_368# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_33/a_27_74#
+ prbs_generator_syn_31/sky130_fd_sc_hs__nand2_1_41/a_117_74# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_69/a_651_503#
+ prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_51/a_293_74# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_21/a_544_485#
+ prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_7/a_138_385# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_32/a_696_458#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_47/a_735_102# prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_33/a_112_119#
+ prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_59/a_222_392# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_17/a_1141_508#
+ prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_55/a_52_123# prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_3/a_293_74#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_7/a_651_503# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_29/a_1226_296#
+ prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_23/a_376_368# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_8/a_544_485#
+ prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_47/B prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_47/a_1178_124#
+ prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_15/a_138_385# prbs_generator_syn_31/sky130_fd_sc_hs__sdlclkp_2_1/a_1195_374#
+ prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_53/a_138_385# prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_37/a_132_392#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_29/a_206_368# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_39/a_437_503#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_59/a_651_503# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_37/a_735_102#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_67/a_1141_508# prbs_generator_syn_31/sky130_fd_sc_hs__and2b_2_1/a_27_74#
+ prbs_generator_syn_31/sky130_fd_sc_hs__conb_1_1/a_165_290# prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_55/a_293_74#
+ prbs_generator_syn_31/sky130_fd_sc_hs__nand2_1_45/a_117_74# prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_63/a_112_119#
+ prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_49/a_222_392# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_37/a_1034_424#
+ prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_23/a_293_74# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_15/a_1141_508#
+ prbs_generator_syn_31/sky130_fd_sc_hs__nand2_1_5/a_117_74# prbs_generator_syn_31/m3_13600_13485#
+ prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_5/a_112_119# prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_13/a_376_368#
+ prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_51/a_376_368# prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_7/a_293_74#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_19/a_206_368# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_57/a_206_368#
+ prbs_generator_syn_31/sky130_fd_sc_hs__sdlclkp_2_1/a_318_74# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_29/a_437_503#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_49/a_651_503# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_25/a_27_74#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_5/a_1226_296# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_41/a_544_485#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_27/a_735_102# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_65/a_1141_508#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_65/a_735_102# prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_3/a_230_79#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_35/a_1034_424# prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_13/a_230_79#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_41/a_27_74# prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_3/a_132_392#
+ prbs_generator_syn_31/sky130_fd_sc_hs__nand2_1_49/a_117_74# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_27/a_1226_296#
+ prbs_generator_syn_31/sky130_fd_sc_hs__nand2_1_15/a_117_74# prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_41/a_376_368#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_45/a_1178_124# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_4/a_735_102#
+ prbs_generator_syn_31/sky130_fd_sc_hs__nand2_1_9/a_117_74# prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_33/a_138_385#
+ prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_17/a_132_392# prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_55/a_132_392#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_9/a_1141_508# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_19/a_437_503#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_57/a_437_503# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_4/a_1226_296#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_32/a_544_485# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_17/a_735_102#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_55/a_735_102# prbs_generator_syn_31/m3_13600_2261#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_65/a_27_74# prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_29/a_222_392#
+ prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_43/a_112_119# prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_19/X
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_25/a_1226_296# prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_31/a_376_368#
+ prbs_generator_syn_31/sky130_fd_sc_hs__or2_1_1/a_63_368# prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_17/a_230_79#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_4/a_27_74# prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_61/a_230_79#
+ prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_63/a_138_385# prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_5/a_222_392#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_8/a_1141_508# prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_41/a_293_74#
+ prbs_generator_syn_31/sky130_fd_sc_hs__nand2_1_31/a_117_74# prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_5/a_138_385#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_63/a_1141_508# prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_19/a_222_392#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_13/a_1141_508# prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_3/a_52_123#
+ prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_13/a_52_123# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_43/a_1178_124#
+ prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_61/a_376_368# prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_35/a_132_392#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_67/a_206_368# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_1/a_1226_296#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_69/a_696_458# prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_31/a_230_79#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_35/a_735_102# prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_23/a_112_119#
+ prbs_generator_syn_31/sky130_fd_sc_hs__nand2_1_35/a_117_74# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_59/a_27_74#
+ prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_13/a_293_74# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_5/a_206_368#
+ prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_50/a_376_368# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_7/a_696_458#
+ prbs_generator_syn_31/sky130_fd_sc_hs__nor2b_1_7/a_278_368# prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_17/a_52_123#
+ prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_43/a_138_385# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_7/a_1141_508#
+ prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_61/a_52_123# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_67/a_437_503#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_61/a_1141_508# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_25/a_735_102#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_59/a_696_458# prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_13/a_112_119#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_33/a_1034_424# prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_51/a_112_119#
+ prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_35/a_230_79# prbs_generator_syn_31/m3_13600_4091#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_23/a_1226_296# prbs_generator_syn_31/sky130_fd_sc_hs__nand2_1_39/a_117_74#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_29/a_27_74# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_5/a_437_503#
+ prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_17/a_293_74# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_41/a_1178_124#
+ prbs_generator_syn_31/sky130_fd_sc_hs__or2_1_1/a_152_368# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_59/a_1178_124#
+ prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_61/a_293_74# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_47/a_206_368#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_39/a_651_503# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_49/a_696_458#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_15/a_735_102# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_32/a_1034_424#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_73/a_1226_296# prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_27/a_222_392#
+ prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_41/a_112_119# prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_31/a_52_123#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_49/a_1034_424# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_29/a_1141_508#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_21/a_1226_296# prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_39/a_230_79#
+ prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_23/a_138_385# prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_51/a_230_79#
+ prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_45/a_132_392# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_37/a_206_368#
+ prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_65/a_293_74# prbs_generator_syn_31/sky130_fd_sc_hs__nand2_1_53/a_117_74#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_47/a_437_503# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_29/a_651_503#
+ prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_31/a_293_74# prbs_generator_syn_31/sky130_fd_sc_hs__nand2_1_21/a_117_74#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_69/a_544_485# prbs_generator_syn_31/sky130_fd_sc_hs__clkbuf_16_1/a_114_74#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_45/a_735_102# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_13/a_27_74#
+ prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_31/a_112_119# prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_57/a_222_392#
+ prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_35/a_52_123# prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_21/a_376_368#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_7/a_544_485# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_57/a_1178_124#
+ prbs_generator_syn_31/m3_13600_6043# prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_13/a_138_385#
+ prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_51/a_138_385# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_5/a_1141_508#
+ prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_3/a_376_368# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_27/a_206_368#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_65/a_206_368# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_37/a_437_503#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_19/a_651_503# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_57/a_651_503#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_59/a_544_485# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_71/a_1226_296#
+ prbs_generator_syn_31/sky130_fd_sc_hs__nand2_1_25/a_117_74# prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_61/a_112_119#
+ prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_47/a_222_392# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_27/a_1141_508#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_53/a_27_74# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_4/a_206_368#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_39/a_1226_296# prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_11/a_376_368#
+ prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_39/a_52_123# prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_41/a_138_385#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_4/a_1141_508# prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_25/a_132_392#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_17/a_206_368# prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_41/A
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_55/a_206_368# prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_51/a_52_123#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_27/a_437_503# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_65/a_437_503#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_49/a_544_485# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_63/a_735_102#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_47/a_1034_424# prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_50/a_112_119#
+ prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_37/a_222_392# prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_59/a_230_79#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_25/a_1141_508# prbs_generator_syn_31/sky130_fd_sc_hs__nor2b_1_4/a_27_112#
+ prbs_generator_syn_31/sky130_fd_sc_hs__sdlclkp_2_1/a_685_81# prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_1/a_132_392#
+ prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_39/a_293_74# prbs_generator_syn_31/sky130_fd_sc_hs__nand2_1_29/a_117_74#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_4/a_437_503# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_55/a_1178_124#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_21/a_27_74# prbs_generator_syn_31/m3_13600_12875#
+ prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_50/a_293_74# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_1/a_735_102#
+ prbs_generator_syn_31/sky130_fd_sc_hs__xnor2_1_31/a_138_385# prbs_generator_syn_31/sky130_fd_sc_hs__a22o_1_15/a_132_392#
+ prbs_generator_syn_31/sky130_fd_sc_hs__nand2_1_1/a_117_74# prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_17/a_437_503#
+ prbs_generator_syn_31/sky130_fd_sc_hs__dfxtp_4_55/a_437_503# prbs_generator_syn
Xsky130_fd_sc_hs__buf_2_140 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__buf_2_37/X sky130_fd_sc_hs__buf_2_141/X
+ sky130_fd_sc_hs__buf_2_141/a_21_260# sky130_fd_sc_hs__buf_2
Xsky130_fd_sc_hs__buf_2_151 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__buf_2_151/A sky130_fd_sc_hs__buf_2_151/X
+ sky130_fd_sc_hs__buf_2_151/a_21_260# sky130_fd_sc_hs__buf_2
Xsky130_fd_sc_hs__buf_2_162 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__buf_2_67/X sky130_fd_sc_hs__buf_2_163/X
+ sky130_fd_sc_hs__buf_2_163/a_21_260# sky130_fd_sc_hs__buf_2
Xsky130_fd_sc_hs__einvp_2_30 DVSS: DVDD: DVDD: DVSS: dout_n sky130_fd_sc_hs__buf_8_1/A
+ sky130_fd_sc_hs__dlrtp_1_27/Q sky130_fd_sc_hs__einvp_2_31/a_263_323# sky130_fd_sc_hs__einvp_2_31/a_36_74#
+ sky130_fd_sc_hs__einvp_2_31/a_27_368# sky130_fd_sc_hs__einvp_2
Xsky130_fd_sc_hs__einvp_2_41 DVSS: DVDD: DVDD: DVSS: dout_n sky130_fd_sc_hs__buf_8_1/A
+ sky130_fd_sc_hs__dlrtp_1_35/Q sky130_fd_sc_hs__einvp_2_41/a_263_323# sky130_fd_sc_hs__einvp_2_41/a_36_74#
+ sky130_fd_sc_hs__einvp_2_41/a_27_368# sky130_fd_sc_hs__einvp_2
Xsky130_fd_sc_hs__einvp_2_52 DVSS: DVDD: DVDD: DVSS: dout_p sky130_fd_sc_hs__inv_4_9/Y
+ sky130_fd_sc_hs__dlrtp_1_45/Q sky130_fd_sc_hs__einvp_2_53/a_263_323# sky130_fd_sc_hs__einvp_2_53/a_36_74#
+ sky130_fd_sc_hs__einvp_2_53/a_27_368# sky130_fd_sc_hs__einvp_2
Xsky130_fd_sc_hs__clkbuf_4_8 DVSS: DVDD: DVDD: DVSS: pi1_con[0] sky130_fd_sc_hs__clkbuf_8_5/A
+ sky130_fd_sc_hs__clkbuf_4_9/a_83_270# sky130_fd_sc_hs__clkbuf_4
Xsky130_fd_sc_hs__einvp_2_63 DVSS: DVDD: DVDD: DVSS: dout_p sky130_fd_sc_hs__einvp_2_65/A
+ sky130_fd_sc_hs__dlrtp_1_49/Q sky130_fd_sc_hs__einvp_2_63/a_263_323# sky130_fd_sc_hs__einvp_2_63/a_36_74#
+ sky130_fd_sc_hs__einvp_2_63/a_27_368# sky130_fd_sc_hs__einvp_2
Xsky130_fd_sc_hs__einvp_2_74 DVSS: DVDD: DVDD: DVSS: dout_p sky130_fd_sc_hs__einvp_2_99/A
+ sky130_fd_sc_hs__einvp_2_75/TE sky130_fd_sc_hs__einvp_2_75/a_263_323# sky130_fd_sc_hs__einvp_2_75/a_36_74#
+ sky130_fd_sc_hs__einvp_2_75/a_27_368# sky130_fd_sc_hs__einvp_2
Xsky130_fd_sc_hs__einvp_2_85 DVSS: DVDD: DVDD: DVSS: dout_p sky130_fd_sc_hs__einvp_2_97/A
+ sky130_fd_sc_hs__dlrtp_1_69/Q sky130_fd_sc_hs__einvp_2_85/a_263_323# sky130_fd_sc_hs__einvp_2_85/a_36_74#
+ sky130_fd_sc_hs__einvp_2_85/a_27_368# sky130_fd_sc_hs__einvp_2
Xsky130_fd_sc_hs__einvp_2_96 DVSS: DVDD: DVDD: DVSS: dout_p sky130_fd_sc_hs__einvp_2_97/A
+ sky130_fd_sc_hs__dlrtp_1_79/Q sky130_fd_sc_hs__einvp_2_97/a_263_323# sky130_fd_sc_hs__einvp_2_97/a_36_74#
+ sky130_fd_sc_hs__einvp_2_97/a_27_368# sky130_fd_sc_hs__einvp_2
Xsky130_fd_sc_hs__or2b_2_0 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__or2b_2_1/X sky130_fd_sc_hs__nor2_4_1/Y
+ sky130_fd_sc_hs__or2b_2_1/A sky130_fd_sc_hs__or2b_2_1/a_470_368# sky130_fd_sc_hs__or2b_2_1/a_27_368#
+ sky130_fd_sc_hs__or2b_2_1/a_187_48# sky130_fd_sc_hs__or2b_2
Xsky130_fd_sc_hs__clkinv_4_8 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__nor2_4_1/B sky130_fd_sc_hs__o21ai_4_1/A1
+ sky130_fd_sc_hs__clkinv_4
Xsky130_fd_sc_hs__conb_1_40 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__conb_1_41/LO
+ sky130_fd_sc_hs__conb_1_41/HI sky130_fd_sc_hs__conb_1_41/a_165_290# sky130_fd_sc_hs__conb_1_41/a_21_290#
+ sky130_fd_sc_hs__conb_1
Xsky130_fd_sc_hs__conb_1_51 DVSS: DVDD: DVDD: DVSS: prbs_generator_syn_7/eqn[9] sky130_fd_sc_hs__conb_1_51/HI
+ sky130_fd_sc_hs__conb_1_51/a_165_290# sky130_fd_sc_hs__conb_1_51/a_21_290# sky130_fd_sc_hs__conb_1
Xsky130_fd_sc_hs__conb_1_62 DVSS: DVDD: DVDD: DVSS: prbs_generator_syn_7/eqn[0] sky130_fd_sc_hs__conb_1_63/HI
+ sky130_fd_sc_hs__conb_1_63/a_165_290# sky130_fd_sc_hs__conb_1_63/a_21_290# sky130_fd_sc_hs__conb_1
Xsky130_fd_sc_hs__conb_1_73 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__conb_1_73/LO
+ sky130_fd_sc_hs__conb_1_73/HI sky130_fd_sc_hs__conb_1_73/a_165_290# sky130_fd_sc_hs__conb_1_73/a_21_290#
+ sky130_fd_sc_hs__conb_1
Xsky130_fd_sc_hs__conb_1_84 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__conb_1_85/LO
+ sky130_fd_sc_hs__conb_1_85/HI sky130_fd_sc_hs__conb_1_85/a_165_290# sky130_fd_sc_hs__conb_1_85/a_21_290#
+ sky130_fd_sc_hs__conb_1
Xsky130_fd_sc_hs__conb_1_95 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__conb_1_95/LO
+ sky130_fd_sc_hs__conb_1_95/HI sky130_fd_sc_hs__conb_1_95/a_165_290# sky130_fd_sc_hs__conb_1_95/a_21_290#
+ sky130_fd_sc_hs__conb_1
Xsky130_fd_sc_hs__inv_4_80 DVSS: DVDD: DVDD: DVSS: hr_16t4_mux_top_3/din[8] hr_16t4_mux_top_1/din[8]
+ sky130_fd_sc_hs__inv_4
Xsky130_fd_sc_hs__dlrtp_1_107 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__einvp_2_27/TE
+ sky130_fd_sc_hs__dlrtp_1_9/GATE sky130_fd_sc_hs__conb_1_133/HI sky130_fd_sc_hs__dlrtp_1_107/D
+ sky130_fd_sc_hs__dlrtp_1_107/a_216_424# sky130_fd_sc_hs__dlrtp_1_107/a_759_508#
+ sky130_fd_sc_hs__dlrtp_1_107/a_565_74# sky130_fd_sc_hs__dlrtp_1_107/a_27_424# sky130_fd_sc_hs__dlrtp_1_107/a_1045_74#
+ sky130_fd_sc_hs__dlrtp_1_107/a_643_74# sky130_fd_sc_hs__dlrtp_1_107/a_817_48# sky130_fd_sc_hs__dlrtp_1_107/a_568_392#
+ sky130_fd_sc_hs__dlrtp_1_107/a_363_74# sky130_fd_sc_hs__dlrtp_1_107/a_769_74# sky130_fd_sc_hs__dlrtp_1
Xsky130_fd_sc_hs__dlrtp_1_118 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__dlrtp_1_119/Q
+ sky130_fd_sc_hs__dlrtp_1_9/GATE sky130_fd_sc_hs__conb_1_131/HI sky130_fd_sc_hs__buf_2_117/X
+ sky130_fd_sc_hs__dlrtp_1_119/a_216_424# sky130_fd_sc_hs__dlrtp_1_119/a_759_508#
+ sky130_fd_sc_hs__dlrtp_1_119/a_565_74# sky130_fd_sc_hs__dlrtp_1_119/a_27_424# sky130_fd_sc_hs__dlrtp_1_119/a_1045_74#
+ sky130_fd_sc_hs__dlrtp_1_119/a_643_74# sky130_fd_sc_hs__dlrtp_1_119/a_817_48# sky130_fd_sc_hs__dlrtp_1_119/a_568_392#
+ sky130_fd_sc_hs__dlrtp_1_119/a_363_74# sky130_fd_sc_hs__dlrtp_1_119/a_769_74# sky130_fd_sc_hs__dlrtp_1
Xsky130_fd_sc_hs__dlrtp_1_129 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__buf_2_17/A
+ sky130_fd_sc_hs__clkbuf_2_3/A sky130_fd_sc_hs__conb_1_121/HI sky130_fd_sc_hs__buf_2_137/X
+ sky130_fd_sc_hs__dlrtp_1_129/a_216_424# sky130_fd_sc_hs__dlrtp_1_129/a_759_508#
+ sky130_fd_sc_hs__dlrtp_1_129/a_565_74# sky130_fd_sc_hs__dlrtp_1_129/a_27_424# sky130_fd_sc_hs__dlrtp_1_129/a_1045_74#
+ sky130_fd_sc_hs__dlrtp_1_129/a_643_74# sky130_fd_sc_hs__dlrtp_1_129/a_817_48# sky130_fd_sc_hs__dlrtp_1_129/a_568_392#
+ sky130_fd_sc_hs__dlrtp_1_129/a_363_74# sky130_fd_sc_hs__dlrtp_1_129/a_769_74# sky130_fd_sc_hs__dlrtp_1
Xsky130_fd_sc_hs__dlrtp_1_20 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__dlrtp_1_21/Q
+ sky130_fd_sc_hs__clkbuf_2_3/X sky130_fd_sc_hs__conb_1_119/HI sky130_fd_sc_hs__dlrtp_1_21/D
+ sky130_fd_sc_hs__dlrtp_1_21/a_216_424# sky130_fd_sc_hs__dlrtp_1_21/a_759_508# sky130_fd_sc_hs__dlrtp_1_21/a_565_74#
+ sky130_fd_sc_hs__dlrtp_1_21/a_27_424# sky130_fd_sc_hs__dlrtp_1_21/a_1045_74# sky130_fd_sc_hs__dlrtp_1_21/a_643_74#
+ sky130_fd_sc_hs__dlrtp_1_21/a_817_48# sky130_fd_sc_hs__dlrtp_1_21/a_568_392# sky130_fd_sc_hs__dlrtp_1_21/a_363_74#
+ sky130_fd_sc_hs__dlrtp_1_21/a_769_74# sky130_fd_sc_hs__dlrtp_1
Xsky130_fd_sc_hs__dlrtp_1_31 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__dlrtp_1_31/Q
+ sky130_fd_sc_hs__clkbuf_2_3/A sky130_fd_sc_hs__conb_1_121/HI sky130_fd_sc_hs__buf_2_133/X
+ sky130_fd_sc_hs__dlrtp_1_31/a_216_424# sky130_fd_sc_hs__dlrtp_1_31/a_759_508# sky130_fd_sc_hs__dlrtp_1_31/a_565_74#
+ sky130_fd_sc_hs__dlrtp_1_31/a_27_424# sky130_fd_sc_hs__dlrtp_1_31/a_1045_74# sky130_fd_sc_hs__dlrtp_1_31/a_643_74#
+ sky130_fd_sc_hs__dlrtp_1_31/a_817_48# sky130_fd_sc_hs__dlrtp_1_31/a_568_392# sky130_fd_sc_hs__dlrtp_1_31/a_363_74#
+ sky130_fd_sc_hs__dlrtp_1_31/a_769_74# sky130_fd_sc_hs__dlrtp_1
Xsky130_fd_sc_hs__dlrtp_1_42 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__dlrtp_1_43/Q
+ sky130_fd_sc_hs__clkbuf_16_53/A sky130_fd_sc_hs__conb_1_135/HI sky130_fd_sc_hs__buf_2_23/X
+ sky130_fd_sc_hs__dlrtp_1_43/a_216_424# sky130_fd_sc_hs__dlrtp_1_43/a_759_508# sky130_fd_sc_hs__dlrtp_1_43/a_565_74#
+ sky130_fd_sc_hs__dlrtp_1_43/a_27_424# sky130_fd_sc_hs__dlrtp_1_43/a_1045_74# sky130_fd_sc_hs__dlrtp_1_43/a_643_74#
+ sky130_fd_sc_hs__dlrtp_1_43/a_817_48# sky130_fd_sc_hs__dlrtp_1_43/a_568_392# sky130_fd_sc_hs__dlrtp_1_43/a_363_74#
+ sky130_fd_sc_hs__dlrtp_1_43/a_769_74# sky130_fd_sc_hs__dlrtp_1
Xsky130_fd_sc_hs__dlrtp_1_53 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__dlrtp_1_53/Q
+ sky130_fd_sc_hs__clkbuf_16_53/A sky130_fd_sc_hs__conb_1_123/HI sky130_fd_sc_hs__dlrtp_1_53/D
+ sky130_fd_sc_hs__dlrtp_1_53/a_216_424# sky130_fd_sc_hs__dlrtp_1_53/a_759_508# sky130_fd_sc_hs__dlrtp_1_53/a_565_74#
+ sky130_fd_sc_hs__dlrtp_1_53/a_27_424# sky130_fd_sc_hs__dlrtp_1_53/a_1045_74# sky130_fd_sc_hs__dlrtp_1_53/a_643_74#
+ sky130_fd_sc_hs__dlrtp_1_53/a_817_48# sky130_fd_sc_hs__dlrtp_1_53/a_568_392# sky130_fd_sc_hs__dlrtp_1_53/a_363_74#
+ sky130_fd_sc_hs__dlrtp_1_53/a_769_74# sky130_fd_sc_hs__dlrtp_1
Xsky130_fd_sc_hs__dlrtp_1_64 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__dlrtp_1_65/Q
+ sky130_fd_sc_hs__clkbuf_16_53/A sky130_fd_sc_hs__conb_1_129/HI sky130_fd_sc_hs__dlrtp_1_65/D
+ sky130_fd_sc_hs__dlrtp_1_65/a_216_424# sky130_fd_sc_hs__dlrtp_1_65/a_759_508# sky130_fd_sc_hs__dlrtp_1_65/a_565_74#
+ sky130_fd_sc_hs__dlrtp_1_65/a_27_424# sky130_fd_sc_hs__dlrtp_1_65/a_1045_74# sky130_fd_sc_hs__dlrtp_1_65/a_643_74#
+ sky130_fd_sc_hs__dlrtp_1_65/a_817_48# sky130_fd_sc_hs__dlrtp_1_65/a_568_392# sky130_fd_sc_hs__dlrtp_1_65/a_363_74#
+ sky130_fd_sc_hs__dlrtp_1_65/a_769_74# sky130_fd_sc_hs__dlrtp_1
Xsky130_fd_sc_hs__dlrtp_1_75 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__dlrtp_1_75/Q
+ sky130_fd_sc_hs__clkbuf_16_53/X sky130_fd_sc_hs__conb_1_129/HI sky130_fd_sc_hs__buf_2_47/X
+ sky130_fd_sc_hs__dlrtp_1_75/a_216_424# sky130_fd_sc_hs__dlrtp_1_75/a_759_508# sky130_fd_sc_hs__dlrtp_1_75/a_565_74#
+ sky130_fd_sc_hs__dlrtp_1_75/a_27_424# sky130_fd_sc_hs__dlrtp_1_75/a_1045_74# sky130_fd_sc_hs__dlrtp_1_75/a_643_74#
+ sky130_fd_sc_hs__dlrtp_1_75/a_817_48# sky130_fd_sc_hs__dlrtp_1_75/a_568_392# sky130_fd_sc_hs__dlrtp_1_75/a_363_74#
+ sky130_fd_sc_hs__dlrtp_1_75/a_769_74# sky130_fd_sc_hs__dlrtp_1
Xsky130_fd_sc_hs__dlrtp_1_86 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__buf_2_159/A
+ sky130_fd_sc_hs__clkbuf_16_53/X sky130_fd_sc_hs__conb_1_137/HI sky130_fd_sc_hs__dlrtp_1_87/D
+ sky130_fd_sc_hs__dlrtp_1_87/a_216_424# sky130_fd_sc_hs__dlrtp_1_87/a_759_508# sky130_fd_sc_hs__dlrtp_1_87/a_565_74#
+ sky130_fd_sc_hs__dlrtp_1_87/a_27_424# sky130_fd_sc_hs__dlrtp_1_87/a_1045_74# sky130_fd_sc_hs__dlrtp_1_87/a_643_74#
+ sky130_fd_sc_hs__dlrtp_1_87/a_817_48# sky130_fd_sc_hs__dlrtp_1_87/a_568_392# sky130_fd_sc_hs__dlrtp_1_87/a_363_74#
+ sky130_fd_sc_hs__dlrtp_1_87/a_769_74# sky130_fd_sc_hs__dlrtp_1
Xsky130_fd_sc_hs__dlrtp_1_97 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__dlrtp_1_97/Q
+ sky130_fd_sc_hs__dlrtp_1_9/GATE sky130_fd_sc_hs__conb_1_133/HI sky130_fd_sc_hs__buf_2_98/X
+ sky130_fd_sc_hs__dlrtp_1_97/a_216_424# sky130_fd_sc_hs__dlrtp_1_97/a_759_508# sky130_fd_sc_hs__dlrtp_1_97/a_565_74#
+ sky130_fd_sc_hs__dlrtp_1_97/a_27_424# sky130_fd_sc_hs__dlrtp_1_97/a_1045_74# sky130_fd_sc_hs__dlrtp_1_97/a_643_74#
+ sky130_fd_sc_hs__dlrtp_1_97/a_817_48# sky130_fd_sc_hs__dlrtp_1_97/a_568_392# sky130_fd_sc_hs__dlrtp_1_97/a_363_74#
+ sky130_fd_sc_hs__dlrtp_1_97/a_769_74# sky130_fd_sc_hs__dlrtp_1
Xsky130_fd_sc_hs__einvp_2_2 DVSS: DVDD: DVDD: DVSS: dout_n sky130_fd_sc_hs__einvp_2_9/A
+ sky130_fd_sc_hs__einvp_2_3/TE sky130_fd_sc_hs__einvp_2_3/a_263_323# sky130_fd_sc_hs__einvp_2_3/a_36_74#
+ sky130_fd_sc_hs__einvp_2_3/a_27_368# sky130_fd_sc_hs__einvp_2
Xsky130_fd_sc_hs__clkbuf_2_5 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__dlrtp_1_53/D
+ sky130_fd_sc_hs__buf_2_45/X sky130_fd_sc_hs__clkbuf_2_5/a_43_192# sky130_fd_sc_hs__clkbuf_2
Xsky130_fd_sc_hs__clkbuf_2_16 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__dlrtp_1_69/D
+ sky130_fd_sc_hs__buf_2_69/X sky130_fd_sc_hs__clkbuf_2_17/a_43_192# sky130_fd_sc_hs__clkbuf_2
Xsky130_fd_sc_hs__clkbuf_2_27 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__o21ai_2_23/A2
+ sky130_fd_sc_hs__or2b_4_5/A sky130_fd_sc_hs__clkbuf_2_29/a_43_192# sky130_fd_sc_hs__clkbuf_2
Xsky130_fd_sc_hs__clkbuf_2_38 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__dlrtp_1_99/D
+ sky130_fd_sc_hs__buf_2_129/X sky130_fd_sc_hs__clkbuf_2_39/a_43_192# sky130_fd_sc_hs__clkbuf_2
Xsky130_fd_sc_hs__clkbuf_2_49 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__dlrtp_1_25/D
+ sky130_fd_sc_hs__o21ai_2_37/Y sky130_fd_sc_hs__clkbuf_2_49/a_43_192# sky130_fd_sc_hs__clkbuf_2
Xsky130_fd_sc_hs__buf_2_7 DVSS: DVDD: DVDD: DVSS: manual_control_osc[3] sky130_fd_sc_hs__buf_2_7/X
+ sky130_fd_sc_hs__buf_2_7/a_21_260# sky130_fd_sc_hs__buf_2
Xsky130_fd_sc_hs__dlrtp_1_9 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__dlrtp_1_9/Q sky130_fd_sc_hs__dlrtp_1_9/GATE
+ sky130_fd_sc_hs__conb_1_117/HI sky130_fd_sc_hs__dlrtp_1_9/D sky130_fd_sc_hs__dlrtp_1_9/a_216_424#
+ sky130_fd_sc_hs__dlrtp_1_9/a_759_508# sky130_fd_sc_hs__dlrtp_1_9/a_565_74# sky130_fd_sc_hs__dlrtp_1_9/a_27_424#
+ sky130_fd_sc_hs__dlrtp_1_9/a_1045_74# sky130_fd_sc_hs__dlrtp_1_9/a_643_74# sky130_fd_sc_hs__dlrtp_1_9/a_817_48#
+ sky130_fd_sc_hs__dlrtp_1_9/a_568_392# sky130_fd_sc_hs__dlrtp_1_9/a_363_74# sky130_fd_sc_hs__dlrtp_1_9/a_769_74#
+ sky130_fd_sc_hs__dlrtp_1
Xsky130_fd_sc_hs__buf_2_12 DVSS: DVDD: DVDD: DVSS: manual_control_osc[1] sky130_fd_sc_hs__buf_2_13/X
+ sky130_fd_sc_hs__buf_2_13/a_21_260# sky130_fd_sc_hs__buf_2
Xsky130_fd_sc_hs__buf_2_23 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__buf_2_41/X sky130_fd_sc_hs__buf_2_23/X
+ sky130_fd_sc_hs__buf_2_23/a_21_260# sky130_fd_sc_hs__buf_2
Xsky130_fd_sc_hs__buf_2_34 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__buf_2_35/A sky130_fd_sc_hs__buf_2_35/X
+ sky130_fd_sc_hs__buf_2_35/a_21_260# sky130_fd_sc_hs__buf_2
Xsky130_fd_sc_hs__buf_2_45 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__buf_2_45/A sky130_fd_sc_hs__buf_2_45/X
+ sky130_fd_sc_hs__buf_2_45/a_21_260# sky130_fd_sc_hs__buf_2
Xsky130_fd_sc_hs__buf_2_56 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__buf_2_57/A sky130_fd_sc_hs__buf_2_57/X
+ sky130_fd_sc_hs__buf_2_57/a_21_260# sky130_fd_sc_hs__buf_2
Xsky130_fd_sc_hs__buf_2_67 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__buf_2_67/A sky130_fd_sc_hs__buf_2_67/X
+ sky130_fd_sc_hs__buf_2_67/a_21_260# sky130_fd_sc_hs__buf_2
Xsky130_fd_sc_hs__buf_2_78 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__buf_2_79/A sky130_fd_sc_hs__buf_2_79/X
+ sky130_fd_sc_hs__buf_2_79/a_21_260# sky130_fd_sc_hs__buf_2
Xsky130_fd_sc_hs__buf_2_89 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__buf_2_89/A sky130_fd_sc_hs__buf_2_89/X
+ sky130_fd_sc_hs__buf_2_89/a_21_260# sky130_fd_sc_hs__buf_2
Xsky130_fd_sc_hs__o21bai_2_14 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__nand2_2_7/A
+ sky130_fd_sc_hs__o21bai_2_3/A2 sky130_fd_sc_hs__dlrtp_1_87/D sky130_fd_sc_hs__buf_2_67/A
+ sky130_fd_sc_hs__o21bai_2_15/a_27_74# sky130_fd_sc_hs__o21bai_2_15/a_225_74# sky130_fd_sc_hs__o21bai_2_15/a_507_368#
+ sky130_fd_sc_hs__o21bai_2
Xsky130_fd_sc_hs__o21bai_2_25 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__buf_8_3/X sky130_fd_sc_hs__clkbuf_4_81/X
+ sky130_fd_sc_hs__buf_2_101/X sky130_fd_sc_hs__buf_2_98/A sky130_fd_sc_hs__o21bai_2_25/a_27_74#
+ sky130_fd_sc_hs__o21bai_2_25/a_225_74# sky130_fd_sc_hs__o21bai_2_25/a_507_368# sky130_fd_sc_hs__o21bai_2
Xsky130_fd_sc_hs__o21bai_2_36 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__o21ai_4_1/A1
+ sky130_fd_sc_hs__clkinv_4_3/Y sky130_fd_sc_hs__dlrtp_1_21/D sky130_fd_sc_hs__o21bai_2_37/Y
+ sky130_fd_sc_hs__o21bai_2_37/a_27_74# sky130_fd_sc_hs__o21bai_2_37/a_225_74# sky130_fd_sc_hs__o21bai_2_37/a_507_368#
+ sky130_fd_sc_hs__o21bai_2
Xsky130_fd_sc_hs__o21bai_2_47 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__clkinv_4_3/Y
+ sky130_fd_sc_hs__or2b_2_1/X sky130_fd_sc_hs__dlrtp_1_115/D sky130_fd_sc_hs__buf_2_121/A
+ sky130_fd_sc_hs__o21bai_2_47/a_27_74# sky130_fd_sc_hs__o21bai_2_47/a_225_74# sky130_fd_sc_hs__o21bai_2_47/a_507_368#
+ sky130_fd_sc_hs__o21bai_2
Xsky130_fd_sc_hs__o21bai_2_58 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__nand2_2_9/B
+ sky130_fd_sc_hs__o21bai_2_3/A2 sky130_fd_sc_hs__clkbuf_2_7/X sky130_fd_sc_hs__buf_2_37/A
+ sky130_fd_sc_hs__o21bai_2_59/a_27_74# sky130_fd_sc_hs__o21bai_2_59/a_225_74# sky130_fd_sc_hs__o21bai_2_59/a_507_368#
+ sky130_fd_sc_hs__o21bai_2
Xsky130_fd_sc_hs__o21bai_2_69 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__inv_8_1/Y sky130_fd_sc_hs__nand2_2_9/B
+ sky130_fd_sc_hs__dlrtp_1_153/D sky130_fd_sc_hs__o21bai_2_69/Y sky130_fd_sc_hs__o21bai_2_69/a_27_74#
+ sky130_fd_sc_hs__o21bai_2_69/a_225_74# sky130_fd_sc_hs__o21bai_2_69/a_507_368# sky130_fd_sc_hs__o21bai_2
Xsky130_fd_sc_hs__o21bai_4_3 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__o21bai_4_3/Y
+ sky130_fd_sc_hs__nand2_2_15/B sky130_fd_sc_hs__o21bai_4_3/A2 sky130_fd_sc_hs__dlrtp_1_25/D
+ sky130_fd_sc_hs__o21bai_4_3/a_28_368# sky130_fd_sc_hs__o21bai_4_3/a_27_74# sky130_fd_sc_hs__o21bai_4_3/a_828_48#
+ sky130_fd_sc_hs__o21bai_4
Xsky130_fd_sc_hs__conb_1_201 DVSS: DVDD: DVDD: DVSS: prbs_generator_syn_19/eqn[30]
+ sky130_fd_sc_hs__conb_1_201/HI sky130_fd_sc_hs__conb_1_201/a_165_290# sky130_fd_sc_hs__conb_1_201/a_21_290#
+ sky130_fd_sc_hs__conb_1
Xsky130_fd_sc_hs__conb_1_212 DVSS: DVDD: DVDD: DVSS: prbs_generator_syn_21/eqn[31]
+ prbs_generator_syn_21/cke sky130_fd_sc_hs__conb_1_213/a_165_290# sky130_fd_sc_hs__conb_1_213/a_21_290#
+ sky130_fd_sc_hs__conb_1
Xsky130_fd_sc_hs__conb_1_223 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__conb_1_223/LO
+ sky130_fd_sc_hs__conb_1_223/HI sky130_fd_sc_hs__conb_1_223/a_165_290# sky130_fd_sc_hs__conb_1_223/a_21_290#
+ sky130_fd_sc_hs__conb_1
Xsky130_fd_sc_hs__conb_1_234 DVSS: DVDD: DVDD: DVSS: prbs_generator_syn_27/eqn[8]
+ prbs_generator_syn_27/eqn[1] sky130_fd_sc_hs__conb_1_235/a_165_290# sky130_fd_sc_hs__conb_1_235/a_21_290#
+ sky130_fd_sc_hs__conb_1
Xsky130_fd_sc_hs__conb_1_245 DVSS: DVDD: DVDD: DVSS: prbs_generator_syn_31/eqn[21]
+ prbs_generator_syn_31/eqn[20] sky130_fd_sc_hs__conb_1_245/a_165_290# sky130_fd_sc_hs__conb_1_245/a_21_290#
+ sky130_fd_sc_hs__conb_1
Xsky130_fd_sc_hs__conb_1_256 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__conb_1_257/LO
+ sky130_fd_sc_hs__conb_1_257/HI sky130_fd_sc_hs__conb_1_257/a_165_290# sky130_fd_sc_hs__conb_1_257/a_21_290#
+ sky130_fd_sc_hs__conb_1
Xsky130_fd_sc_hs__conb_1_267 DVSS: DVDD: DVDD: DVSS: prbs_generator_syn_31/eqn[8]
+ sky130_fd_sc_hs__conb_1_267/HI sky130_fd_sc_hs__conb_1_267/a_165_290# sky130_fd_sc_hs__conb_1_267/a_21_290#
+ sky130_fd_sc_hs__conb_1
Xsky130_fd_sc_hs__clkbuf_8_15 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__clkbuf_8_15/X
+ sky130_fd_sc_hs__clkbuf_8_15/A sky130_fd_sc_hs__clkbuf_8_15/a_125_368# sky130_fd_sc_hs__clkbuf_8
Xsky130_fd_sc_hs__clkbuf_8_26 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__clkbuf_8_27/X
+ sky130_fd_sc_hs__clkbuf_8_27/A sky130_fd_sc_hs__clkbuf_8_27/a_125_368# sky130_fd_sc_hs__clkbuf_8
Xsky130_fd_sc_hs__clkbuf_8_37 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__nand2_2_15/B
+ sky130_fd_sc_hs__or2b_2_1/X sky130_fd_sc_hs__clkbuf_8_37/a_125_368# sky130_fd_sc_hs__clkbuf_8
Xsky130_fd_sc_hs__clkbuf_8_48 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__nand2_2_5/B
+ sky130_fd_sc_hs__or2b_4_3/X sky130_fd_sc_hs__clkbuf_8_49/a_125_368# sky130_fd_sc_hs__clkbuf_8
Xsky130_fd_sc_hs__clkbuf_8_59 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__or4_2_1/A sky130_fd_sc_hs__clkbuf_8_59/A
+ sky130_fd_sc_hs__clkbuf_8_59/a_125_368# sky130_fd_sc_hs__clkbuf_8
Xsky130_fd_sc_hs__o21bai_2_0 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__o21bai_2_3/A2
+ sky130_fd_sc_hs__nand2_2_3/B sky130_fd_sc_hs__dlrtp_1_53/D sky130_fd_sc_hs__buf_2_25/A
+ sky130_fd_sc_hs__o21bai_2_1/a_27_74# sky130_fd_sc_hs__o21bai_2_1/a_225_74# sky130_fd_sc_hs__o21bai_2_1/a_507_368#
+ sky130_fd_sc_hs__o21bai_2
Xsky130_fd_sc_hs__nand2_2_8 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__inv_4_15/A sky130_fd_sc_hs__nand2_2_9/B
+ sky130_fd_sc_hs__buf_2_65/X sky130_fd_sc_hs__nand2_2_9/a_27_74# sky130_fd_sc_hs__nand2_2
Xsky130_fd_sc_hs__or2b_4_4 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__or2b_4_5/A sky130_fd_sc_hs__or4_2_1/A
+ sky130_fd_sc_hs__or2b_4_5/X sky130_fd_sc_hs__or2b_4_5/a_676_48# sky130_fd_sc_hs__or2b_4_5/a_489_392#
+ sky130_fd_sc_hs__or2b_4_5/a_81_296# sky130_fd_sc_hs__or2b_4
Xprbs_generator_syn_10 prbs_generator_syn_9/clk prbs_generator_syn_9/rst prbs_generator_syn_11/cke
+ sky130_fd_sc_hs__conb_1_91/LO sky130_fd_sc_hs__conb_1_91/LO sky130_fd_sc_hs__conb_1_91/LO
+ sky130_fd_sc_hs__conb_1_91/LO sky130_fd_sc_hs__conb_1_91/HI sky130_fd_sc_hs__conb_1_91/HI
+ sky130_fd_sc_hs__conb_1_91/HI sky130_fd_sc_hs__conb_1_91/HI sky130_fd_sc_hs__conb_1_91/HI
+ sky130_fd_sc_hs__conb_1_91/HI sky130_fd_sc_hs__conb_1_91/HI prbs_generator_syn_11/cke
+ prbs_generator_syn_11/cke prbs_generator_syn_11/cke sky130_fd_sc_hs__conb_1_81/LO
+ prbs_generator_syn_11/cke sky130_fd_sc_hs__conb_1_81/LO prbs_generator_syn_11/cke
+ prbs_generator_syn_11/eqn[2] prbs_generator_syn_11/eqn[2] prbs_generator_syn_11/eqn[2]
+ prbs_generator_syn_11/eqn[2] prbs_generator_syn_11/eqn[2] prbs_generator_syn_11/eqn[2]
+ sky130_fd_sc_hs__conb_1_89/LO sky130_fd_sc_hs__conb_1_89/HI sky130_fd_sc_hs__conb_1_89/HI
+ sky130_fd_sc_hs__conb_1_89/LO sky130_fd_sc_hs__conb_1_89/LO sky130_fd_sc_hs__conb_1_89/HI
+ sky130_fd_sc_hs__conb_1_89/HI sky130_fd_sc_hs__conb_1_89/LO sky130_fd_sc_hs__conb_1_81/LO
+ sky130_fd_sc_hs__conb_1_79/LO sky130_fd_sc_hs__conb_1_79/LO sky130_fd_sc_hs__conb_1_77/LO
+ sky130_fd_sc_hs__conb_1_77/LO sky130_fd_sc_hs__conb_1_77/LO sky130_fd_sc_hs__conb_1_77/LO
+ sky130_fd_sc_hs__conb_1_77/LO sky130_fd_sc_hs__conb_1_65/LO sky130_fd_sc_hs__conb_1_65/LO
+ sky130_fd_sc_hs__conb_1_65/LO sky130_fd_sc_hs__conb_1_65/HI sky130_fd_sc_hs__conb_1_65/LO
+ sky130_fd_sc_hs__conb_1_65/LO sky130_fd_sc_hs__conb_1_65/LO sky130_fd_sc_hs__conb_1_65/LO
+ prbs_generator_syn_7/eqn[0] prbs_generator_syn_7/eqn[0] prbs_generator_syn_7/eqn[0]
+ prbs_generator_syn_7/eqn[0] prbs_generator_syn_7/eqn[0] prbs_generator_syn_7/eqn[0]
+ prbs_generator_syn_11/eqn[9] prbs_generator_syn_11/eqn[9] prbs_generator_syn_11/eqn[9]
+ prbs_generator_syn_11/eqn[9] prbs_generator_syn_11/eqn[9] prbs_generator_syn_11/eqn[9]
+ prbs_generator_syn_11/eqn[9] prbs_generator_syn_11/eqn[2] prbs_generator_syn_11/eqn[1]
+ prbs_generator_syn_11/eqn[2] prbs_generator_syn_9/inj_err sky130_fd_sc_hs__conb_1_81/LO
+ sky130_fd_sc_hs__conb_1_81/LO prbs_generator_syn_11/out DVSS: DVDD: prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_1/a_293_74#
+ prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_15/X prbs_generator_syn_11/sky130_fd_sc_hs__nand2_1_35/B
+ prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_51/Y prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_9/A
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_9/CLK prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_47/a_27_74#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_37/a_1226_296# prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_3/B
+ prbs_generator_syn_11/sky130_fd_sc_hs__nor2b_1_7/a_27_112# prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_29/B
+ prbs_generator_syn_11/sky130_fd_sc_hs__sdlclkp_2_1/a_580_74# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_1/a_1141_508#
+ prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_5/Y prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_41/a_230_79#
+ prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_61/a_138_385# prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_43/a_132_392#
+ prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_3/a_222_392# prbs_generator_syn_11/sky130_fd_sc_hs__nor2b_1_9/a_27_112#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_61/a_27_74# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_35/a_206_368#
+ prbs_generator_syn_11/sky130_fd_sc_hs__nand2_2_3/Y prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_25/B
+ prbs_generator_syn_11/sky130_fd_sc_hs__nand2_1_11/a_117_74# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_67/a_651_503#
+ prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_45/X prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_39/a_696_458#
+ prbs_generator_syn_11/sky130_fd_sc_hs__sdlclkp_2_1/a_1198_74# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_45/a_1034_424#
+ prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_17/a_222_392# prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_55/a_222_392#
+ prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_53/Y prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_35/A
+ prbs_generator_syn_11/m3_13600_1651# prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_59/a_52_123#
+ prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_5/a_293_74# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_35/a_1226_296#
+ prbs_generator_syn_11/sky130_fd_sc_hs__nand2_1_51/B prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_5/a_651_503#
+ prbs_generator_syn_11/sky130_fd_sc_hs__nand2_1_21/B prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_8/a_27_74#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_15/a_27_74# prbs_generator_syn_11/sky130_fd_sc_hs__and2b_2_1/X
+ prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_13/X prbs_generator_syn_11/sky130_fd_sc_hs__nand2_2_3/a_27_74#
+ prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_50/a_138_385# prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_33/a_132_392#
+ prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_1/a_376_368# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_25/a_206_368#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_35/a_437_503# prbs_generator_syn_11/sky130_fd_sc_hs__sdlclkp_2_1/a_708_451#
+ prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_45/a_230_79# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_29/a_696_458#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_32/a_27_74# prbs_generator_syn_11/sky130_fd_sc_hs__nor2b_1_4/Y
+ prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_59/a_293_74# prbs_generator_syn_11/sky130_fd_sc_hs__nand2_1_47/a_117_74#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_73/a_735_102# prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_21/a_112_119#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_23/a_1141_508# prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_25/a_293_74#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_7/Q prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_3/a_112_119#
+ prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_35/B prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_51/X
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_53/a_1178_124# prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_23/a_132_392#
+ prbs_generator_syn_11/sky130_fd_sc_hs__nand2_1_3/B prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_15/a_206_368#
+ prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_63/a_132_392# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_55/a_27_74#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_25/a_437_503# prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_41/a_52_123#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_47/a_651_503# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_73/a_1141_508#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_19/a_696_458# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_57/a_696_458#
+ prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_7/X prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_43/a_1034_424#
+ prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_55/A prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_11/a_112_119#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_21/a_1141_508# prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_35/a_222_392#
+ prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_49/a_230_79# prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_67/Y
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_71/a_27_74# prbs_generator_syn_11/sky130_fd_sc_hs__nand2_1_33/B
+ prbs_generator_syn_11/sky130_fd_sc_hs__conb_1_1/LO prbs_generator_syn_11/sky130_fd_sc_hs__nand2_1_19/a_117_74#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_51/a_1178_124# prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_33/X
+ prbs_generator_syn_11/sky130_fd_sc_hs__nand2_1_29/B prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_41/Y
+ prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_53/a_132_392# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_45/a_206_368#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_15/a_437_503# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_37/a_651_503#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_39/a_544_485# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_53/a_735_102#
+ prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_45/a_52_123# prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_1/B
+ prbs_generator_syn_11/sky130_fd_sc_hs__nand2_2_3/B prbs_generator_syn_11/sky130_fd_sc_hs__clkbuf_16_1/A
+ prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_21/X prbs_generator_syn_11/sky130_fd_sc_hs__nand2_1_25/B
+ prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_39/a_376_368# prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_63/X
+ prbs_generator_syn_11/m3_13600_3481# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_69/a_1178_124#
+ prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_21/a_138_385# prbs_generator_syn_11/sky130_fd_sc_hs__nor2b_1_8/Y
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_19/a_1178_124# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_49/a_27_74#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_45/a_437_503# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_27/a_651_503#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_71/a_1141_508# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_65/a_651_503#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_29/a_544_485# prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_3/a_138_385#
+ prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_55/X prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_43/a_735_102#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_41/a_1034_424# prbs_generator_syn_11/sky130_fd_sc_hs__nand2_1_9/B
+ prbs_generator_syn_11/sky130_fd_sc_hs__nor2b_1_9/Y prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_59/a_1034_424#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_39/a_1141_508# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_33/a_1226_296#
+ prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_49/a_52_123# prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_47/Y
+ prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_43/Y prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_4/a_651_503#
+ prbs_generator_syn_11/sky130_fd_sc_hs__nand2_1_49/B prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_19/A
+ prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_11/a_138_385# prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_5/X
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_63/a_206_368# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_17/a_651_503#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_19/a_544_485# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_55/a_651_503#
+ prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_9/Y prbs_generator_syn_11/sky130_fd_sc_hs__nand2_1_17/B
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_57/a_544_485# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_67/a_696_458#
+ prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_35/X prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_19/a_27_74#
+ prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_45/a_222_392# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_32/a_1226_296#
+ prbs_generator_syn_11/sky130_fd_sc_hs__nand2_1_43/B prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_25/A
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_1/a_206_368# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_49/a_1226_296#
+ prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_1/a_112_119# prbs_generator_syn_11/sky130_fd_sc_hs__or2_1_1/X
+ prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_59/a_376_368# prbs_generator_syn_11/sky130_fd_sc_hs__nand2_1_19/B
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_5/a_696_458# prbs_generator_syn_11/sky130_fd_sc_hs__nor2b_1_1/Y
+ prbs_generator_syn_11/sky130_fd_sc_hs__nor2b_1_5/a_278_368# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_17/a_1178_124#
+ prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_39/X prbs_generator_syn_11/m3_13600_5433#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_63/a_437_503# prbs_generator_syn_11/sky130_fd_sc_hs__nand2_2_5/B
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_23/a_735_102# prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_53/A
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_61/a_735_102# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_57/a_1034_424#
+ prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_63/B prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_37/a_1141_508#
+ prbs_generator_syn_11/sky130_fd_sc_hs__nand2_1_47/B prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_29/X
+ prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_65/Y prbs_generator_syn_11/m3_13600_4701#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_1/a_437_503# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_67/a_1178_124#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_9/a_735_102# prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_13/a_132_392#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_15/a_1178_124# prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_15/A
+ prbs_generator_syn_11/sky130_fd_sc_hs__nand2_1_1/B prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_43/B
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_35/a_651_503# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_8/D
+ prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_29/A prbs_generator_syn_11/sky130_fd_sc_hs__nand2_1_7/B
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_13/a_735_102# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_47/a_696_458#
+ prbs_generator_syn_11/sky130_fd_sc_hs__nand2_1_31/B prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_51/a_735_102#
+ prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_59/X prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_35/a_1141_508#
+ prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_25/a_222_392# prbs_generator_syn_11/sky130_fd_sc_hs__sdlclkp_2_1/a_288_48#
+ prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_55/B prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_17/B
+ prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_43/A prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_7/A
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_65/a_1178_124# prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_59/Y
+ prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_41/X prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_21/a_230_79#
+ prbs_generator_syn_11/sky130_fd_sc_hs__nand2_1_57/a_117_74# prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_1/a_222_392#
+ prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_19/B prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_35/a_293_74#
+ prbs_generator_syn_11/sky130_fd_sc_hs__nand2_1_23/a_117_74# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_73/a_206_368#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_25/a_651_503# prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_1/a_138_385#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_37/a_696_458# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_67/a_544_485#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_43/a_27_74# prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_9/X
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_55/a_1034_424# prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_39/a_112_119#
+ prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_15/a_222_392# prbs_generator_syn_11/sky130_fd_sc_hs__conb_1_1/HI
+ prbs_generator_syn_11/sky130_fd_sc_hs__nand2_1_23/B prbs_generator_syn_11/sky130_fd_sc_hs__nand2_1_53/B
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_9/a_1178_124# prbs_generator_syn_11/sky130_fd_sc_hs__nor2b_1_4/A
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_47/a_1226_296# prbs_generator_syn_11/m3_13600_11045#
+ prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_17/X prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_29/a_376_368#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_5/a_544_485# prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_3/X
+ prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_31/a_132_392# prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_61/A
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_15/a_651_503# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_73/a_437_503#
+ prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_25/a_230_79# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_27/a_696_458#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_65/a_696_458# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_33/a_735_102#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_71/a_735_102# prbs_generator_syn_11/m3_13600_7263#
+ prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_43/a_222_392# prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_50/Y
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_8/a_1178_124# prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_53/B
+ prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_19/a_376_368# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_63/a_1178_124#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_4/a_696_458# prbs_generator_syn_11/sky130_fd_sc_hs__nor2b_1_4/a_278_368#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_13/a_1178_124# prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_61/a_132_392#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_53/a_206_368# prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_21/a_52_123#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_45/a_651_503# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_17/a_696_458#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_47/a_544_485# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_55/a_696_458#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_21/a_735_102# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_37/a_27_74#
+ prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_61/B prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_61/X
+ prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_59/a_112_119# prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_31/A
+ prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_33/a_222_392# prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_29/a_230_79#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_45/a_1226_296# prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_9/a_132_392#
+ prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_5/A prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_57/Y
+ prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_31/X prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_51/a_27_74#
+ prbs_generator_syn_11/sky130_fd_sc_hs__nor2b_1_8/a_27_112# prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_47/a_376_368#
+ prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_53/a_293_74# prbs_generator_syn_11/sky130_fd_sc_hs__nand2_1_43/a_117_74#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_8/a_735_102# prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_21/a_293_74#
+ prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_39/a_138_385# prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_63/Y
+ prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_51/a_132_392# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_43/a_206_368#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_53/a_437_503# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_37/a_544_485#
+ prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_57/X prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_53/a_1034_424#
+ prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_25/a_52_123# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_33/a_1141_508#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_63/Q prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_23/a_222_392#
+ prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_63/a_222_392# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_7/a_1178_124#
+ prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_53/X prbs_generator_syn_11/sky130_fd_sc_hs__nand2_2_5/Y
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_61/a_1178_124# prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_1/a_230_79#
+ prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_43/a_230_79# prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_11/a_230_79#
+ prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_41/a_132_392# prbs_generator_syn_11/sky130_fd_sc_hs__nand2_1_13/a_117_74#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_43/a_437_503# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_27/a_544_485#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_63/a_651_503# prbs_generator_syn_11/sky130_fd_sc_hs__nand2_1_7/a_117_74#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_35/a_696_458# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_65/a_544_485#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_51/a_1034_424# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_41/a_735_102#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_32/a_1141_508# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_49/a_1141_508#
+ prbs_generator_syn_11/sky130_fd_sc_hs__nand2_1_55/B prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_53/a_222_392#
+ prbs_generator_syn_11/sky130_fd_sc_hs__sdlclkp_2_1/a_114_112# prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_9/a_293_74#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_43/a_1226_296# prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_29/a_52_123#
+ prbs_generator_syn_11/sky130_fd_sc_hs__nand2_1_37/B prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_1/a_651_503#
+ prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_27/a_376_368# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_4/a_544_485#
+ prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_67/a_376_368# prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_27/X
+ prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_1/X prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_59/a_138_385#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_29/a_1178_124# prbs_generator_syn_11/m3_13600_2871#
+ prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_5/a_230_79# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_23/a_206_368#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_61/a_206_368# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_17/a_544_485#
+ prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_15/a_230_79# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_25/a_696_458#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_55/a_544_485# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_32/a_735_102#
+ prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_29/a_293_74# prbs_generator_syn_11/sky130_fd_sc_hs__nand2_1_17/a_117_74#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_69/a_1034_424# prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_29/a_112_119#
+ prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_37/X prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_31/B
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_19/a_1034_424# prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_33/A
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_9/a_206_368# prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_57/a_376_368#
+ prbs_generator_syn_11/sky130_fd_sc_hs__sdlclkp_2_1/a_706_317# prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_11/B
+ prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_1/a_52_123# prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_39/B
+ prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_21/a_132_392# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_13/a_206_368#
+ prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_43/a_52_123# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_51/a_206_368#
+ prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_47/X prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_23/a_437_503#
+ prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_11/a_52_123# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_61/a_437_503#
+ prbs_generator_syn_11/sky130_fd_sc_hs__nor2b_1_7/Y prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_51/A
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_15/a_696_458# prbs_generator_syn_11/sky130_fd_sc_hs__nor2b_1_5/Y
+ prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_9/a_230_79# prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_25/X
+ prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_19/a_112_119# prbs_generator_syn_11/sky130_fd_sc_hs__nand2_1_45/B
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_5/a_1178_124# prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_19/a_230_79#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_41/a_1226_296# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_59/a_1226_296#
+ prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_63/a_230_79# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_51/Q
+ prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_7/a_132_392# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_9/a_437_503#
+ prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_46/a_376_368# prbs_generator_syn_11/sky130_fd_sc_hs__nand2_1_33/a_117_74#
+ prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_11/a_293_74# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_27/a_1178_124#
+ prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_11/a_132_392# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_13/a_437_503#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_51/a_437_503# prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_5/a_52_123#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_35/a_544_485# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_73/a_651_503#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_45/a_696_458# prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_15/a_52_123#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_47/a_1141_508# prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_47/a_112_119#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_4/a_1178_124# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_17/a_1034_424#
+ prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_23/B prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_37/a_376_368#
+ prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_15/B prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_7/Y
+ prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_29/a_138_385# prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_33/a_230_79#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_25/a_1178_124# prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_47/a_293_74#
+ prbs_generator_syn_11/sky130_fd_sc_hs__nand2_1_37/a_117_74# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_33/a_206_368#
+ prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_15/a_293_74# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_71/a_206_368#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_25/a_544_485# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_67/a_1034_424#
+ prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_13/a_222_392# prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_9/a_52_123#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_15/a_1034_424# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_57/a_1226_296#
+ prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_19/a_52_123# prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_23/X
+ prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_63/a_52_123# prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_19/a_138_385#
+ prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_9/a_376_368# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_21/a_206_368#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_33/a_437_503# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_71/a_437_503#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_53/a_651_503# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_15/a_544_485#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_63/a_696_458# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_65/a_1034_424#
+ prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_19/a_293_74# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_45/a_1141_508#
+ prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_27/a_112_119# prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_67/a_112_119#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_1/a_1178_124# prbs_generator_syn_11/sky130_fd_sc_hs__conb_1_1/a_21_290#
+ prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_63/a_293_74# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_8/a_206_368#
+ prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_17/a_376_368# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_63/a_27_74#
+ prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_21/A prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_55/a_376_368#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_1/a_696_458# prbs_generator_syn_11/sky130_fd_sc_hs__nor2b_1_1/a_278_368#
+ prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_47/a_138_385# prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_33/a_52_123#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_9/a_1034_424# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_21/a_437_503#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_1/a_27_74# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_43/a_651_503#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_1/Q prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_45/a_544_485#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_69/a_735_102# prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_57/a_112_119#
+ prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_31/a_222_392# prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_13/A
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_55/a_1226_296# prbs_generator_syn_11/sky130_fd_sc_hs__nand2_2_5/a_27_74#
+ prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_53/a_230_79# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_8/a_437_503#
+ prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_67/a_293_74# prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_33/a_293_74#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_7/a_735_102# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_23/a_1178_124#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_41/a_206_368# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_8/a_1034_424#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_63/a_1034_424# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_59/a_735_102#
+ prbs_generator_syn_11/sky130_fd_sc_hs__nand2_1_5/B prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_43/a_1141_508#
+ prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_46/a_112_119# prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_61/a_222_392#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_13/a_1034_424# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_73/a_1178_124#
+ prbs_generator_syn_11/sky130_fd_sc_hs__nand2_1_27/B prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_13/B
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_57/a_27_74# prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_57/a_230_79#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_21/a_1178_124# prbs_generator_syn_11/sky130_fd_sc_hs__nor2b_1_1/a_27_112#
+ prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_27/a_138_385# prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_23/a_230_79#
+ prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_67/a_138_385# prbs_generator_syn_11/sky130_fd_sc_hs__nand2_1_41/B
+ prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_9/a_222_392# prbs_generator_syn_11/sky130_fd_sc_hs__nand2_1_27/a_117_74#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_32/a_206_368# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_23/a_651_503#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_41/a_437_503# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_73/a_27_74#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_61/a_651_503# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_63/a_544_485#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_49/a_735_102# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_73/a_696_458#
+ prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_37/a_112_119# prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_51/a_222_392#
+ prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_43/X prbs_generator_syn_11/sky130_fd_sc_hs__nand2_2_1/B
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_9/a_651_503# prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_53/a_52_123#
+ prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_49/X prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_25/a_376_368#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_1/a_544_485# prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_65/a_376_368#
+ prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_57/a_138_385# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_27/a_27_74#
+ prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_39/a_132_392# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_7/a_1034_424#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_13/a_651_503# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_32/a_437_503#
+ prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_27/a_230_79# prbs_generator_syn_11/m3_13600_12265#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_51/a_651_503# prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_59/B
+ prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_47/A prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_61/a_1034_424#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_41/a_1141_508# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_59/a_1141_508#
+ prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_41/a_222_392# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_53/a_1226_296#
+ prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_3/A prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_71/a_1178_124#
+ prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_9/a_112_119# prbs_generator_syn_11/sky130_fd_sc_hs__nand2_1_3/a_117_74#
+ prbs_generator_syn_11/m3_13600_8483# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_39/a_1178_124#
+ prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_57/a_52_123# prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_46/a_138_385#
+ prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_23/a_52_123# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_67/a_27_74#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_53/a_696_458# prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_17/a_112_119#
+ prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_11/A prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_55/a_112_119#
+ prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_1/A prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_51/a_1226_296#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_29/a_1034_424# prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_59/A
+ prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_23/A prbs_generator_syn_11/sky130_fd_sc_hs__nand2_1_39/B
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_5/a_27_74# prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_57/a_293_74#
+ prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_37/a_138_385# prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_59/a_132_392#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_33/a_651_503# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_71/a_651_503#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_43/a_696_458# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_73/a_544_485#
+ prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_27/a_52_123# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_57/a_1141_508#
+ prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_21/a_222_392# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_35/a_27_74#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_69/a_1226_296# prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_37/B
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_19/a_1226_296# prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_35/a_376_368#
+ prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_47/a_230_79# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_37/a_1178_124#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_5/a_1034_424# prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_49/a_132_392#
+ prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_7/a_222_392# prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_27/a_293_74#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_21/a_651_503# prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_9/a_138_385#
+ prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_11/a_222_392# prbs_generator_syn_11/m3_13600_14095#
+ prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_50/A prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_27/a_1034_424#
+ prbs_generator_syn_11/sky130_fd_sc_hs__nand2_1_13/B prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_8/a_651_503#
+ prbs_generator_syn_11/m3_13600_9703# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_35/a_1178_124#
+ prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_17/a_138_385# prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_55/a_138_385#
+ prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_7/a_230_79# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_4/a_1034_424#
+ prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_7/a_376_368# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_69/a_206_368#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_23/a_696_458# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_53/a_544_485#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_39/a_735_102# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_61/a_696_458#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_55/a_1141_508# prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_25/a_112_119#
+ prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_65/a_112_119# prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_43/a_293_74#
+ prbs_generator_syn_11/sky130_fd_sc_hs__nand2_1_57/B prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_25/a_1034_424#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_7/a_206_368# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_17/a_1226_296#
+ prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_15/a_376_368# prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_53/a_376_368#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_9/a_696_458# prbs_generator_syn_11/m3_13600_431#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_45/a_27_74# prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_47/a_52_123#
+ prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_29/a_132_392# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_59/a_206_368#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_69/a_437_503# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_41/a_651_503#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_43/a_544_485# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_13/a_696_458#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_29/a_735_102# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_51/a_696_458#
+ prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_61/Y prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_67/a_1226_296#
+ prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_5/a_132_392# prbs_generator_syn_11/sky130_fd_sc_hs__and2b_2_1/a_198_48#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_7/a_437_503# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_15/a_1226_296#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_69/a_27_74# prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_46/a_293_74#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_1/a_1034_424# prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_19/a_132_392#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_49/a_206_368# prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_7/a_52_123#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_59/a_437_503# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_32/a_651_503#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_7/a_27_74# prbs_generator_syn_11/sky130_fd_sc_hs__nand2_2_1/a_27_74#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_19/a_735_102# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_57/a_735_102#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_65/a_1226_296# prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_37/A
+ prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_33/a_376_368# prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_37/a_230_79#
+ prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_25/a_138_385# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_39/a_27_74#
+ prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_65/a_138_385# prbs_generator_syn_11/sky130_fd_sc_hs__nor2b_1_9/a_278_368#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_49/a_437_503# prbs_generator_syn_11/sky130_fd_sc_hs__and2b_2_1/a_505_74#
+ prbs_generator_syn_11/sky130_fd_sc_hs__nand2_1_51/a_117_74# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_23/a_544_485#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_33/a_696_458# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_61/a_544_485#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_9/a_1226_296# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_53/a_1141_508#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_71/a_696_458# prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_35/a_112_119#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_23/a_1034_424# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_9/a_544_485#
+ prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_63/a_376_368# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_33/a_1178_124#
+ prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_5/a_376_368# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_13/a_544_485#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_73/a_1034_424# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_21/a_696_458#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_51/a_544_485# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_8/a_1226_296#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_51/a_1141_508# prbs_generator_syn_11/sky130_fd_sc_hs__nand2_1_55/a_117_74#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_21/a_1034_424# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_63/a_1226_296#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_23/a_27_74# prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_7/a_112_119#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_13/a_1226_296# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_8/a_696_458#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_32/a_1178_124# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_49/a_1178_124#
+ prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_37/a_52_123# prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_27/a_132_392#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_71/Q prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_67/a_735_102#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_69/a_1141_508# prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_15/a_112_119#
+ prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_53/a_112_119# prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_39/a_222_392#
+ prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_55/a_230_79# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_19/a_1141_508#
+ prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_37/a_293_74# prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_43/a_376_368#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_5/a_735_102# prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_35/a_138_385#
+ prbs_generator_syn_11/sky130_fd_sc_hs__sdlclkp_2_1/a_114_424# prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_57/a_132_392#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_71/a_1034_424# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_7/a_1226_296#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_33/a_544_485# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_41/a_696_458#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_71/a_544_485# prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_21/B
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_61/a_1226_296# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_39/a_1034_424#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_17/a_27_74# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_9/a_27_74#
+ prbs_generator_syn_11/sky130_fd_sc_hs__nor2b_1_5/a_27_112# prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_47/a_132_392#
+ prbs_generator_syn_11/sky130_fd_sc_hs__nor2b_1_8/a_278_368# prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_9/B
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_39/a_206_368# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_33/a_27_74#
+ prbs_generator_syn_11/sky130_fd_sc_hs__nand2_1_41/a_117_74# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_69/a_651_503#
+ prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_51/a_293_74# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_21/a_544_485#
+ prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_7/a_138_385# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_32/a_696_458#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_47/a_735_102# prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_33/a_112_119#
+ prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_59/a_222_392# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_17/a_1141_508#
+ prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_55/a_52_123# prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_3/a_293_74#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_7/a_651_503# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_29/a_1226_296#
+ prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_23/a_376_368# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_8/a_544_485#
+ prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_47/B prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_47/a_1178_124#
+ prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_15/a_138_385# prbs_generator_syn_11/sky130_fd_sc_hs__sdlclkp_2_1/a_1195_374#
+ prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_53/a_138_385# prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_37/a_132_392#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_29/a_206_368# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_39/a_437_503#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_59/a_651_503# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_37/a_735_102#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_67/a_1141_508# prbs_generator_syn_11/sky130_fd_sc_hs__and2b_2_1/a_27_74#
+ prbs_generator_syn_11/sky130_fd_sc_hs__conb_1_1/a_165_290# prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_55/a_293_74#
+ prbs_generator_syn_11/sky130_fd_sc_hs__nand2_1_45/a_117_74# prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_63/a_112_119#
+ prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_49/a_222_392# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_37/a_1034_424#
+ prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_23/a_293_74# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_15/a_1141_508#
+ prbs_generator_syn_11/sky130_fd_sc_hs__nand2_1_5/a_117_74# prbs_generator_syn_11/m3_13600_13485#
+ prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_5/a_112_119# prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_13/a_376_368#
+ prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_51/a_376_368# prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_7/a_293_74#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_19/a_206_368# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_57/a_206_368#
+ prbs_generator_syn_11/sky130_fd_sc_hs__sdlclkp_2_1/a_318_74# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_29/a_437_503#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_49/a_651_503# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_25/a_27_74#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_5/a_1226_296# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_41/a_544_485#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_27/a_735_102# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_65/a_1141_508#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_65/a_735_102# prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_3/a_230_79#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_35/a_1034_424# prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_13/a_230_79#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_41/a_27_74# prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_3/a_132_392#
+ prbs_generator_syn_11/sky130_fd_sc_hs__nand2_1_49/a_117_74# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_27/a_1226_296#
+ prbs_generator_syn_11/sky130_fd_sc_hs__nand2_1_15/a_117_74# prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_41/a_376_368#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_45/a_1178_124# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_4/a_735_102#
+ prbs_generator_syn_11/sky130_fd_sc_hs__nand2_1_9/a_117_74# prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_33/a_138_385#
+ prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_17/a_132_392# prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_55/a_132_392#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_9/a_1141_508# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_19/a_437_503#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_57/a_437_503# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_4/a_1226_296#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_32/a_544_485# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_17/a_735_102#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_55/a_735_102# prbs_generator_syn_11/m3_13600_2261#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_65/a_27_74# prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_29/a_222_392#
+ prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_43/a_112_119# prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_19/X
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_25/a_1226_296# prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_31/a_376_368#
+ prbs_generator_syn_11/sky130_fd_sc_hs__or2_1_1/a_63_368# prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_17/a_230_79#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_4/a_27_74# prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_61/a_230_79#
+ prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_63/a_138_385# prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_5/a_222_392#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_8/a_1141_508# prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_41/a_293_74#
+ prbs_generator_syn_11/sky130_fd_sc_hs__nand2_1_31/a_117_74# prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_5/a_138_385#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_63/a_1141_508# prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_19/a_222_392#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_13/a_1141_508# prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_3/a_52_123#
+ prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_13/a_52_123# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_43/a_1178_124#
+ prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_61/a_376_368# prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_35/a_132_392#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_67/a_206_368# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_1/a_1226_296#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_69/a_696_458# prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_31/a_230_79#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_35/a_735_102# prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_23/a_112_119#
+ prbs_generator_syn_11/sky130_fd_sc_hs__nand2_1_35/a_117_74# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_59/a_27_74#
+ prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_13/a_293_74# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_5/a_206_368#
+ prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_50/a_376_368# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_7/a_696_458#
+ prbs_generator_syn_11/sky130_fd_sc_hs__nor2b_1_7/a_278_368# prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_17/a_52_123#
+ prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_43/a_138_385# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_7/a_1141_508#
+ prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_61/a_52_123# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_67/a_437_503#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_61/a_1141_508# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_25/a_735_102#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_59/a_696_458# prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_13/a_112_119#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_33/a_1034_424# prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_51/a_112_119#
+ prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_35/a_230_79# prbs_generator_syn_11/m3_13600_4091#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_23/a_1226_296# prbs_generator_syn_11/sky130_fd_sc_hs__nand2_1_39/a_117_74#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_29/a_27_74# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_5/a_437_503#
+ prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_17/a_293_74# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_41/a_1178_124#
+ prbs_generator_syn_11/sky130_fd_sc_hs__or2_1_1/a_152_368# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_59/a_1178_124#
+ prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_61/a_293_74# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_47/a_206_368#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_39/a_651_503# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_49/a_696_458#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_15/a_735_102# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_32/a_1034_424#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_73/a_1226_296# prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_27/a_222_392#
+ prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_41/a_112_119# prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_31/a_52_123#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_49/a_1034_424# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_29/a_1141_508#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_21/a_1226_296# prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_39/a_230_79#
+ prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_23/a_138_385# prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_51/a_230_79#
+ prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_45/a_132_392# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_37/a_206_368#
+ prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_65/a_293_74# prbs_generator_syn_11/sky130_fd_sc_hs__nand2_1_53/a_117_74#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_47/a_437_503# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_29/a_651_503#
+ prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_31/a_293_74# prbs_generator_syn_11/sky130_fd_sc_hs__nand2_1_21/a_117_74#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_69/a_544_485# prbs_generator_syn_11/sky130_fd_sc_hs__clkbuf_16_1/a_114_74#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_45/a_735_102# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_13/a_27_74#
+ prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_31/a_112_119# prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_57/a_222_392#
+ prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_35/a_52_123# prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_21/a_376_368#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_7/a_544_485# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_57/a_1178_124#
+ prbs_generator_syn_11/m3_13600_6043# prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_13/a_138_385#
+ prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_51/a_138_385# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_5/a_1141_508#
+ prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_3/a_376_368# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_27/a_206_368#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_65/a_206_368# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_37/a_437_503#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_19/a_651_503# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_57/a_651_503#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_59/a_544_485# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_71/a_1226_296#
+ prbs_generator_syn_11/sky130_fd_sc_hs__nand2_1_25/a_117_74# prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_61/a_112_119#
+ prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_47/a_222_392# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_27/a_1141_508#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_53/a_27_74# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_4/a_206_368#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_39/a_1226_296# prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_11/a_376_368#
+ prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_39/a_52_123# prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_41/a_138_385#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_4/a_1141_508# prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_25/a_132_392#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_17/a_206_368# prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_41/A
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_55/a_206_368# prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_51/a_52_123#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_27/a_437_503# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_65/a_437_503#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_49/a_544_485# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_63/a_735_102#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_47/a_1034_424# prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_50/a_112_119#
+ prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_37/a_222_392# prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_59/a_230_79#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_25/a_1141_508# prbs_generator_syn_11/sky130_fd_sc_hs__nor2b_1_4/a_27_112#
+ prbs_generator_syn_11/sky130_fd_sc_hs__sdlclkp_2_1/a_685_81# prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_1/a_132_392#
+ prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_39/a_293_74# prbs_generator_syn_11/sky130_fd_sc_hs__nand2_1_29/a_117_74#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_4/a_437_503# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_55/a_1178_124#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_21/a_27_74# prbs_generator_syn_11/m3_13600_12875#
+ prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_50/a_293_74# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_1/a_735_102#
+ prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_31/a_138_385# prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_15/a_132_392#
+ prbs_generator_syn_11/sky130_fd_sc_hs__nand2_1_1/a_117_74# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_17/a_437_503#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_55/a_437_503# prbs_generator_syn
Xprbs_generator_syn_21 prbs_generator_syn_31/clk prbs_generator_syn_31/rst prbs_generator_syn_21/cke
+ sky130_fd_sc_hs__conb_1_223/LO sky130_fd_sc_hs__conb_1_223/LO sky130_fd_sc_hs__conb_1_223/LO
+ prbs_generator_syn_25/eqn[1] prbs_generator_syn_25/eqn[1] prbs_generator_syn_25/eqn[1]
+ prbs_generator_syn_25/eqn[1] prbs_generator_syn_25/eqn[1] sky130_fd_sc_hs__conb_1_223/LO
+ sky130_fd_sc_hs__conb_1_223/LO sky130_fd_sc_hs__conb_1_223/LO prbs_generator_syn_21/eqn[31]
+ prbs_generator_syn_25/eqn[9] sky130_fd_sc_hs__conb_1_215/HI prbs_generator_syn_25/eqn[9]
+ sky130_fd_sc_hs__conb_1_215/HI prbs_generator_syn_25/eqn[9] prbs_generator_syn_21/cke
+ prbs_generator_syn_21/eqn[0] prbs_generator_syn_23/eqn[20] prbs_generator_syn_23/eqn[22]
+ prbs_generator_syn_23/eqn[20] prbs_generator_syn_23/eqn[22] sky130_fd_sc_hs__conb_1_181/HI
+ sky130_fd_sc_hs__conb_1_181/HI prbs_generator_syn_23/eqn[28] prbs_generator_syn_23/eqn[28]
+ sky130_fd_sc_hs__conb_1_227/HI sky130_fd_sc_hs__conb_1_227/HI sky130_fd_sc_hs__conb_1_227/HI
+ sky130_fd_sc_hs__conb_1_227/HI sky130_fd_sc_hs__conb_1_227/HI prbs_generator_syn_21/eqn[31]
+ prbs_generator_syn_21/eqn[30] prbs_generator_syn_21/eqn[30] prbs_generator_syn_21/eqn[30]
+ prbs_generator_syn_21/eqn[30] prbs_generator_syn_21/eqn[30] prbs_generator_syn_21/eqn[30]
+ prbs_generator_syn_21/eqn[30] prbs_generator_syn_21/eqn[30] prbs_generator_syn_21/eqn[22]
+ prbs_generator_syn_21/eqn[22] prbs_generator_syn_21/eqn[20] prbs_generator_syn_21/eqn[22]
+ prbs_generator_syn_21/eqn[22] prbs_generator_syn_21/eqn[22] prbs_generator_syn_21/eqn[22]
+ prbs_generator_syn_21/eqn[22] prbs_generator_syn_21/eqn[22] prbs_generator_syn_21/eqn[9]
+ prbs_generator_syn_21/eqn[9] prbs_generator_syn_21/eqn[9] prbs_generator_syn_21/eqn[9]
+ prbs_generator_syn_21/eqn[9] prbs_generator_syn_21/eqn[8] prbs_generator_syn_21/eqn[8]
+ prbs_generator_syn_21/eqn[8] prbs_generator_syn_21/eqn[8] prbs_generator_syn_21/eqn[8]
+ prbs_generator_syn_21/eqn[8] prbs_generator_syn_21/eqn[8] prbs_generator_syn_21/eqn[1]
+ prbs_generator_syn_21/eqn[0] prbs_generator_syn_31/inj_err prbs_generator_syn_21/eqn[31]
+ prbs_generator_syn_21/eqn[31] prbs_generator_syn_21/out DVSS: DVDD: prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_1/a_293_74#
+ prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_15/X prbs_generator_syn_21/sky130_fd_sc_hs__nand2_1_35/B
+ prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_51/Y prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_9/A
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_9/CLK prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_47/a_27_74#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_37/a_1226_296# prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_3/B
+ prbs_generator_syn_21/sky130_fd_sc_hs__nor2b_1_7/a_27_112# prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_29/B
+ prbs_generator_syn_21/sky130_fd_sc_hs__sdlclkp_2_1/a_580_74# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_1/a_1141_508#
+ prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_5/Y prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_41/a_230_79#
+ prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_61/a_138_385# prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_43/a_132_392#
+ prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_3/a_222_392# prbs_generator_syn_21/sky130_fd_sc_hs__nor2b_1_9/a_27_112#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_61/a_27_74# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_35/a_206_368#
+ prbs_generator_syn_21/sky130_fd_sc_hs__nand2_2_3/Y prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_25/B
+ prbs_generator_syn_21/sky130_fd_sc_hs__nand2_1_11/a_117_74# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_67/a_651_503#
+ prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_45/X prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_39/a_696_458#
+ prbs_generator_syn_21/sky130_fd_sc_hs__sdlclkp_2_1/a_1198_74# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_45/a_1034_424#
+ prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_17/a_222_392# prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_55/a_222_392#
+ prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_53/Y prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_35/A
+ prbs_generator_syn_21/m3_13600_1651# prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_59/a_52_123#
+ prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_5/a_293_74# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_35/a_1226_296#
+ prbs_generator_syn_21/sky130_fd_sc_hs__nand2_1_51/B prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_5/a_651_503#
+ prbs_generator_syn_21/sky130_fd_sc_hs__nand2_1_21/B prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_8/a_27_74#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_15/a_27_74# prbs_generator_syn_21/sky130_fd_sc_hs__and2b_2_1/X
+ prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_13/X prbs_generator_syn_21/sky130_fd_sc_hs__nand2_2_3/a_27_74#
+ prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_50/a_138_385# prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_33/a_132_392#
+ prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_1/a_376_368# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_25/a_206_368#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_35/a_437_503# prbs_generator_syn_21/sky130_fd_sc_hs__sdlclkp_2_1/a_708_451#
+ prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_45/a_230_79# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_29/a_696_458#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_32/a_27_74# prbs_generator_syn_21/sky130_fd_sc_hs__nor2b_1_4/Y
+ prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_59/a_293_74# prbs_generator_syn_21/sky130_fd_sc_hs__nand2_1_47/a_117_74#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_73/a_735_102# prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_21/a_112_119#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_23/a_1141_508# prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_25/a_293_74#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_7/Q prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_3/a_112_119#
+ prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_35/B prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_51/X
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_53/a_1178_124# prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_23/a_132_392#
+ prbs_generator_syn_21/sky130_fd_sc_hs__nand2_1_3/B prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_15/a_206_368#
+ prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_63/a_132_392# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_55/a_27_74#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_25/a_437_503# prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_41/a_52_123#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_47/a_651_503# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_73/a_1141_508#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_19/a_696_458# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_57/a_696_458#
+ prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_7/X prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_43/a_1034_424#
+ prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_55/A prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_11/a_112_119#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_21/a_1141_508# prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_35/a_222_392#
+ prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_49/a_230_79# prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_67/Y
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_71/a_27_74# prbs_generator_syn_21/sky130_fd_sc_hs__nand2_1_33/B
+ prbs_generator_syn_21/sky130_fd_sc_hs__conb_1_1/LO prbs_generator_syn_21/sky130_fd_sc_hs__nand2_1_19/a_117_74#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_51/a_1178_124# prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_33/X
+ prbs_generator_syn_21/sky130_fd_sc_hs__nand2_1_29/B prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_41/Y
+ prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_53/a_132_392# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_45/a_206_368#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_15/a_437_503# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_37/a_651_503#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_39/a_544_485# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_53/a_735_102#
+ prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_45/a_52_123# prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_1/B
+ prbs_generator_syn_21/sky130_fd_sc_hs__nand2_2_3/B prbs_generator_syn_21/sky130_fd_sc_hs__clkbuf_16_1/A
+ prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_21/X prbs_generator_syn_21/sky130_fd_sc_hs__nand2_1_25/B
+ prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_39/a_376_368# prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_63/X
+ prbs_generator_syn_21/m3_13600_3481# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_69/a_1178_124#
+ prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_21/a_138_385# prbs_generator_syn_21/sky130_fd_sc_hs__nor2b_1_8/Y
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_19/a_1178_124# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_49/a_27_74#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_45/a_437_503# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_27/a_651_503#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_71/a_1141_508# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_65/a_651_503#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_29/a_544_485# prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_3/a_138_385#
+ prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_55/X prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_43/a_735_102#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_41/a_1034_424# prbs_generator_syn_21/sky130_fd_sc_hs__nand2_1_9/B
+ prbs_generator_syn_21/sky130_fd_sc_hs__nor2b_1_9/Y prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_59/a_1034_424#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_39/a_1141_508# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_33/a_1226_296#
+ prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_49/a_52_123# prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_47/Y
+ prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_43/Y prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_4/a_651_503#
+ prbs_generator_syn_21/sky130_fd_sc_hs__nand2_1_49/B prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_19/A
+ prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_11/a_138_385# prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_5/X
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_63/a_206_368# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_17/a_651_503#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_19/a_544_485# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_55/a_651_503#
+ prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_9/Y prbs_generator_syn_21/sky130_fd_sc_hs__nand2_1_17/B
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_57/a_544_485# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_67/a_696_458#
+ prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_35/X prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_19/a_27_74#
+ prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_45/a_222_392# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_32/a_1226_296#
+ prbs_generator_syn_21/sky130_fd_sc_hs__nand2_1_43/B prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_25/A
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_1/a_206_368# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_49/a_1226_296#
+ prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_1/a_112_119# prbs_generator_syn_21/sky130_fd_sc_hs__or2_1_1/X
+ prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_59/a_376_368# prbs_generator_syn_21/sky130_fd_sc_hs__nand2_1_19/B
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_5/a_696_458# prbs_generator_syn_21/sky130_fd_sc_hs__nor2b_1_1/Y
+ prbs_generator_syn_21/sky130_fd_sc_hs__nor2b_1_5/a_278_368# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_17/a_1178_124#
+ prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_39/X prbs_generator_syn_21/m3_13600_5433#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_63/a_437_503# prbs_generator_syn_21/sky130_fd_sc_hs__nand2_2_5/B
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_23/a_735_102# prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_53/A
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_61/a_735_102# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_57/a_1034_424#
+ prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_63/B prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_37/a_1141_508#
+ prbs_generator_syn_21/sky130_fd_sc_hs__nand2_1_47/B prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_29/X
+ prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_65/Y prbs_generator_syn_21/m3_13600_4701#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_1/a_437_503# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_67/a_1178_124#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_9/a_735_102# prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_13/a_132_392#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_15/a_1178_124# prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_15/A
+ prbs_generator_syn_21/sky130_fd_sc_hs__nand2_1_1/B prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_43/B
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_35/a_651_503# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_8/D
+ prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_29/A prbs_generator_syn_21/sky130_fd_sc_hs__nand2_1_7/B
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_13/a_735_102# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_47/a_696_458#
+ prbs_generator_syn_21/sky130_fd_sc_hs__nand2_1_31/B prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_51/a_735_102#
+ prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_59/X prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_35/a_1141_508#
+ prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_25/a_222_392# prbs_generator_syn_21/sky130_fd_sc_hs__sdlclkp_2_1/a_288_48#
+ prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_55/B prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_17/B
+ prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_43/A prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_7/A
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_65/a_1178_124# prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_59/Y
+ prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_41/X prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_21/a_230_79#
+ prbs_generator_syn_21/sky130_fd_sc_hs__nand2_1_57/a_117_74# prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_1/a_222_392#
+ prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_19/B prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_35/a_293_74#
+ prbs_generator_syn_21/sky130_fd_sc_hs__nand2_1_23/a_117_74# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_73/a_206_368#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_25/a_651_503# prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_1/a_138_385#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_37/a_696_458# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_67/a_544_485#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_43/a_27_74# prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_9/X
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_55/a_1034_424# prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_39/a_112_119#
+ prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_15/a_222_392# prbs_generator_syn_21/sky130_fd_sc_hs__conb_1_1/HI
+ prbs_generator_syn_21/sky130_fd_sc_hs__nand2_1_23/B prbs_generator_syn_21/sky130_fd_sc_hs__nand2_1_53/B
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_9/a_1178_124# prbs_generator_syn_21/sky130_fd_sc_hs__nor2b_1_4/A
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_47/a_1226_296# prbs_generator_syn_21/m3_13600_11045#
+ prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_17/X prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_29/a_376_368#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_5/a_544_485# prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_3/X
+ prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_31/a_132_392# prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_61/A
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_15/a_651_503# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_73/a_437_503#
+ prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_25/a_230_79# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_27/a_696_458#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_65/a_696_458# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_33/a_735_102#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_71/a_735_102# prbs_generator_syn_21/m3_13600_7263#
+ prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_43/a_222_392# prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_50/Y
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_8/a_1178_124# prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_53/B
+ prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_19/a_376_368# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_63/a_1178_124#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_4/a_696_458# prbs_generator_syn_21/sky130_fd_sc_hs__nor2b_1_4/a_278_368#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_13/a_1178_124# prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_61/a_132_392#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_53/a_206_368# prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_21/a_52_123#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_45/a_651_503# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_17/a_696_458#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_47/a_544_485# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_55/a_696_458#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_21/a_735_102# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_37/a_27_74#
+ prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_61/B prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_61/X
+ prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_59/a_112_119# prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_31/A
+ prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_33/a_222_392# prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_29/a_230_79#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_45/a_1226_296# prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_9/a_132_392#
+ prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_5/A prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_57/Y
+ prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_31/X prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_51/a_27_74#
+ prbs_generator_syn_21/sky130_fd_sc_hs__nor2b_1_8/a_27_112# prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_47/a_376_368#
+ prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_53/a_293_74# prbs_generator_syn_21/sky130_fd_sc_hs__nand2_1_43/a_117_74#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_8/a_735_102# prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_21/a_293_74#
+ prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_39/a_138_385# prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_63/Y
+ prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_51/a_132_392# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_43/a_206_368#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_53/a_437_503# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_37/a_544_485#
+ prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_57/X prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_53/a_1034_424#
+ prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_25/a_52_123# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_33/a_1141_508#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_63/Q prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_23/a_222_392#
+ prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_63/a_222_392# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_7/a_1178_124#
+ prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_53/X prbs_generator_syn_21/sky130_fd_sc_hs__nand2_2_5/Y
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_61/a_1178_124# prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_1/a_230_79#
+ prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_43/a_230_79# prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_11/a_230_79#
+ prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_41/a_132_392# prbs_generator_syn_21/sky130_fd_sc_hs__nand2_1_13/a_117_74#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_43/a_437_503# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_27/a_544_485#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_63/a_651_503# prbs_generator_syn_21/sky130_fd_sc_hs__nand2_1_7/a_117_74#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_35/a_696_458# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_65/a_544_485#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_51/a_1034_424# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_41/a_735_102#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_32/a_1141_508# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_49/a_1141_508#
+ prbs_generator_syn_21/sky130_fd_sc_hs__nand2_1_55/B prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_53/a_222_392#
+ prbs_generator_syn_21/sky130_fd_sc_hs__sdlclkp_2_1/a_114_112# prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_9/a_293_74#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_43/a_1226_296# prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_29/a_52_123#
+ prbs_generator_syn_21/sky130_fd_sc_hs__nand2_1_37/B prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_1/a_651_503#
+ prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_27/a_376_368# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_4/a_544_485#
+ prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_67/a_376_368# prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_27/X
+ prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_1/X prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_59/a_138_385#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_29/a_1178_124# prbs_generator_syn_21/m3_13600_2871#
+ prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_5/a_230_79# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_23/a_206_368#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_61/a_206_368# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_17/a_544_485#
+ prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_15/a_230_79# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_25/a_696_458#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_55/a_544_485# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_32/a_735_102#
+ prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_29/a_293_74# prbs_generator_syn_21/sky130_fd_sc_hs__nand2_1_17/a_117_74#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_69/a_1034_424# prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_29/a_112_119#
+ prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_37/X prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_31/B
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_19/a_1034_424# prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_33/A
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_9/a_206_368# prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_57/a_376_368#
+ prbs_generator_syn_21/sky130_fd_sc_hs__sdlclkp_2_1/a_706_317# prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_11/B
+ prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_1/a_52_123# prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_39/B
+ prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_21/a_132_392# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_13/a_206_368#
+ prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_43/a_52_123# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_51/a_206_368#
+ prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_47/X prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_23/a_437_503#
+ prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_11/a_52_123# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_61/a_437_503#
+ prbs_generator_syn_21/sky130_fd_sc_hs__nor2b_1_7/Y prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_51/A
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_15/a_696_458# prbs_generator_syn_21/sky130_fd_sc_hs__nor2b_1_5/Y
+ prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_9/a_230_79# prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_25/X
+ prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_19/a_112_119# prbs_generator_syn_21/sky130_fd_sc_hs__nand2_1_45/B
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_5/a_1178_124# prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_19/a_230_79#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_41/a_1226_296# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_59/a_1226_296#
+ prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_63/a_230_79# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_51/Q
+ prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_7/a_132_392# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_9/a_437_503#
+ prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_46/a_376_368# prbs_generator_syn_21/sky130_fd_sc_hs__nand2_1_33/a_117_74#
+ prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_11/a_293_74# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_27/a_1178_124#
+ prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_11/a_132_392# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_13/a_437_503#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_51/a_437_503# prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_5/a_52_123#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_35/a_544_485# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_73/a_651_503#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_45/a_696_458# prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_15/a_52_123#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_47/a_1141_508# prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_47/a_112_119#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_4/a_1178_124# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_17/a_1034_424#
+ prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_23/B prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_37/a_376_368#
+ prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_15/B prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_7/Y
+ prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_29/a_138_385# prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_33/a_230_79#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_25/a_1178_124# prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_47/a_293_74#
+ prbs_generator_syn_21/sky130_fd_sc_hs__nand2_1_37/a_117_74# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_33/a_206_368#
+ prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_15/a_293_74# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_71/a_206_368#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_25/a_544_485# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_67/a_1034_424#
+ prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_13/a_222_392# prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_9/a_52_123#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_15/a_1034_424# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_57/a_1226_296#
+ prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_19/a_52_123# prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_23/X
+ prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_63/a_52_123# prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_19/a_138_385#
+ prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_9/a_376_368# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_21/a_206_368#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_33/a_437_503# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_71/a_437_503#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_53/a_651_503# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_15/a_544_485#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_63/a_696_458# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_65/a_1034_424#
+ prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_19/a_293_74# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_45/a_1141_508#
+ prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_27/a_112_119# prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_67/a_112_119#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_1/a_1178_124# prbs_generator_syn_21/sky130_fd_sc_hs__conb_1_1/a_21_290#
+ prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_63/a_293_74# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_8/a_206_368#
+ prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_17/a_376_368# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_63/a_27_74#
+ prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_21/A prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_55/a_376_368#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_1/a_696_458# prbs_generator_syn_21/sky130_fd_sc_hs__nor2b_1_1/a_278_368#
+ prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_47/a_138_385# prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_33/a_52_123#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_9/a_1034_424# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_21/a_437_503#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_1/a_27_74# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_43/a_651_503#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_1/Q prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_45/a_544_485#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_69/a_735_102# prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_57/a_112_119#
+ prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_31/a_222_392# prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_13/A
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_55/a_1226_296# prbs_generator_syn_21/sky130_fd_sc_hs__nand2_2_5/a_27_74#
+ prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_53/a_230_79# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_8/a_437_503#
+ prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_67/a_293_74# prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_33/a_293_74#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_7/a_735_102# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_23/a_1178_124#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_41/a_206_368# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_8/a_1034_424#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_63/a_1034_424# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_59/a_735_102#
+ prbs_generator_syn_21/sky130_fd_sc_hs__nand2_1_5/B prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_43/a_1141_508#
+ prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_46/a_112_119# prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_61/a_222_392#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_13/a_1034_424# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_73/a_1178_124#
+ prbs_generator_syn_21/sky130_fd_sc_hs__nand2_1_27/B prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_13/B
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_57/a_27_74# prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_57/a_230_79#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_21/a_1178_124# prbs_generator_syn_21/sky130_fd_sc_hs__nor2b_1_1/a_27_112#
+ prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_27/a_138_385# prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_23/a_230_79#
+ prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_67/a_138_385# prbs_generator_syn_21/sky130_fd_sc_hs__nand2_1_41/B
+ prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_9/a_222_392# prbs_generator_syn_21/sky130_fd_sc_hs__nand2_1_27/a_117_74#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_32/a_206_368# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_23/a_651_503#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_41/a_437_503# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_73/a_27_74#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_61/a_651_503# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_63/a_544_485#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_49/a_735_102# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_73/a_696_458#
+ prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_37/a_112_119# prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_51/a_222_392#
+ prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_43/X prbs_generator_syn_21/sky130_fd_sc_hs__nand2_2_1/B
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_9/a_651_503# prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_53/a_52_123#
+ prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_49/X prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_25/a_376_368#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_1/a_544_485# prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_65/a_376_368#
+ prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_57/a_138_385# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_27/a_27_74#
+ prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_39/a_132_392# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_7/a_1034_424#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_13/a_651_503# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_32/a_437_503#
+ prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_27/a_230_79# prbs_generator_syn_21/m3_13600_12265#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_51/a_651_503# prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_59/B
+ prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_47/A prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_61/a_1034_424#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_41/a_1141_508# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_59/a_1141_508#
+ prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_41/a_222_392# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_53/a_1226_296#
+ prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_3/A prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_71/a_1178_124#
+ prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_9/a_112_119# prbs_generator_syn_21/sky130_fd_sc_hs__nand2_1_3/a_117_74#
+ prbs_generator_syn_21/m3_13600_8483# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_39/a_1178_124#
+ prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_57/a_52_123# prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_46/a_138_385#
+ prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_23/a_52_123# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_67/a_27_74#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_53/a_696_458# prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_17/a_112_119#
+ prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_11/A prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_55/a_112_119#
+ prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_1/A prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_51/a_1226_296#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_29/a_1034_424# prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_59/A
+ prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_23/A prbs_generator_syn_21/sky130_fd_sc_hs__nand2_1_39/B
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_5/a_27_74# prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_57/a_293_74#
+ prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_37/a_138_385# prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_59/a_132_392#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_33/a_651_503# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_71/a_651_503#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_43/a_696_458# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_73/a_544_485#
+ prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_27/a_52_123# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_57/a_1141_508#
+ prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_21/a_222_392# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_35/a_27_74#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_69/a_1226_296# prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_37/B
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_19/a_1226_296# prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_35/a_376_368#
+ prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_47/a_230_79# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_37/a_1178_124#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_5/a_1034_424# prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_49/a_132_392#
+ prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_7/a_222_392# prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_27/a_293_74#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_21/a_651_503# prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_9/a_138_385#
+ prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_11/a_222_392# prbs_generator_syn_21/m3_13600_14095#
+ prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_50/A prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_27/a_1034_424#
+ prbs_generator_syn_21/sky130_fd_sc_hs__nand2_1_13/B prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_8/a_651_503#
+ prbs_generator_syn_21/m3_13600_9703# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_35/a_1178_124#
+ prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_17/a_138_385# prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_55/a_138_385#
+ prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_7/a_230_79# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_4/a_1034_424#
+ prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_7/a_376_368# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_69/a_206_368#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_23/a_696_458# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_53/a_544_485#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_39/a_735_102# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_61/a_696_458#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_55/a_1141_508# prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_25/a_112_119#
+ prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_65/a_112_119# prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_43/a_293_74#
+ prbs_generator_syn_21/sky130_fd_sc_hs__nand2_1_57/B prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_25/a_1034_424#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_7/a_206_368# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_17/a_1226_296#
+ prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_15/a_376_368# prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_53/a_376_368#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_9/a_696_458# prbs_generator_syn_21/m3_13600_431#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_45/a_27_74# prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_47/a_52_123#
+ prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_29/a_132_392# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_59/a_206_368#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_69/a_437_503# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_41/a_651_503#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_43/a_544_485# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_13/a_696_458#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_29/a_735_102# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_51/a_696_458#
+ prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_61/Y prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_67/a_1226_296#
+ prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_5/a_132_392# prbs_generator_syn_21/sky130_fd_sc_hs__and2b_2_1/a_198_48#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_7/a_437_503# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_15/a_1226_296#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_69/a_27_74# prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_46/a_293_74#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_1/a_1034_424# prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_19/a_132_392#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_49/a_206_368# prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_7/a_52_123#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_59/a_437_503# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_32/a_651_503#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_7/a_27_74# prbs_generator_syn_21/sky130_fd_sc_hs__nand2_2_1/a_27_74#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_19/a_735_102# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_57/a_735_102#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_65/a_1226_296# prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_37/A
+ prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_33/a_376_368# prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_37/a_230_79#
+ prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_25/a_138_385# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_39/a_27_74#
+ prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_65/a_138_385# prbs_generator_syn_21/sky130_fd_sc_hs__nor2b_1_9/a_278_368#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_49/a_437_503# prbs_generator_syn_21/sky130_fd_sc_hs__and2b_2_1/a_505_74#
+ prbs_generator_syn_21/sky130_fd_sc_hs__nand2_1_51/a_117_74# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_23/a_544_485#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_33/a_696_458# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_61/a_544_485#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_9/a_1226_296# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_53/a_1141_508#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_71/a_696_458# prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_35/a_112_119#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_23/a_1034_424# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_9/a_544_485#
+ prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_63/a_376_368# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_33/a_1178_124#
+ prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_5/a_376_368# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_13/a_544_485#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_73/a_1034_424# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_21/a_696_458#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_51/a_544_485# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_8/a_1226_296#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_51/a_1141_508# prbs_generator_syn_21/sky130_fd_sc_hs__nand2_1_55/a_117_74#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_21/a_1034_424# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_63/a_1226_296#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_23/a_27_74# prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_7/a_112_119#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_13/a_1226_296# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_8/a_696_458#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_32/a_1178_124# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_49/a_1178_124#
+ prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_37/a_52_123# prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_27/a_132_392#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_71/Q prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_67/a_735_102#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_69/a_1141_508# prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_15/a_112_119#
+ prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_53/a_112_119# prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_39/a_222_392#
+ prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_55/a_230_79# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_19/a_1141_508#
+ prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_37/a_293_74# prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_43/a_376_368#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_5/a_735_102# prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_35/a_138_385#
+ prbs_generator_syn_21/sky130_fd_sc_hs__sdlclkp_2_1/a_114_424# prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_57/a_132_392#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_71/a_1034_424# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_7/a_1226_296#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_33/a_544_485# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_41/a_696_458#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_71/a_544_485# prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_21/B
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_61/a_1226_296# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_39/a_1034_424#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_17/a_27_74# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_9/a_27_74#
+ prbs_generator_syn_21/sky130_fd_sc_hs__nor2b_1_5/a_27_112# prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_47/a_132_392#
+ prbs_generator_syn_21/sky130_fd_sc_hs__nor2b_1_8/a_278_368# prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_9/B
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_39/a_206_368# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_33/a_27_74#
+ prbs_generator_syn_21/sky130_fd_sc_hs__nand2_1_41/a_117_74# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_69/a_651_503#
+ prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_51/a_293_74# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_21/a_544_485#
+ prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_7/a_138_385# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_32/a_696_458#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_47/a_735_102# prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_33/a_112_119#
+ prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_59/a_222_392# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_17/a_1141_508#
+ prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_55/a_52_123# prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_3/a_293_74#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_7/a_651_503# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_29/a_1226_296#
+ prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_23/a_376_368# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_8/a_544_485#
+ prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_47/B prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_47/a_1178_124#
+ prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_15/a_138_385# prbs_generator_syn_21/sky130_fd_sc_hs__sdlclkp_2_1/a_1195_374#
+ prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_53/a_138_385# prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_37/a_132_392#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_29/a_206_368# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_39/a_437_503#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_59/a_651_503# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_37/a_735_102#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_67/a_1141_508# prbs_generator_syn_21/sky130_fd_sc_hs__and2b_2_1/a_27_74#
+ prbs_generator_syn_21/sky130_fd_sc_hs__conb_1_1/a_165_290# prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_55/a_293_74#
+ prbs_generator_syn_21/sky130_fd_sc_hs__nand2_1_45/a_117_74# prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_63/a_112_119#
+ prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_49/a_222_392# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_37/a_1034_424#
+ prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_23/a_293_74# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_15/a_1141_508#
+ prbs_generator_syn_21/sky130_fd_sc_hs__nand2_1_5/a_117_74# prbs_generator_syn_21/m3_13600_13485#
+ prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_5/a_112_119# prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_13/a_376_368#
+ prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_51/a_376_368# prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_7/a_293_74#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_19/a_206_368# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_57/a_206_368#
+ prbs_generator_syn_21/sky130_fd_sc_hs__sdlclkp_2_1/a_318_74# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_29/a_437_503#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_49/a_651_503# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_25/a_27_74#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_5/a_1226_296# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_41/a_544_485#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_27/a_735_102# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_65/a_1141_508#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_65/a_735_102# prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_3/a_230_79#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_35/a_1034_424# prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_13/a_230_79#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_41/a_27_74# prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_3/a_132_392#
+ prbs_generator_syn_21/sky130_fd_sc_hs__nand2_1_49/a_117_74# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_27/a_1226_296#
+ prbs_generator_syn_21/sky130_fd_sc_hs__nand2_1_15/a_117_74# prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_41/a_376_368#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_45/a_1178_124# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_4/a_735_102#
+ prbs_generator_syn_21/sky130_fd_sc_hs__nand2_1_9/a_117_74# prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_33/a_138_385#
+ prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_17/a_132_392# prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_55/a_132_392#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_9/a_1141_508# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_19/a_437_503#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_57/a_437_503# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_4/a_1226_296#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_32/a_544_485# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_17/a_735_102#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_55/a_735_102# prbs_generator_syn_21/m3_13600_2261#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_65/a_27_74# prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_29/a_222_392#
+ prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_43/a_112_119# prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_19/X
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_25/a_1226_296# prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_31/a_376_368#
+ prbs_generator_syn_21/sky130_fd_sc_hs__or2_1_1/a_63_368# prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_17/a_230_79#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_4/a_27_74# prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_61/a_230_79#
+ prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_63/a_138_385# prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_5/a_222_392#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_8/a_1141_508# prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_41/a_293_74#
+ prbs_generator_syn_21/sky130_fd_sc_hs__nand2_1_31/a_117_74# prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_5/a_138_385#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_63/a_1141_508# prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_19/a_222_392#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_13/a_1141_508# prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_3/a_52_123#
+ prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_13/a_52_123# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_43/a_1178_124#
+ prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_61/a_376_368# prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_35/a_132_392#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_67/a_206_368# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_1/a_1226_296#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_69/a_696_458# prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_31/a_230_79#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_35/a_735_102# prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_23/a_112_119#
+ prbs_generator_syn_21/sky130_fd_sc_hs__nand2_1_35/a_117_74# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_59/a_27_74#
+ prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_13/a_293_74# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_5/a_206_368#
+ prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_50/a_376_368# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_7/a_696_458#
+ prbs_generator_syn_21/sky130_fd_sc_hs__nor2b_1_7/a_278_368# prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_17/a_52_123#
+ prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_43/a_138_385# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_7/a_1141_508#
+ prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_61/a_52_123# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_67/a_437_503#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_61/a_1141_508# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_25/a_735_102#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_59/a_696_458# prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_13/a_112_119#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_33/a_1034_424# prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_51/a_112_119#
+ prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_35/a_230_79# prbs_generator_syn_21/m3_13600_4091#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_23/a_1226_296# prbs_generator_syn_21/sky130_fd_sc_hs__nand2_1_39/a_117_74#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_29/a_27_74# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_5/a_437_503#
+ prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_17/a_293_74# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_41/a_1178_124#
+ prbs_generator_syn_21/sky130_fd_sc_hs__or2_1_1/a_152_368# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_59/a_1178_124#
+ prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_61/a_293_74# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_47/a_206_368#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_39/a_651_503# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_49/a_696_458#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_15/a_735_102# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_32/a_1034_424#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_73/a_1226_296# prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_27/a_222_392#
+ prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_41/a_112_119# prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_31/a_52_123#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_49/a_1034_424# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_29/a_1141_508#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_21/a_1226_296# prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_39/a_230_79#
+ prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_23/a_138_385# prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_51/a_230_79#
+ prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_45/a_132_392# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_37/a_206_368#
+ prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_65/a_293_74# prbs_generator_syn_21/sky130_fd_sc_hs__nand2_1_53/a_117_74#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_47/a_437_503# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_29/a_651_503#
+ prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_31/a_293_74# prbs_generator_syn_21/sky130_fd_sc_hs__nand2_1_21/a_117_74#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_69/a_544_485# prbs_generator_syn_21/sky130_fd_sc_hs__clkbuf_16_1/a_114_74#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_45/a_735_102# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_13/a_27_74#
+ prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_31/a_112_119# prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_57/a_222_392#
+ prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_35/a_52_123# prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_21/a_376_368#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_7/a_544_485# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_57/a_1178_124#
+ prbs_generator_syn_21/m3_13600_6043# prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_13/a_138_385#
+ prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_51/a_138_385# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_5/a_1141_508#
+ prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_3/a_376_368# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_27/a_206_368#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_65/a_206_368# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_37/a_437_503#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_19/a_651_503# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_57/a_651_503#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_59/a_544_485# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_71/a_1226_296#
+ prbs_generator_syn_21/sky130_fd_sc_hs__nand2_1_25/a_117_74# prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_61/a_112_119#
+ prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_47/a_222_392# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_27/a_1141_508#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_53/a_27_74# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_4/a_206_368#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_39/a_1226_296# prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_11/a_376_368#
+ prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_39/a_52_123# prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_41/a_138_385#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_4/a_1141_508# prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_25/a_132_392#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_17/a_206_368# prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_41/A
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_55/a_206_368# prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_51/a_52_123#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_27/a_437_503# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_65/a_437_503#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_49/a_544_485# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_63/a_735_102#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_47/a_1034_424# prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_50/a_112_119#
+ prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_37/a_222_392# prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_59/a_230_79#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_25/a_1141_508# prbs_generator_syn_21/sky130_fd_sc_hs__nor2b_1_4/a_27_112#
+ prbs_generator_syn_21/sky130_fd_sc_hs__sdlclkp_2_1/a_685_81# prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_1/a_132_392#
+ prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_39/a_293_74# prbs_generator_syn_21/sky130_fd_sc_hs__nand2_1_29/a_117_74#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_4/a_437_503# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_55/a_1178_124#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_21/a_27_74# prbs_generator_syn_21/m3_13600_12875#
+ prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_50/a_293_74# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_1/a_735_102#
+ prbs_generator_syn_21/sky130_fd_sc_hs__xnor2_1_31/a_138_385# prbs_generator_syn_21/sky130_fd_sc_hs__a22o_1_15/a_132_392#
+ prbs_generator_syn_21/sky130_fd_sc_hs__nand2_1_1/a_117_74# prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_17/a_437_503#
+ prbs_generator_syn_21/sky130_fd_sc_hs__dfxtp_4_55/a_437_503# prbs_generator_syn
Xsky130_fd_sc_hs__conb_1_1 DVSS: DVDD: DVDD: DVSS: prbs_generator_syn_1/eqn[9] sky130_fd_sc_hs__conb_1_1/HI
+ sky130_fd_sc_hs__conb_1_1/a_165_290# sky130_fd_sc_hs__conb_1_1/a_21_290# sky130_fd_sc_hs__conb_1
Xsky130_fd_sc_hs__buf_2_130 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__buf_2_131/A sky130_fd_sc_hs__buf_2_131/X
+ sky130_fd_sc_hs__buf_2_131/a_21_260# sky130_fd_sc_hs__buf_2
Xsky130_fd_sc_hs__buf_2_141 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__buf_2_37/X sky130_fd_sc_hs__buf_2_141/X
+ sky130_fd_sc_hs__buf_2_141/a_21_260# sky130_fd_sc_hs__buf_2
Xsky130_fd_sc_hs__buf_2_152 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__buf_2_153/A sky130_fd_sc_hs__buf_2_153/X
+ sky130_fd_sc_hs__buf_2_153/a_21_260# sky130_fd_sc_hs__buf_2
Xsky130_fd_sc_hs__buf_2_163 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__buf_2_67/X sky130_fd_sc_hs__buf_2_163/X
+ sky130_fd_sc_hs__buf_2_163/a_21_260# sky130_fd_sc_hs__buf_2
Xsky130_fd_sc_hs__einvp_2_20 DVSS: DVDD: DVDD: DVSS: dout_n sky130_fd_sc_hs__buf_8_1/A
+ sky130_fd_sc_hs__dlrtp_1_21/Q sky130_fd_sc_hs__einvp_2_21/a_263_323# sky130_fd_sc_hs__einvp_2_21/a_36_74#
+ sky130_fd_sc_hs__einvp_2_21/a_27_368# sky130_fd_sc_hs__einvp_2
Xsky130_fd_sc_hs__einvp_2_31 DVSS: DVDD: DVDD: DVSS: dout_n sky130_fd_sc_hs__buf_8_1/A
+ sky130_fd_sc_hs__dlrtp_1_27/Q sky130_fd_sc_hs__einvp_2_31/a_263_323# sky130_fd_sc_hs__einvp_2_31/a_36_74#
+ sky130_fd_sc_hs__einvp_2_31/a_27_368# sky130_fd_sc_hs__einvp_2
Xsky130_fd_sc_hs__einvp_2_42 DVSS: DVDD: DVDD: DVSS: dout_n sky130_fd_sc_hs__buf_8_1/X
+ sky130_fd_sc_hs__dlrtp_1_31/Q sky130_fd_sc_hs__einvp_2_43/a_263_323# sky130_fd_sc_hs__einvp_2_43/a_36_74#
+ sky130_fd_sc_hs__einvp_2_43/a_27_368# sky130_fd_sc_hs__einvp_2
Xsky130_fd_sc_hs__clkbuf_4_9 DVSS: DVDD: DVDD: DVSS: pi1_con[0] sky130_fd_sc_hs__clkbuf_8_5/A
+ sky130_fd_sc_hs__clkbuf_4_9/a_83_270# sky130_fd_sc_hs__clkbuf_4
Xsky130_fd_sc_hs__einvp_2_53 DVSS: DVDD: DVDD: DVSS: dout_p sky130_fd_sc_hs__inv_4_9/Y
+ sky130_fd_sc_hs__dlrtp_1_45/Q sky130_fd_sc_hs__einvp_2_53/a_263_323# sky130_fd_sc_hs__einvp_2_53/a_36_74#
+ sky130_fd_sc_hs__einvp_2_53/a_27_368# sky130_fd_sc_hs__einvp_2
Xsky130_fd_sc_hs__einvp_2_64 DVSS: DVDD: DVDD: DVSS: dout_p sky130_fd_sc_hs__einvp_2_65/A
+ sky130_fd_sc_hs__dlrtp_1_53/Q sky130_fd_sc_hs__einvp_2_65/a_263_323# sky130_fd_sc_hs__einvp_2_65/a_36_74#
+ sky130_fd_sc_hs__einvp_2_65/a_27_368# sky130_fd_sc_hs__einvp_2
Xsky130_fd_sc_hs__einvp_2_75 DVSS: DVDD: DVDD: DVSS: dout_p sky130_fd_sc_hs__einvp_2_99/A
+ sky130_fd_sc_hs__einvp_2_75/TE sky130_fd_sc_hs__einvp_2_75/a_263_323# sky130_fd_sc_hs__einvp_2_75/a_36_74#
+ sky130_fd_sc_hs__einvp_2_75/a_27_368# sky130_fd_sc_hs__einvp_2
Xsky130_fd_sc_hs__einvp_2_86 DVSS: DVDD: DVDD: DVSS: dout_p sky130_fd_sc_hs__einvp_2_97/A
+ sky130_fd_sc_hs__dlrtp_1_63/Q sky130_fd_sc_hs__einvp_2_87/a_263_323# sky130_fd_sc_hs__einvp_2_87/a_36_74#
+ sky130_fd_sc_hs__einvp_2_87/a_27_368# sky130_fd_sc_hs__einvp_2
Xsky130_fd_sc_hs__einvp_2_97 DVSS: DVDD: DVDD: DVSS: dout_p sky130_fd_sc_hs__einvp_2_97/A
+ sky130_fd_sc_hs__dlrtp_1_79/Q sky130_fd_sc_hs__einvp_2_97/a_263_323# sky130_fd_sc_hs__einvp_2_97/a_36_74#
+ sky130_fd_sc_hs__einvp_2_97/a_27_368# sky130_fd_sc_hs__einvp_2
Xsky130_fd_sc_hs__or2b_2_1 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__or2b_2_1/X sky130_fd_sc_hs__nor2_4_1/Y
+ sky130_fd_sc_hs__or2b_2_1/A sky130_fd_sc_hs__or2b_2_1/a_470_368# sky130_fd_sc_hs__or2b_2_1/a_27_368#
+ sky130_fd_sc_hs__or2b_2_1/a_187_48# sky130_fd_sc_hs__or2b_2
Xsky130_fd_sc_hs__clkinv_4_9 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__nor2_4_1/B sky130_fd_sc_hs__o21ai_4_1/A1
+ sky130_fd_sc_hs__clkinv_4
Xsky130_fd_sc_hs__conb_1_30 DVSS: DVDD: DVDD: DVSS: prbs_generator_syn_5/eqn[23] prbs_generator_syn_5/eqn[20]
+ sky130_fd_sc_hs__conb_1_31/a_165_290# sky130_fd_sc_hs__conb_1_31/a_21_290# sky130_fd_sc_hs__conb_1
Xsky130_fd_sc_hs__conb_1_41 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__conb_1_41/LO
+ sky130_fd_sc_hs__conb_1_41/HI sky130_fd_sc_hs__conb_1_41/a_165_290# sky130_fd_sc_hs__conb_1_41/a_21_290#
+ sky130_fd_sc_hs__conb_1
Xsky130_fd_sc_hs__conb_1_52 DVSS: DVDD: DVDD: DVSS: prbs_generator_syn_7/eqn[21] prbs_generator_syn_7/eqn[20]
+ sky130_fd_sc_hs__conb_1_53/a_165_290# sky130_fd_sc_hs__conb_1_53/a_21_290# sky130_fd_sc_hs__conb_1
Xsky130_fd_sc_hs__conb_1_63 DVSS: DVDD: DVDD: DVSS: prbs_generator_syn_7/eqn[0] sky130_fd_sc_hs__conb_1_63/HI
+ sky130_fd_sc_hs__conb_1_63/a_165_290# sky130_fd_sc_hs__conb_1_63/a_21_290# sky130_fd_sc_hs__conb_1
Xsky130_fd_sc_hs__conb_1_74 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__conb_1_75/LO
+ sky130_fd_sc_hs__conb_1_75/HI sky130_fd_sc_hs__conb_1_75/a_165_290# sky130_fd_sc_hs__conb_1_75/a_21_290#
+ sky130_fd_sc_hs__conb_1
Xsky130_fd_sc_hs__conb_1_85 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__conb_1_85/LO
+ sky130_fd_sc_hs__conb_1_85/HI sky130_fd_sc_hs__conb_1_85/a_165_290# sky130_fd_sc_hs__conb_1_85/a_21_290#
+ sky130_fd_sc_hs__conb_1
Xsky130_fd_sc_hs__conb_1_96 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__conb_1_97/LO
+ sky130_fd_sc_hs__conb_1_97/HI sky130_fd_sc_hs__conb_1_97/a_165_290# sky130_fd_sc_hs__conb_1_97/a_21_290#
+ sky130_fd_sc_hs__conb_1
Xsky130_fd_sc_hs__inv_4_70 DVSS: DVDD: DVDD: DVSS: osc_core_1/pi5_r[0] osc_core_1/pi5_l[0]
+ sky130_fd_sc_hs__inv_4
Xsky130_fd_sc_hs__inv_4_81 DVSS: DVDD: DVDD: DVSS: hr_16t4_mux_top_3/din[8] hr_16t4_mux_top_1/din[8]
+ sky130_fd_sc_hs__inv_4
Xsky130_fd_sc_hs__dlrtp_1_108 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__buf_2_115/A
+ sky130_fd_sc_hs__dlrtp_1_9/GATE sky130_fd_sc_hs__conb_1_133/HI sky130_fd_sc_hs__inv_4_23/A
+ sky130_fd_sc_hs__dlrtp_1_109/a_216_424# sky130_fd_sc_hs__dlrtp_1_109/a_759_508#
+ sky130_fd_sc_hs__dlrtp_1_109/a_565_74# sky130_fd_sc_hs__dlrtp_1_109/a_27_424# sky130_fd_sc_hs__dlrtp_1_109/a_1045_74#
+ sky130_fd_sc_hs__dlrtp_1_109/a_643_74# sky130_fd_sc_hs__dlrtp_1_109/a_817_48# sky130_fd_sc_hs__dlrtp_1_109/a_568_392#
+ sky130_fd_sc_hs__dlrtp_1_109/a_363_74# sky130_fd_sc_hs__dlrtp_1_109/a_769_74# sky130_fd_sc_hs__dlrtp_1
Xsky130_fd_sc_hs__dlrtp_1_119 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__dlrtp_1_119/Q
+ sky130_fd_sc_hs__dlrtp_1_9/GATE sky130_fd_sc_hs__conb_1_131/HI sky130_fd_sc_hs__buf_2_117/X
+ sky130_fd_sc_hs__dlrtp_1_119/a_216_424# sky130_fd_sc_hs__dlrtp_1_119/a_759_508#
+ sky130_fd_sc_hs__dlrtp_1_119/a_565_74# sky130_fd_sc_hs__dlrtp_1_119/a_27_424# sky130_fd_sc_hs__dlrtp_1_119/a_1045_74#
+ sky130_fd_sc_hs__dlrtp_1_119/a_643_74# sky130_fd_sc_hs__dlrtp_1_119/a_817_48# sky130_fd_sc_hs__dlrtp_1_119/a_568_392#
+ sky130_fd_sc_hs__dlrtp_1_119/a_363_74# sky130_fd_sc_hs__dlrtp_1_119/a_769_74# sky130_fd_sc_hs__dlrtp_1
Xsky130_fd_sc_hs__dlrtp_1_10 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__dlrtp_1_8/Q
+ sky130_fd_sc_hs__dlrtp_1_9/GATE sky130_fd_sc_hs__conb_1_117/HI sky130_fd_sc_hs__dlrtp_1_8/D
+ sky130_fd_sc_hs__dlrtp_1_8/a_216_424# sky130_fd_sc_hs__dlrtp_1_8/a_759_508# sky130_fd_sc_hs__dlrtp_1_8/a_565_74#
+ sky130_fd_sc_hs__dlrtp_1_8/a_27_424# sky130_fd_sc_hs__dlrtp_1_8/a_1045_74# sky130_fd_sc_hs__dlrtp_1_8/a_643_74#
+ sky130_fd_sc_hs__dlrtp_1_8/a_817_48# sky130_fd_sc_hs__dlrtp_1_8/a_568_392# sky130_fd_sc_hs__dlrtp_1_8/a_363_74#
+ sky130_fd_sc_hs__dlrtp_1_8/a_769_74# sky130_fd_sc_hs__dlrtp_1
Xsky130_fd_sc_hs__dlrtp_1_21 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__dlrtp_1_21/Q
+ sky130_fd_sc_hs__clkbuf_2_3/X sky130_fd_sc_hs__conb_1_119/HI sky130_fd_sc_hs__dlrtp_1_21/D
+ sky130_fd_sc_hs__dlrtp_1_21/a_216_424# sky130_fd_sc_hs__dlrtp_1_21/a_759_508# sky130_fd_sc_hs__dlrtp_1_21/a_565_74#
+ sky130_fd_sc_hs__dlrtp_1_21/a_27_424# sky130_fd_sc_hs__dlrtp_1_21/a_1045_74# sky130_fd_sc_hs__dlrtp_1_21/a_643_74#
+ sky130_fd_sc_hs__dlrtp_1_21/a_817_48# sky130_fd_sc_hs__dlrtp_1_21/a_568_392# sky130_fd_sc_hs__dlrtp_1_21/a_363_74#
+ sky130_fd_sc_hs__dlrtp_1_21/a_769_74# sky130_fd_sc_hs__dlrtp_1
Xsky130_fd_sc_hs__dlrtp_1_32 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__dlrtp_1_33/Q
+ sky130_fd_sc_hs__clkbuf_2_3/A sky130_fd_sc_hs__conb_1_123/HI sky130_fd_sc_hs__buf_2_15/X
+ sky130_fd_sc_hs__dlrtp_1_33/a_216_424# sky130_fd_sc_hs__dlrtp_1_33/a_759_508# sky130_fd_sc_hs__dlrtp_1_33/a_565_74#
+ sky130_fd_sc_hs__dlrtp_1_33/a_27_424# sky130_fd_sc_hs__dlrtp_1_33/a_1045_74# sky130_fd_sc_hs__dlrtp_1_33/a_643_74#
+ sky130_fd_sc_hs__dlrtp_1_33/a_817_48# sky130_fd_sc_hs__dlrtp_1_33/a_568_392# sky130_fd_sc_hs__dlrtp_1_33/a_363_74#
+ sky130_fd_sc_hs__dlrtp_1_33/a_769_74# sky130_fd_sc_hs__dlrtp_1
Xsky130_fd_sc_hs__dlrtp_1_43 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__dlrtp_1_43/Q
+ sky130_fd_sc_hs__clkbuf_16_53/A sky130_fd_sc_hs__conb_1_135/HI sky130_fd_sc_hs__buf_2_23/X
+ sky130_fd_sc_hs__dlrtp_1_43/a_216_424# sky130_fd_sc_hs__dlrtp_1_43/a_759_508# sky130_fd_sc_hs__dlrtp_1_43/a_565_74#
+ sky130_fd_sc_hs__dlrtp_1_43/a_27_424# sky130_fd_sc_hs__dlrtp_1_43/a_1045_74# sky130_fd_sc_hs__dlrtp_1_43/a_643_74#
+ sky130_fd_sc_hs__dlrtp_1_43/a_817_48# sky130_fd_sc_hs__dlrtp_1_43/a_568_392# sky130_fd_sc_hs__dlrtp_1_43/a_363_74#
+ sky130_fd_sc_hs__dlrtp_1_43/a_769_74# sky130_fd_sc_hs__dlrtp_1
Xsky130_fd_sc_hs__dlrtp_1_54 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__dlrtp_1_55/Q
+ sky130_fd_sc_hs__clkbuf_16_53/A sky130_fd_sc_hs__conb_1_135/HI sky130_fd_sc_hs__dlrtp_1_55/D
+ sky130_fd_sc_hs__dlrtp_1_55/a_216_424# sky130_fd_sc_hs__dlrtp_1_55/a_759_508# sky130_fd_sc_hs__dlrtp_1_55/a_565_74#
+ sky130_fd_sc_hs__dlrtp_1_55/a_27_424# sky130_fd_sc_hs__dlrtp_1_55/a_1045_74# sky130_fd_sc_hs__dlrtp_1_55/a_643_74#
+ sky130_fd_sc_hs__dlrtp_1_55/a_817_48# sky130_fd_sc_hs__dlrtp_1_55/a_568_392# sky130_fd_sc_hs__dlrtp_1_55/a_363_74#
+ sky130_fd_sc_hs__dlrtp_1_55/a_769_74# sky130_fd_sc_hs__dlrtp_1
Xsky130_fd_sc_hs__dlrtp_1_65 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__dlrtp_1_65/Q
+ sky130_fd_sc_hs__clkbuf_16_53/A sky130_fd_sc_hs__conb_1_129/HI sky130_fd_sc_hs__dlrtp_1_65/D
+ sky130_fd_sc_hs__dlrtp_1_65/a_216_424# sky130_fd_sc_hs__dlrtp_1_65/a_759_508# sky130_fd_sc_hs__dlrtp_1_65/a_565_74#
+ sky130_fd_sc_hs__dlrtp_1_65/a_27_424# sky130_fd_sc_hs__dlrtp_1_65/a_1045_74# sky130_fd_sc_hs__dlrtp_1_65/a_643_74#
+ sky130_fd_sc_hs__dlrtp_1_65/a_817_48# sky130_fd_sc_hs__dlrtp_1_65/a_568_392# sky130_fd_sc_hs__dlrtp_1_65/a_363_74#
+ sky130_fd_sc_hs__dlrtp_1_65/a_769_74# sky130_fd_sc_hs__dlrtp_1
Xsky130_fd_sc_hs__dlrtp_1_76 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__dlrtp_1_77/Q
+ sky130_fd_sc_hs__clkbuf_16_53/A sky130_fd_sc_hs__conb_1_129/HI sky130_fd_sc_hs__inv_4_15/A
+ sky130_fd_sc_hs__dlrtp_1_77/a_216_424# sky130_fd_sc_hs__dlrtp_1_77/a_759_508# sky130_fd_sc_hs__dlrtp_1_77/a_565_74#
+ sky130_fd_sc_hs__dlrtp_1_77/a_27_424# sky130_fd_sc_hs__dlrtp_1_77/a_1045_74# sky130_fd_sc_hs__dlrtp_1_77/a_643_74#
+ sky130_fd_sc_hs__dlrtp_1_77/a_817_48# sky130_fd_sc_hs__dlrtp_1_77/a_568_392# sky130_fd_sc_hs__dlrtp_1_77/a_363_74#
+ sky130_fd_sc_hs__dlrtp_1_77/a_769_74# sky130_fd_sc_hs__dlrtp_1
Xsky130_fd_sc_hs__dlrtp_1_87 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__buf_2_159/A
+ sky130_fd_sc_hs__clkbuf_16_53/X sky130_fd_sc_hs__conb_1_137/HI sky130_fd_sc_hs__dlrtp_1_87/D
+ sky130_fd_sc_hs__dlrtp_1_87/a_216_424# sky130_fd_sc_hs__dlrtp_1_87/a_759_508# sky130_fd_sc_hs__dlrtp_1_87/a_565_74#
+ sky130_fd_sc_hs__dlrtp_1_87/a_27_424# sky130_fd_sc_hs__dlrtp_1_87/a_1045_74# sky130_fd_sc_hs__dlrtp_1_87/a_643_74#
+ sky130_fd_sc_hs__dlrtp_1_87/a_817_48# sky130_fd_sc_hs__dlrtp_1_87/a_568_392# sky130_fd_sc_hs__dlrtp_1_87/a_363_74#
+ sky130_fd_sc_hs__dlrtp_1_87/a_769_74# sky130_fd_sc_hs__dlrtp_1
Xsky130_fd_sc_hs__dlrtp_1_98 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__dlrtp_1_98/Q
+ sky130_fd_sc_hs__dlrtp_1_9/GATE sky130_fd_sc_hs__conb_1_95/HI sky130_fd_sc_hs__dlrtp_1_98/D
+ sky130_fd_sc_hs__dlrtp_1_98/a_216_424# sky130_fd_sc_hs__dlrtp_1_98/a_759_508# sky130_fd_sc_hs__dlrtp_1_98/a_565_74#
+ sky130_fd_sc_hs__dlrtp_1_98/a_27_424# sky130_fd_sc_hs__dlrtp_1_98/a_1045_74# sky130_fd_sc_hs__dlrtp_1_98/a_643_74#
+ sky130_fd_sc_hs__dlrtp_1_98/a_817_48# sky130_fd_sc_hs__dlrtp_1_98/a_568_392# sky130_fd_sc_hs__dlrtp_1_98/a_363_74#
+ sky130_fd_sc_hs__dlrtp_1_98/a_769_74# sky130_fd_sc_hs__dlrtp_1
Xsky130_fd_sc_hs__einvp_2_3 DVSS: DVDD: DVDD: DVSS: dout_n sky130_fd_sc_hs__einvp_2_9/A
+ sky130_fd_sc_hs__einvp_2_3/TE sky130_fd_sc_hs__einvp_2_3/a_263_323# sky130_fd_sc_hs__einvp_2_3/a_36_74#
+ sky130_fd_sc_hs__einvp_2_3/a_27_368# sky130_fd_sc_hs__einvp_2
Xsky130_fd_sc_hs__clkbuf_2_6 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__clkbuf_2_7/X
+ sky130_fd_sc_hs__o21ai_2_5/Y sky130_fd_sc_hs__clkbuf_2_7/a_43_192# sky130_fd_sc_hs__clkbuf_2
Xsky130_fd_sc_hs__clkbuf_2_17 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__dlrtp_1_69/D
+ sky130_fd_sc_hs__buf_2_69/X sky130_fd_sc_hs__clkbuf_2_17/a_43_192# sky130_fd_sc_hs__clkbuf_2
Xsky130_fd_sc_hs__clkbuf_2_28 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__dlrtp_1_79/D
+ sky130_fd_sc_hs__o21ai_2_23/Y sky130_fd_sc_hs__clkbuf_2_28/a_43_192# sky130_fd_sc_hs__clkbuf_2
Xsky130_fd_sc_hs__clkbuf_2_39 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__dlrtp_1_99/D
+ sky130_fd_sc_hs__buf_2_129/X sky130_fd_sc_hs__clkbuf_2_39/a_43_192# sky130_fd_sc_hs__clkbuf_2
Xsky130_fd_sc_hs__buf_2_8 DVSS: DVDD: DVDD: DVSS: manual_control_osc[11] sky130_fd_sc_hs__buf_2_9/X
+ sky130_fd_sc_hs__buf_2_9/a_21_260# sky130_fd_sc_hs__buf_2
Xsky130_fd_sc_hs__buf_2_13 DVSS: DVDD: DVDD: DVSS: manual_control_osc[1] sky130_fd_sc_hs__buf_2_13/X
+ sky130_fd_sc_hs__buf_2_13/a_21_260# sky130_fd_sc_hs__buf_2
Xsky130_fd_sc_hs__buf_2_24 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__buf_2_25/A sky130_fd_sc_hs__buf_2_25/X
+ sky130_fd_sc_hs__buf_2_25/a_21_260# sky130_fd_sc_hs__buf_2
Xsky130_fd_sc_hs__buf_2_35 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__buf_2_35/A sky130_fd_sc_hs__buf_2_35/X
+ sky130_fd_sc_hs__buf_2_35/a_21_260# sky130_fd_sc_hs__buf_2
Xsky130_fd_sc_hs__buf_2_46 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__buf_2_47/A sky130_fd_sc_hs__buf_2_47/X
+ sky130_fd_sc_hs__buf_2_47/a_21_260# sky130_fd_sc_hs__buf_2
Xsky130_fd_sc_hs__buf_2_57 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__buf_2_57/A sky130_fd_sc_hs__buf_2_57/X
+ sky130_fd_sc_hs__buf_2_57/a_21_260# sky130_fd_sc_hs__buf_2
Xsky130_fd_sc_hs__buf_2_68 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__buf_2_69/A sky130_fd_sc_hs__buf_2_69/X
+ sky130_fd_sc_hs__buf_2_69/a_21_260# sky130_fd_sc_hs__buf_2
Xsky130_fd_sc_hs__buf_2_79 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__buf_2_79/A sky130_fd_sc_hs__buf_2_79/X
+ sky130_fd_sc_hs__buf_2_79/a_21_260# sky130_fd_sc_hs__buf_2
Xsky130_fd_sc_hs__o21bai_2_15 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__nand2_2_7/A
+ sky130_fd_sc_hs__o21bai_2_3/A2 sky130_fd_sc_hs__dlrtp_1_87/D sky130_fd_sc_hs__buf_2_67/A
+ sky130_fd_sc_hs__o21bai_2_15/a_27_74# sky130_fd_sc_hs__o21bai_2_15/a_225_74# sky130_fd_sc_hs__o21bai_2_15/a_507_368#
+ sky130_fd_sc_hs__o21bai_2
Xsky130_fd_sc_hs__o21bai_2_26 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__or2b_2_3/A
+ sky130_fd_sc_hs__clkbuf_4_81/X sky130_fd_sc_hs__dlrtp_1_99/D sky130_fd_sc_hs__buf_2_105/A
+ sky130_fd_sc_hs__o21bai_2_27/a_27_74# sky130_fd_sc_hs__o21bai_2_27/a_225_74# sky130_fd_sc_hs__o21bai_2_27/a_507_368#
+ sky130_fd_sc_hs__o21bai_2
Xsky130_fd_sc_hs__o21bai_2_37 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__o21ai_4_1/A1
+ sky130_fd_sc_hs__clkinv_4_3/Y sky130_fd_sc_hs__dlrtp_1_21/D sky130_fd_sc_hs__o21bai_2_37/Y
+ sky130_fd_sc_hs__o21bai_2_37/a_27_74# sky130_fd_sc_hs__o21bai_2_37/a_225_74# sky130_fd_sc_hs__o21bai_2_37/a_507_368#
+ sky130_fd_sc_hs__o21bai_2
Xsky130_fd_sc_hs__o21bai_2_48 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__nand2_8_1/Y
+ sky130_fd_sc_hs__nand2_2_21/B sky130_fd_sc_hs__dlrtp_1_121/D sky130_fd_sc_hs__o21bai_2_49/Y
+ sky130_fd_sc_hs__o21bai_2_49/a_27_74# sky130_fd_sc_hs__o21bai_2_49/a_225_74# sky130_fd_sc_hs__o21bai_2_49/a_507_368#
+ sky130_fd_sc_hs__o21bai_2
Xsky130_fd_sc_hs__o21bai_2_59 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__nand2_2_9/B
+ sky130_fd_sc_hs__o21bai_2_3/A2 sky130_fd_sc_hs__clkbuf_2_7/X sky130_fd_sc_hs__buf_2_37/A
+ sky130_fd_sc_hs__o21bai_2_59/a_27_74# sky130_fd_sc_hs__o21bai_2_59/a_225_74# sky130_fd_sc_hs__o21bai_2_59/a_507_368#
+ sky130_fd_sc_hs__o21bai_2
Xsky130_fd_sc_hs__o21bai_4_4 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__buf_2_143/A
+ sky130_fd_sc_hs__nand2_2_5/B sky130_fd_sc_hs__o21bai_4_7/A1 sky130_fd_sc_hs__buf_2_153/X
+ sky130_fd_sc_hs__o21bai_4_5/a_28_368# sky130_fd_sc_hs__o21bai_4_5/a_27_74# sky130_fd_sc_hs__o21bai_4_5/a_828_48#
+ sky130_fd_sc_hs__o21bai_4
Xsky130_fd_sc_hs__conb_1_202 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__conb_1_203/LO
+ sky130_fd_sc_hs__conb_1_203/HI sky130_fd_sc_hs__conb_1_203/a_165_290# sky130_fd_sc_hs__conb_1_203/a_21_290#
+ sky130_fd_sc_hs__conb_1
Xsky130_fd_sc_hs__conb_1_213 DVSS: DVDD: DVDD: DVSS: prbs_generator_syn_21/eqn[31]
+ prbs_generator_syn_21/cke sky130_fd_sc_hs__conb_1_213/a_165_290# sky130_fd_sc_hs__conb_1_213/a_21_290#
+ sky130_fd_sc_hs__conb_1
Xsky130_fd_sc_hs__conb_1_224 DVSS: DVDD: DVDD: DVSS: prbs_generator_syn_25/eqn[8]
+ prbs_generator_syn_25/eqn[1] sky130_fd_sc_hs__conb_1_225/a_165_290# sky130_fd_sc_hs__conb_1_225/a_21_290#
+ sky130_fd_sc_hs__conb_1
Xsky130_fd_sc_hs__conb_1_235 DVSS: DVDD: DVDD: DVSS: prbs_generator_syn_27/eqn[8]
+ prbs_generator_syn_27/eqn[1] sky130_fd_sc_hs__conb_1_235/a_165_290# sky130_fd_sc_hs__conb_1_235/a_21_290#
+ sky130_fd_sc_hs__conb_1
Xsky130_fd_sc_hs__conb_1_246 DVSS: DVDD: DVDD: DVSS: prbs_generator_syn_31/eqn[28]
+ sky130_fd_sc_hs__conb_1_247/HI sky130_fd_sc_hs__conb_1_247/a_165_290# sky130_fd_sc_hs__conb_1_247/a_21_290#
+ sky130_fd_sc_hs__conb_1
Xsky130_fd_sc_hs__conb_1_257 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__conb_1_257/LO
+ sky130_fd_sc_hs__conb_1_257/HI sky130_fd_sc_hs__conb_1_257/a_165_290# sky130_fd_sc_hs__conb_1_257/a_21_290#
+ sky130_fd_sc_hs__conb_1
Xsky130_fd_sc_hs__conb_1_268 DVSS: DVDD: DVDD: DVSS: prbs_generator_syn_31/eqn[2]
+ prbs_generator_syn_31/eqn[1] sky130_fd_sc_hs__conb_1_269/a_165_290# sky130_fd_sc_hs__conb_1_269/a_21_290#
+ sky130_fd_sc_hs__conb_1
Xsky130_fd_sc_hs__clkbuf_8_16 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__clkbuf_8_17/X
+ sky130_fd_sc_hs__buf_2_9/X sky130_fd_sc_hs__clkbuf_8_17/a_125_368# sky130_fd_sc_hs__clkbuf_8
Xsky130_fd_sc_hs__clkbuf_8_27 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__clkbuf_8_27/X
+ sky130_fd_sc_hs__clkbuf_8_27/A sky130_fd_sc_hs__clkbuf_8_27/a_125_368# sky130_fd_sc_hs__clkbuf_8
Xsky130_fd_sc_hs__clkbuf_8_38 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__nand2_2_21/B
+ sky130_fd_sc_hs__or2b_2_3/X sky130_fd_sc_hs__clkbuf_8_39/a_125_368# sky130_fd_sc_hs__clkbuf_8
Xsky130_fd_sc_hs__clkbuf_8_49 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__nand2_2_5/B
+ sky130_fd_sc_hs__or2b_4_3/X sky130_fd_sc_hs__clkbuf_8_49/a_125_368# sky130_fd_sc_hs__clkbuf_8
Xsky130_fd_sc_hs__o21bai_2_1 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__o21bai_2_3/A2
+ sky130_fd_sc_hs__nand2_2_3/B sky130_fd_sc_hs__dlrtp_1_53/D sky130_fd_sc_hs__buf_2_25/A
+ sky130_fd_sc_hs__o21bai_2_1/a_27_74# sky130_fd_sc_hs__o21bai_2_1/a_225_74# sky130_fd_sc_hs__o21bai_2_1/a_507_368#
+ sky130_fd_sc_hs__o21bai_2
Xsky130_fd_sc_hs__nand2_2_9 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__inv_4_15/A sky130_fd_sc_hs__nand2_2_9/B
+ sky130_fd_sc_hs__buf_2_65/X sky130_fd_sc_hs__nand2_2_9/a_27_74# sky130_fd_sc_hs__nand2_2
Xsky130_fd_sc_hs__o21ai_2_50 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__inv_4_25/Y sky130_fd_sc_hs__or2b_4_1/A
+ sky130_fd_sc_hs__o21ai_2_51/A1 sky130_fd_sc_hs__o21ai_2_51/Y sky130_fd_sc_hs__o21ai_2_51/a_116_368#
+ sky130_fd_sc_hs__o21ai_2_51/a_27_74# sky130_fd_sc_hs__o21ai_2
Xsky130_fd_sc_hs__or2b_4_5 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__or2b_4_5/A sky130_fd_sc_hs__or4_2_1/A
+ sky130_fd_sc_hs__or2b_4_5/X sky130_fd_sc_hs__or2b_4_5/a_676_48# sky130_fd_sc_hs__or2b_4_5/a_489_392#
+ sky130_fd_sc_hs__or2b_4_5/a_81_296# sky130_fd_sc_hs__or2b_4
Xprbs_generator_syn_11 prbs_generator_syn_9/clk prbs_generator_syn_9/rst prbs_generator_syn_11/cke
+ sky130_fd_sc_hs__conb_1_91/LO sky130_fd_sc_hs__conb_1_91/LO sky130_fd_sc_hs__conb_1_91/LO
+ sky130_fd_sc_hs__conb_1_91/LO sky130_fd_sc_hs__conb_1_91/HI sky130_fd_sc_hs__conb_1_91/HI
+ sky130_fd_sc_hs__conb_1_91/HI sky130_fd_sc_hs__conb_1_91/HI sky130_fd_sc_hs__conb_1_91/HI
+ sky130_fd_sc_hs__conb_1_91/HI sky130_fd_sc_hs__conb_1_91/HI prbs_generator_syn_11/cke
+ prbs_generator_syn_11/cke prbs_generator_syn_11/cke sky130_fd_sc_hs__conb_1_81/LO
+ prbs_generator_syn_11/cke sky130_fd_sc_hs__conb_1_81/LO prbs_generator_syn_11/cke
+ prbs_generator_syn_11/eqn[2] prbs_generator_syn_11/eqn[2] prbs_generator_syn_11/eqn[2]
+ prbs_generator_syn_11/eqn[2] prbs_generator_syn_11/eqn[2] prbs_generator_syn_11/eqn[2]
+ sky130_fd_sc_hs__conb_1_89/LO sky130_fd_sc_hs__conb_1_89/HI sky130_fd_sc_hs__conb_1_89/HI
+ sky130_fd_sc_hs__conb_1_89/LO sky130_fd_sc_hs__conb_1_89/LO sky130_fd_sc_hs__conb_1_89/HI
+ sky130_fd_sc_hs__conb_1_89/HI sky130_fd_sc_hs__conb_1_89/LO sky130_fd_sc_hs__conb_1_81/LO
+ sky130_fd_sc_hs__conb_1_79/LO sky130_fd_sc_hs__conb_1_79/LO sky130_fd_sc_hs__conb_1_77/LO
+ sky130_fd_sc_hs__conb_1_77/LO sky130_fd_sc_hs__conb_1_77/LO sky130_fd_sc_hs__conb_1_77/LO
+ sky130_fd_sc_hs__conb_1_77/LO sky130_fd_sc_hs__conb_1_65/LO sky130_fd_sc_hs__conb_1_65/LO
+ sky130_fd_sc_hs__conb_1_65/LO sky130_fd_sc_hs__conb_1_65/HI sky130_fd_sc_hs__conb_1_65/LO
+ sky130_fd_sc_hs__conb_1_65/LO sky130_fd_sc_hs__conb_1_65/LO sky130_fd_sc_hs__conb_1_65/LO
+ prbs_generator_syn_7/eqn[0] prbs_generator_syn_7/eqn[0] prbs_generator_syn_7/eqn[0]
+ prbs_generator_syn_7/eqn[0] prbs_generator_syn_7/eqn[0] prbs_generator_syn_7/eqn[0]
+ prbs_generator_syn_11/eqn[9] prbs_generator_syn_11/eqn[9] prbs_generator_syn_11/eqn[9]
+ prbs_generator_syn_11/eqn[9] prbs_generator_syn_11/eqn[9] prbs_generator_syn_11/eqn[9]
+ prbs_generator_syn_11/eqn[9] prbs_generator_syn_11/eqn[2] prbs_generator_syn_11/eqn[1]
+ prbs_generator_syn_11/eqn[2] prbs_generator_syn_9/inj_err sky130_fd_sc_hs__conb_1_81/LO
+ sky130_fd_sc_hs__conb_1_81/LO prbs_generator_syn_11/out DVSS: DVDD: prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_1/a_293_74#
+ prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_15/X prbs_generator_syn_11/sky130_fd_sc_hs__nand2_1_35/B
+ prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_51/Y prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_9/A
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_9/CLK prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_47/a_27_74#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_37/a_1226_296# prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_3/B
+ prbs_generator_syn_11/sky130_fd_sc_hs__nor2b_1_7/a_27_112# prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_29/B
+ prbs_generator_syn_11/sky130_fd_sc_hs__sdlclkp_2_1/a_580_74# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_1/a_1141_508#
+ prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_5/Y prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_41/a_230_79#
+ prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_61/a_138_385# prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_43/a_132_392#
+ prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_3/a_222_392# prbs_generator_syn_11/sky130_fd_sc_hs__nor2b_1_9/a_27_112#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_61/a_27_74# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_35/a_206_368#
+ prbs_generator_syn_11/sky130_fd_sc_hs__nand2_2_3/Y prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_25/B
+ prbs_generator_syn_11/sky130_fd_sc_hs__nand2_1_11/a_117_74# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_67/a_651_503#
+ prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_45/X prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_39/a_696_458#
+ prbs_generator_syn_11/sky130_fd_sc_hs__sdlclkp_2_1/a_1198_74# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_45/a_1034_424#
+ prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_17/a_222_392# prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_55/a_222_392#
+ prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_53/Y prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_35/A
+ prbs_generator_syn_11/m3_13600_1651# prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_59/a_52_123#
+ prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_5/a_293_74# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_35/a_1226_296#
+ prbs_generator_syn_11/sky130_fd_sc_hs__nand2_1_51/B prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_5/a_651_503#
+ prbs_generator_syn_11/sky130_fd_sc_hs__nand2_1_21/B prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_8/a_27_74#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_15/a_27_74# prbs_generator_syn_11/sky130_fd_sc_hs__and2b_2_1/X
+ prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_13/X prbs_generator_syn_11/sky130_fd_sc_hs__nand2_2_3/a_27_74#
+ prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_50/a_138_385# prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_33/a_132_392#
+ prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_1/a_376_368# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_25/a_206_368#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_35/a_437_503# prbs_generator_syn_11/sky130_fd_sc_hs__sdlclkp_2_1/a_708_451#
+ prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_45/a_230_79# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_29/a_696_458#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_32/a_27_74# prbs_generator_syn_11/sky130_fd_sc_hs__nor2b_1_4/Y
+ prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_59/a_293_74# prbs_generator_syn_11/sky130_fd_sc_hs__nand2_1_47/a_117_74#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_73/a_735_102# prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_21/a_112_119#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_23/a_1141_508# prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_25/a_293_74#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_7/Q prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_3/a_112_119#
+ prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_35/B prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_51/X
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_53/a_1178_124# prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_23/a_132_392#
+ prbs_generator_syn_11/sky130_fd_sc_hs__nand2_1_3/B prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_15/a_206_368#
+ prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_63/a_132_392# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_55/a_27_74#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_25/a_437_503# prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_41/a_52_123#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_47/a_651_503# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_73/a_1141_508#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_19/a_696_458# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_57/a_696_458#
+ prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_7/X prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_43/a_1034_424#
+ prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_55/A prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_11/a_112_119#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_21/a_1141_508# prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_35/a_222_392#
+ prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_49/a_230_79# prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_67/Y
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_71/a_27_74# prbs_generator_syn_11/sky130_fd_sc_hs__nand2_1_33/B
+ prbs_generator_syn_11/sky130_fd_sc_hs__conb_1_1/LO prbs_generator_syn_11/sky130_fd_sc_hs__nand2_1_19/a_117_74#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_51/a_1178_124# prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_33/X
+ prbs_generator_syn_11/sky130_fd_sc_hs__nand2_1_29/B prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_41/Y
+ prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_53/a_132_392# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_45/a_206_368#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_15/a_437_503# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_37/a_651_503#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_39/a_544_485# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_53/a_735_102#
+ prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_45/a_52_123# prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_1/B
+ prbs_generator_syn_11/sky130_fd_sc_hs__nand2_2_3/B prbs_generator_syn_11/sky130_fd_sc_hs__clkbuf_16_1/A
+ prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_21/X prbs_generator_syn_11/sky130_fd_sc_hs__nand2_1_25/B
+ prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_39/a_376_368# prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_63/X
+ prbs_generator_syn_11/m3_13600_3481# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_69/a_1178_124#
+ prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_21/a_138_385# prbs_generator_syn_11/sky130_fd_sc_hs__nor2b_1_8/Y
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_19/a_1178_124# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_49/a_27_74#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_45/a_437_503# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_27/a_651_503#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_71/a_1141_508# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_65/a_651_503#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_29/a_544_485# prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_3/a_138_385#
+ prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_55/X prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_43/a_735_102#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_41/a_1034_424# prbs_generator_syn_11/sky130_fd_sc_hs__nand2_1_9/B
+ prbs_generator_syn_11/sky130_fd_sc_hs__nor2b_1_9/Y prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_59/a_1034_424#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_39/a_1141_508# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_33/a_1226_296#
+ prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_49/a_52_123# prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_47/Y
+ prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_43/Y prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_4/a_651_503#
+ prbs_generator_syn_11/sky130_fd_sc_hs__nand2_1_49/B prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_19/A
+ prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_11/a_138_385# prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_5/X
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_63/a_206_368# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_17/a_651_503#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_19/a_544_485# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_55/a_651_503#
+ prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_9/Y prbs_generator_syn_11/sky130_fd_sc_hs__nand2_1_17/B
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_57/a_544_485# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_67/a_696_458#
+ prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_35/X prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_19/a_27_74#
+ prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_45/a_222_392# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_32/a_1226_296#
+ prbs_generator_syn_11/sky130_fd_sc_hs__nand2_1_43/B prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_25/A
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_1/a_206_368# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_49/a_1226_296#
+ prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_1/a_112_119# prbs_generator_syn_11/sky130_fd_sc_hs__or2_1_1/X
+ prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_59/a_376_368# prbs_generator_syn_11/sky130_fd_sc_hs__nand2_1_19/B
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_5/a_696_458# prbs_generator_syn_11/sky130_fd_sc_hs__nor2b_1_1/Y
+ prbs_generator_syn_11/sky130_fd_sc_hs__nor2b_1_5/a_278_368# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_17/a_1178_124#
+ prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_39/X prbs_generator_syn_11/m3_13600_5433#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_63/a_437_503# prbs_generator_syn_11/sky130_fd_sc_hs__nand2_2_5/B
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_23/a_735_102# prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_53/A
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_61/a_735_102# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_57/a_1034_424#
+ prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_63/B prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_37/a_1141_508#
+ prbs_generator_syn_11/sky130_fd_sc_hs__nand2_1_47/B prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_29/X
+ prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_65/Y prbs_generator_syn_11/m3_13600_4701#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_1/a_437_503# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_67/a_1178_124#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_9/a_735_102# prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_13/a_132_392#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_15/a_1178_124# prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_15/A
+ prbs_generator_syn_11/sky130_fd_sc_hs__nand2_1_1/B prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_43/B
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_35/a_651_503# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_8/D
+ prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_29/A prbs_generator_syn_11/sky130_fd_sc_hs__nand2_1_7/B
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_13/a_735_102# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_47/a_696_458#
+ prbs_generator_syn_11/sky130_fd_sc_hs__nand2_1_31/B prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_51/a_735_102#
+ prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_59/X prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_35/a_1141_508#
+ prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_25/a_222_392# prbs_generator_syn_11/sky130_fd_sc_hs__sdlclkp_2_1/a_288_48#
+ prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_55/B prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_17/B
+ prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_43/A prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_7/A
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_65/a_1178_124# prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_59/Y
+ prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_41/X prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_21/a_230_79#
+ prbs_generator_syn_11/sky130_fd_sc_hs__nand2_1_57/a_117_74# prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_1/a_222_392#
+ prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_19/B prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_35/a_293_74#
+ prbs_generator_syn_11/sky130_fd_sc_hs__nand2_1_23/a_117_74# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_73/a_206_368#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_25/a_651_503# prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_1/a_138_385#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_37/a_696_458# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_67/a_544_485#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_43/a_27_74# prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_9/X
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_55/a_1034_424# prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_39/a_112_119#
+ prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_15/a_222_392# prbs_generator_syn_11/sky130_fd_sc_hs__conb_1_1/HI
+ prbs_generator_syn_11/sky130_fd_sc_hs__nand2_1_23/B prbs_generator_syn_11/sky130_fd_sc_hs__nand2_1_53/B
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_9/a_1178_124# prbs_generator_syn_11/sky130_fd_sc_hs__nor2b_1_4/A
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_47/a_1226_296# prbs_generator_syn_11/m3_13600_11045#
+ prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_17/X prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_29/a_376_368#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_5/a_544_485# prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_3/X
+ prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_31/a_132_392# prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_61/A
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_15/a_651_503# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_73/a_437_503#
+ prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_25/a_230_79# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_27/a_696_458#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_65/a_696_458# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_33/a_735_102#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_71/a_735_102# prbs_generator_syn_11/m3_13600_7263#
+ prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_43/a_222_392# prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_50/Y
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_8/a_1178_124# prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_53/B
+ prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_19/a_376_368# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_63/a_1178_124#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_4/a_696_458# prbs_generator_syn_11/sky130_fd_sc_hs__nor2b_1_4/a_278_368#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_13/a_1178_124# prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_61/a_132_392#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_53/a_206_368# prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_21/a_52_123#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_45/a_651_503# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_17/a_696_458#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_47/a_544_485# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_55/a_696_458#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_21/a_735_102# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_37/a_27_74#
+ prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_61/B prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_61/X
+ prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_59/a_112_119# prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_31/A
+ prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_33/a_222_392# prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_29/a_230_79#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_45/a_1226_296# prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_9/a_132_392#
+ prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_5/A prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_57/Y
+ prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_31/X prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_51/a_27_74#
+ prbs_generator_syn_11/sky130_fd_sc_hs__nor2b_1_8/a_27_112# prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_47/a_376_368#
+ prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_53/a_293_74# prbs_generator_syn_11/sky130_fd_sc_hs__nand2_1_43/a_117_74#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_8/a_735_102# prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_21/a_293_74#
+ prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_39/a_138_385# prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_63/Y
+ prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_51/a_132_392# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_43/a_206_368#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_53/a_437_503# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_37/a_544_485#
+ prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_57/X prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_53/a_1034_424#
+ prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_25/a_52_123# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_33/a_1141_508#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_63/Q prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_23/a_222_392#
+ prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_63/a_222_392# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_7/a_1178_124#
+ prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_53/X prbs_generator_syn_11/sky130_fd_sc_hs__nand2_2_5/Y
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_61/a_1178_124# prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_1/a_230_79#
+ prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_43/a_230_79# prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_11/a_230_79#
+ prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_41/a_132_392# prbs_generator_syn_11/sky130_fd_sc_hs__nand2_1_13/a_117_74#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_43/a_437_503# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_27/a_544_485#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_63/a_651_503# prbs_generator_syn_11/sky130_fd_sc_hs__nand2_1_7/a_117_74#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_35/a_696_458# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_65/a_544_485#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_51/a_1034_424# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_41/a_735_102#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_32/a_1141_508# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_49/a_1141_508#
+ prbs_generator_syn_11/sky130_fd_sc_hs__nand2_1_55/B prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_53/a_222_392#
+ prbs_generator_syn_11/sky130_fd_sc_hs__sdlclkp_2_1/a_114_112# prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_9/a_293_74#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_43/a_1226_296# prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_29/a_52_123#
+ prbs_generator_syn_11/sky130_fd_sc_hs__nand2_1_37/B prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_1/a_651_503#
+ prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_27/a_376_368# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_4/a_544_485#
+ prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_67/a_376_368# prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_27/X
+ prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_1/X prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_59/a_138_385#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_29/a_1178_124# prbs_generator_syn_11/m3_13600_2871#
+ prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_5/a_230_79# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_23/a_206_368#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_61/a_206_368# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_17/a_544_485#
+ prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_15/a_230_79# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_25/a_696_458#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_55/a_544_485# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_32/a_735_102#
+ prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_29/a_293_74# prbs_generator_syn_11/sky130_fd_sc_hs__nand2_1_17/a_117_74#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_69/a_1034_424# prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_29/a_112_119#
+ prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_37/X prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_31/B
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_19/a_1034_424# prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_33/A
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_9/a_206_368# prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_57/a_376_368#
+ prbs_generator_syn_11/sky130_fd_sc_hs__sdlclkp_2_1/a_706_317# prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_11/B
+ prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_1/a_52_123# prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_39/B
+ prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_21/a_132_392# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_13/a_206_368#
+ prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_43/a_52_123# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_51/a_206_368#
+ prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_47/X prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_23/a_437_503#
+ prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_11/a_52_123# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_61/a_437_503#
+ prbs_generator_syn_11/sky130_fd_sc_hs__nor2b_1_7/Y prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_51/A
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_15/a_696_458# prbs_generator_syn_11/sky130_fd_sc_hs__nor2b_1_5/Y
+ prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_9/a_230_79# prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_25/X
+ prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_19/a_112_119# prbs_generator_syn_11/sky130_fd_sc_hs__nand2_1_45/B
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_5/a_1178_124# prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_19/a_230_79#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_41/a_1226_296# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_59/a_1226_296#
+ prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_63/a_230_79# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_51/Q
+ prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_7/a_132_392# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_9/a_437_503#
+ prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_46/a_376_368# prbs_generator_syn_11/sky130_fd_sc_hs__nand2_1_33/a_117_74#
+ prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_11/a_293_74# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_27/a_1178_124#
+ prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_11/a_132_392# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_13/a_437_503#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_51/a_437_503# prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_5/a_52_123#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_35/a_544_485# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_73/a_651_503#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_45/a_696_458# prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_15/a_52_123#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_47/a_1141_508# prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_47/a_112_119#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_4/a_1178_124# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_17/a_1034_424#
+ prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_23/B prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_37/a_376_368#
+ prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_15/B prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_7/Y
+ prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_29/a_138_385# prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_33/a_230_79#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_25/a_1178_124# prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_47/a_293_74#
+ prbs_generator_syn_11/sky130_fd_sc_hs__nand2_1_37/a_117_74# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_33/a_206_368#
+ prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_15/a_293_74# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_71/a_206_368#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_25/a_544_485# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_67/a_1034_424#
+ prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_13/a_222_392# prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_9/a_52_123#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_15/a_1034_424# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_57/a_1226_296#
+ prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_19/a_52_123# prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_23/X
+ prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_63/a_52_123# prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_19/a_138_385#
+ prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_9/a_376_368# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_21/a_206_368#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_33/a_437_503# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_71/a_437_503#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_53/a_651_503# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_15/a_544_485#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_63/a_696_458# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_65/a_1034_424#
+ prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_19/a_293_74# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_45/a_1141_508#
+ prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_27/a_112_119# prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_67/a_112_119#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_1/a_1178_124# prbs_generator_syn_11/sky130_fd_sc_hs__conb_1_1/a_21_290#
+ prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_63/a_293_74# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_8/a_206_368#
+ prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_17/a_376_368# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_63/a_27_74#
+ prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_21/A prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_55/a_376_368#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_1/a_696_458# prbs_generator_syn_11/sky130_fd_sc_hs__nor2b_1_1/a_278_368#
+ prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_47/a_138_385# prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_33/a_52_123#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_9/a_1034_424# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_21/a_437_503#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_1/a_27_74# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_43/a_651_503#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_1/Q prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_45/a_544_485#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_69/a_735_102# prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_57/a_112_119#
+ prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_31/a_222_392# prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_13/A
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_55/a_1226_296# prbs_generator_syn_11/sky130_fd_sc_hs__nand2_2_5/a_27_74#
+ prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_53/a_230_79# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_8/a_437_503#
+ prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_67/a_293_74# prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_33/a_293_74#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_7/a_735_102# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_23/a_1178_124#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_41/a_206_368# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_8/a_1034_424#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_63/a_1034_424# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_59/a_735_102#
+ prbs_generator_syn_11/sky130_fd_sc_hs__nand2_1_5/B prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_43/a_1141_508#
+ prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_46/a_112_119# prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_61/a_222_392#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_13/a_1034_424# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_73/a_1178_124#
+ prbs_generator_syn_11/sky130_fd_sc_hs__nand2_1_27/B prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_13/B
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_57/a_27_74# prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_57/a_230_79#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_21/a_1178_124# prbs_generator_syn_11/sky130_fd_sc_hs__nor2b_1_1/a_27_112#
+ prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_27/a_138_385# prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_23/a_230_79#
+ prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_67/a_138_385# prbs_generator_syn_11/sky130_fd_sc_hs__nand2_1_41/B
+ prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_9/a_222_392# prbs_generator_syn_11/sky130_fd_sc_hs__nand2_1_27/a_117_74#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_32/a_206_368# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_23/a_651_503#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_41/a_437_503# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_73/a_27_74#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_61/a_651_503# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_63/a_544_485#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_49/a_735_102# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_73/a_696_458#
+ prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_37/a_112_119# prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_51/a_222_392#
+ prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_43/X prbs_generator_syn_11/sky130_fd_sc_hs__nand2_2_1/B
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_9/a_651_503# prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_53/a_52_123#
+ prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_49/X prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_25/a_376_368#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_1/a_544_485# prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_65/a_376_368#
+ prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_57/a_138_385# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_27/a_27_74#
+ prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_39/a_132_392# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_7/a_1034_424#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_13/a_651_503# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_32/a_437_503#
+ prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_27/a_230_79# prbs_generator_syn_11/m3_13600_12265#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_51/a_651_503# prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_59/B
+ prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_47/A prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_61/a_1034_424#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_41/a_1141_508# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_59/a_1141_508#
+ prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_41/a_222_392# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_53/a_1226_296#
+ prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_3/A prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_71/a_1178_124#
+ prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_9/a_112_119# prbs_generator_syn_11/sky130_fd_sc_hs__nand2_1_3/a_117_74#
+ prbs_generator_syn_11/m3_13600_8483# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_39/a_1178_124#
+ prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_57/a_52_123# prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_46/a_138_385#
+ prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_23/a_52_123# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_67/a_27_74#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_53/a_696_458# prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_17/a_112_119#
+ prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_11/A prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_55/a_112_119#
+ prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_1/A prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_51/a_1226_296#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_29/a_1034_424# prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_59/A
+ prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_23/A prbs_generator_syn_11/sky130_fd_sc_hs__nand2_1_39/B
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_5/a_27_74# prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_57/a_293_74#
+ prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_37/a_138_385# prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_59/a_132_392#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_33/a_651_503# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_71/a_651_503#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_43/a_696_458# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_73/a_544_485#
+ prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_27/a_52_123# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_57/a_1141_508#
+ prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_21/a_222_392# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_35/a_27_74#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_69/a_1226_296# prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_37/B
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_19/a_1226_296# prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_35/a_376_368#
+ prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_47/a_230_79# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_37/a_1178_124#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_5/a_1034_424# prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_49/a_132_392#
+ prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_7/a_222_392# prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_27/a_293_74#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_21/a_651_503# prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_9/a_138_385#
+ prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_11/a_222_392# prbs_generator_syn_11/m3_13600_14095#
+ prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_50/A prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_27/a_1034_424#
+ prbs_generator_syn_11/sky130_fd_sc_hs__nand2_1_13/B prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_8/a_651_503#
+ prbs_generator_syn_11/m3_13600_9703# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_35/a_1178_124#
+ prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_17/a_138_385# prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_55/a_138_385#
+ prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_7/a_230_79# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_4/a_1034_424#
+ prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_7/a_376_368# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_69/a_206_368#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_23/a_696_458# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_53/a_544_485#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_39/a_735_102# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_61/a_696_458#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_55/a_1141_508# prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_25/a_112_119#
+ prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_65/a_112_119# prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_43/a_293_74#
+ prbs_generator_syn_11/sky130_fd_sc_hs__nand2_1_57/B prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_25/a_1034_424#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_7/a_206_368# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_17/a_1226_296#
+ prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_15/a_376_368# prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_53/a_376_368#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_9/a_696_458# prbs_generator_syn_11/m3_13600_431#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_45/a_27_74# prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_47/a_52_123#
+ prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_29/a_132_392# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_59/a_206_368#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_69/a_437_503# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_41/a_651_503#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_43/a_544_485# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_13/a_696_458#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_29/a_735_102# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_51/a_696_458#
+ prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_61/Y prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_67/a_1226_296#
+ prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_5/a_132_392# prbs_generator_syn_11/sky130_fd_sc_hs__and2b_2_1/a_198_48#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_7/a_437_503# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_15/a_1226_296#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_69/a_27_74# prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_46/a_293_74#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_1/a_1034_424# prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_19/a_132_392#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_49/a_206_368# prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_7/a_52_123#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_59/a_437_503# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_32/a_651_503#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_7/a_27_74# prbs_generator_syn_11/sky130_fd_sc_hs__nand2_2_1/a_27_74#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_19/a_735_102# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_57/a_735_102#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_65/a_1226_296# prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_37/A
+ prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_33/a_376_368# prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_37/a_230_79#
+ prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_25/a_138_385# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_39/a_27_74#
+ prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_65/a_138_385# prbs_generator_syn_11/sky130_fd_sc_hs__nor2b_1_9/a_278_368#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_49/a_437_503# prbs_generator_syn_11/sky130_fd_sc_hs__and2b_2_1/a_505_74#
+ prbs_generator_syn_11/sky130_fd_sc_hs__nand2_1_51/a_117_74# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_23/a_544_485#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_33/a_696_458# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_61/a_544_485#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_9/a_1226_296# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_53/a_1141_508#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_71/a_696_458# prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_35/a_112_119#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_23/a_1034_424# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_9/a_544_485#
+ prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_63/a_376_368# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_33/a_1178_124#
+ prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_5/a_376_368# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_13/a_544_485#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_73/a_1034_424# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_21/a_696_458#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_51/a_544_485# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_8/a_1226_296#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_51/a_1141_508# prbs_generator_syn_11/sky130_fd_sc_hs__nand2_1_55/a_117_74#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_21/a_1034_424# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_63/a_1226_296#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_23/a_27_74# prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_7/a_112_119#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_13/a_1226_296# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_8/a_696_458#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_32/a_1178_124# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_49/a_1178_124#
+ prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_37/a_52_123# prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_27/a_132_392#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_71/Q prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_67/a_735_102#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_69/a_1141_508# prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_15/a_112_119#
+ prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_53/a_112_119# prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_39/a_222_392#
+ prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_55/a_230_79# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_19/a_1141_508#
+ prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_37/a_293_74# prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_43/a_376_368#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_5/a_735_102# prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_35/a_138_385#
+ prbs_generator_syn_11/sky130_fd_sc_hs__sdlclkp_2_1/a_114_424# prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_57/a_132_392#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_71/a_1034_424# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_7/a_1226_296#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_33/a_544_485# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_41/a_696_458#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_71/a_544_485# prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_21/B
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_61/a_1226_296# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_39/a_1034_424#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_17/a_27_74# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_9/a_27_74#
+ prbs_generator_syn_11/sky130_fd_sc_hs__nor2b_1_5/a_27_112# prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_47/a_132_392#
+ prbs_generator_syn_11/sky130_fd_sc_hs__nor2b_1_8/a_278_368# prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_9/B
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_39/a_206_368# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_33/a_27_74#
+ prbs_generator_syn_11/sky130_fd_sc_hs__nand2_1_41/a_117_74# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_69/a_651_503#
+ prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_51/a_293_74# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_21/a_544_485#
+ prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_7/a_138_385# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_32/a_696_458#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_47/a_735_102# prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_33/a_112_119#
+ prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_59/a_222_392# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_17/a_1141_508#
+ prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_55/a_52_123# prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_3/a_293_74#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_7/a_651_503# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_29/a_1226_296#
+ prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_23/a_376_368# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_8/a_544_485#
+ prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_47/B prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_47/a_1178_124#
+ prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_15/a_138_385# prbs_generator_syn_11/sky130_fd_sc_hs__sdlclkp_2_1/a_1195_374#
+ prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_53/a_138_385# prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_37/a_132_392#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_29/a_206_368# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_39/a_437_503#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_59/a_651_503# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_37/a_735_102#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_67/a_1141_508# prbs_generator_syn_11/sky130_fd_sc_hs__and2b_2_1/a_27_74#
+ prbs_generator_syn_11/sky130_fd_sc_hs__conb_1_1/a_165_290# prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_55/a_293_74#
+ prbs_generator_syn_11/sky130_fd_sc_hs__nand2_1_45/a_117_74# prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_63/a_112_119#
+ prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_49/a_222_392# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_37/a_1034_424#
+ prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_23/a_293_74# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_15/a_1141_508#
+ prbs_generator_syn_11/sky130_fd_sc_hs__nand2_1_5/a_117_74# prbs_generator_syn_11/m3_13600_13485#
+ prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_5/a_112_119# prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_13/a_376_368#
+ prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_51/a_376_368# prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_7/a_293_74#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_19/a_206_368# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_57/a_206_368#
+ prbs_generator_syn_11/sky130_fd_sc_hs__sdlclkp_2_1/a_318_74# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_29/a_437_503#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_49/a_651_503# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_25/a_27_74#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_5/a_1226_296# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_41/a_544_485#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_27/a_735_102# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_65/a_1141_508#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_65/a_735_102# prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_3/a_230_79#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_35/a_1034_424# prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_13/a_230_79#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_41/a_27_74# prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_3/a_132_392#
+ prbs_generator_syn_11/sky130_fd_sc_hs__nand2_1_49/a_117_74# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_27/a_1226_296#
+ prbs_generator_syn_11/sky130_fd_sc_hs__nand2_1_15/a_117_74# prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_41/a_376_368#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_45/a_1178_124# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_4/a_735_102#
+ prbs_generator_syn_11/sky130_fd_sc_hs__nand2_1_9/a_117_74# prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_33/a_138_385#
+ prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_17/a_132_392# prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_55/a_132_392#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_9/a_1141_508# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_19/a_437_503#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_57/a_437_503# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_4/a_1226_296#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_32/a_544_485# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_17/a_735_102#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_55/a_735_102# prbs_generator_syn_11/m3_13600_2261#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_65/a_27_74# prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_29/a_222_392#
+ prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_43/a_112_119# prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_19/X
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_25/a_1226_296# prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_31/a_376_368#
+ prbs_generator_syn_11/sky130_fd_sc_hs__or2_1_1/a_63_368# prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_17/a_230_79#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_4/a_27_74# prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_61/a_230_79#
+ prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_63/a_138_385# prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_5/a_222_392#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_8/a_1141_508# prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_41/a_293_74#
+ prbs_generator_syn_11/sky130_fd_sc_hs__nand2_1_31/a_117_74# prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_5/a_138_385#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_63/a_1141_508# prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_19/a_222_392#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_13/a_1141_508# prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_3/a_52_123#
+ prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_13/a_52_123# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_43/a_1178_124#
+ prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_61/a_376_368# prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_35/a_132_392#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_67/a_206_368# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_1/a_1226_296#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_69/a_696_458# prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_31/a_230_79#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_35/a_735_102# prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_23/a_112_119#
+ prbs_generator_syn_11/sky130_fd_sc_hs__nand2_1_35/a_117_74# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_59/a_27_74#
+ prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_13/a_293_74# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_5/a_206_368#
+ prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_50/a_376_368# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_7/a_696_458#
+ prbs_generator_syn_11/sky130_fd_sc_hs__nor2b_1_7/a_278_368# prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_17/a_52_123#
+ prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_43/a_138_385# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_7/a_1141_508#
+ prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_61/a_52_123# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_67/a_437_503#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_61/a_1141_508# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_25/a_735_102#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_59/a_696_458# prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_13/a_112_119#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_33/a_1034_424# prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_51/a_112_119#
+ prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_35/a_230_79# prbs_generator_syn_11/m3_13600_4091#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_23/a_1226_296# prbs_generator_syn_11/sky130_fd_sc_hs__nand2_1_39/a_117_74#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_29/a_27_74# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_5/a_437_503#
+ prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_17/a_293_74# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_41/a_1178_124#
+ prbs_generator_syn_11/sky130_fd_sc_hs__or2_1_1/a_152_368# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_59/a_1178_124#
+ prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_61/a_293_74# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_47/a_206_368#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_39/a_651_503# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_49/a_696_458#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_15/a_735_102# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_32/a_1034_424#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_73/a_1226_296# prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_27/a_222_392#
+ prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_41/a_112_119# prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_31/a_52_123#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_49/a_1034_424# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_29/a_1141_508#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_21/a_1226_296# prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_39/a_230_79#
+ prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_23/a_138_385# prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_51/a_230_79#
+ prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_45/a_132_392# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_37/a_206_368#
+ prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_65/a_293_74# prbs_generator_syn_11/sky130_fd_sc_hs__nand2_1_53/a_117_74#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_47/a_437_503# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_29/a_651_503#
+ prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_31/a_293_74# prbs_generator_syn_11/sky130_fd_sc_hs__nand2_1_21/a_117_74#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_69/a_544_485# prbs_generator_syn_11/sky130_fd_sc_hs__clkbuf_16_1/a_114_74#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_45/a_735_102# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_13/a_27_74#
+ prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_31/a_112_119# prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_57/a_222_392#
+ prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_35/a_52_123# prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_21/a_376_368#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_7/a_544_485# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_57/a_1178_124#
+ prbs_generator_syn_11/m3_13600_6043# prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_13/a_138_385#
+ prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_51/a_138_385# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_5/a_1141_508#
+ prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_3/a_376_368# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_27/a_206_368#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_65/a_206_368# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_37/a_437_503#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_19/a_651_503# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_57/a_651_503#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_59/a_544_485# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_71/a_1226_296#
+ prbs_generator_syn_11/sky130_fd_sc_hs__nand2_1_25/a_117_74# prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_61/a_112_119#
+ prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_47/a_222_392# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_27/a_1141_508#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_53/a_27_74# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_4/a_206_368#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_39/a_1226_296# prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_11/a_376_368#
+ prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_39/a_52_123# prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_41/a_138_385#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_4/a_1141_508# prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_25/a_132_392#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_17/a_206_368# prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_41/A
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_55/a_206_368# prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_51/a_52_123#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_27/a_437_503# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_65/a_437_503#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_49/a_544_485# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_63/a_735_102#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_47/a_1034_424# prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_50/a_112_119#
+ prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_37/a_222_392# prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_59/a_230_79#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_25/a_1141_508# prbs_generator_syn_11/sky130_fd_sc_hs__nor2b_1_4/a_27_112#
+ prbs_generator_syn_11/sky130_fd_sc_hs__sdlclkp_2_1/a_685_81# prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_1/a_132_392#
+ prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_39/a_293_74# prbs_generator_syn_11/sky130_fd_sc_hs__nand2_1_29/a_117_74#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_4/a_437_503# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_55/a_1178_124#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_21/a_27_74# prbs_generator_syn_11/m3_13600_12875#
+ prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_50/a_293_74# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_1/a_735_102#
+ prbs_generator_syn_11/sky130_fd_sc_hs__xnor2_1_31/a_138_385# prbs_generator_syn_11/sky130_fd_sc_hs__a22o_1_15/a_132_392#
+ prbs_generator_syn_11/sky130_fd_sc_hs__nand2_1_1/a_117_74# prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_17/a_437_503#
+ prbs_generator_syn_11/sky130_fd_sc_hs__dfxtp_4_55/a_437_503# prbs_generator_syn
Xprbs_generator_syn_22 prbs_generator_syn_31/clk prbs_generator_syn_31/rst prbs_generator_syn_23/cke
+ sky130_fd_sc_hs__conb_1_231/LO sky130_fd_sc_hs__conb_1_231/LO sky130_fd_sc_hs__conb_1_231/HI
+ prbs_generator_syn_27/eqn[1] prbs_generator_syn_27/eqn[8] sky130_fd_sc_hs__conb_1_231/LO
+ sky130_fd_sc_hs__conb_1_231/LO sky130_fd_sc_hs__conb_1_231/LO sky130_fd_sc_hs__conb_1_231/LO
+ sky130_fd_sc_hs__conb_1_231/LO sky130_fd_sc_hs__conb_1_231/LO prbs_generator_syn_23/eqn[31]
+ prbs_generator_syn_23/cke prbs_generator_syn_23/eqn[31] sky130_fd_sc_hs__conb_1_233/HI
+ sky130_fd_sc_hs__conb_1_233/HI sky130_fd_sc_hs__conb_1_233/HI prbs_generator_syn_27/eqn[9]
+ sky130_fd_sc_hs__conb_1_187/HI prbs_generator_syn_29/eqn[22] prbs_generator_syn_29/eqn[20]
+ prbs_generator_syn_29/eqn[22] prbs_generator_syn_29/eqn[20] sky130_fd_sc_hs__conb_1_191/HI
+ prbs_generator_syn_29/eqn[28] sky130_fd_sc_hs__conb_1_191/HI prbs_generator_syn_29/eqn[28]
+ prbs_generator_syn_29/cke prbs_generator_syn_29/eqn[31] prbs_generator_syn_29/cke
+ prbs_generator_syn_29/eqn[31] prbs_generator_syn_29/cke prbs_generator_syn_23/eqn[31]
+ prbs_generator_syn_23/eqn[30] prbs_generator_syn_23/eqn[30] prbs_generator_syn_23/eqn[28]
+ prbs_generator_syn_23/eqn[28] prbs_generator_syn_23/eqn[28] prbs_generator_syn_23/eqn[28]
+ prbs_generator_syn_23/eqn[28] prbs_generator_syn_23/eqn[28] prbs_generator_syn_23/eqn[22]
+ prbs_generator_syn_23/eqn[22] prbs_generator_syn_23/eqn[20] prbs_generator_syn_23/eqn[22]
+ prbs_generator_syn_23/eqn[22] prbs_generator_syn_23/eqn[22] prbs_generator_syn_23/eqn[22]
+ prbs_generator_syn_21/eqn[0] prbs_generator_syn_21/eqn[0] prbs_generator_syn_21/eqn[0]
+ prbs_generator_syn_21/eqn[0] prbs_generator_syn_21/eqn[0] prbs_generator_syn_21/eqn[0]
+ prbs_generator_syn_23/eqn[9] prbs_generator_syn_23/eqn[8] prbs_generator_syn_23/eqn[8]
+ prbs_generator_syn_23/eqn[8] prbs_generator_syn_23/eqn[8] prbs_generator_syn_23/eqn[8]
+ prbs_generator_syn_23/eqn[8] prbs_generator_syn_23/eqn[8] prbs_generator_syn_23/eqn[1]
+ prbs_generator_syn_23/eqn[0] prbs_generator_syn_31/inj_err prbs_generator_syn_23/eqn[31]
+ prbs_generator_syn_23/eqn[31] hr_16t4_mux_top_1/din[2] DVSS: DVDD: prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_1/a_293_74#
+ prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_15/X prbs_generator_syn_23/sky130_fd_sc_hs__nand2_1_35/B
+ prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_51/Y prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_9/A
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_9/CLK prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_47/a_27_74#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_37/a_1226_296# prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_3/B
+ prbs_generator_syn_23/sky130_fd_sc_hs__nor2b_1_7/a_27_112# prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_29/B
+ prbs_generator_syn_23/sky130_fd_sc_hs__sdlclkp_2_1/a_580_74# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_1/a_1141_508#
+ prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_5/Y prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_41/a_230_79#
+ prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_61/a_138_385# prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_43/a_132_392#
+ prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_3/a_222_392# prbs_generator_syn_23/sky130_fd_sc_hs__nor2b_1_9/a_27_112#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_61/a_27_74# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_35/a_206_368#
+ prbs_generator_syn_23/sky130_fd_sc_hs__nand2_2_3/Y prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_25/B
+ prbs_generator_syn_23/sky130_fd_sc_hs__nand2_1_11/a_117_74# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_67/a_651_503#
+ prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_45/X prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_39/a_696_458#
+ prbs_generator_syn_23/sky130_fd_sc_hs__sdlclkp_2_1/a_1198_74# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_45/a_1034_424#
+ prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_17/a_222_392# prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_55/a_222_392#
+ prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_53/Y prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_35/A
+ prbs_generator_syn_23/m3_13600_1651# prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_59/a_52_123#
+ prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_5/a_293_74# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_35/a_1226_296#
+ prbs_generator_syn_23/sky130_fd_sc_hs__nand2_1_51/B prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_5/a_651_503#
+ prbs_generator_syn_23/sky130_fd_sc_hs__nand2_1_21/B prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_8/a_27_74#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_15/a_27_74# prbs_generator_syn_23/sky130_fd_sc_hs__and2b_2_1/X
+ prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_13/X prbs_generator_syn_23/sky130_fd_sc_hs__nand2_2_3/a_27_74#
+ prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_50/a_138_385# prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_33/a_132_392#
+ prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_1/a_376_368# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_25/a_206_368#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_35/a_437_503# prbs_generator_syn_23/sky130_fd_sc_hs__sdlclkp_2_1/a_708_451#
+ prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_45/a_230_79# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_29/a_696_458#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_32/a_27_74# prbs_generator_syn_23/sky130_fd_sc_hs__nor2b_1_4/Y
+ prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_59/a_293_74# prbs_generator_syn_23/sky130_fd_sc_hs__nand2_1_47/a_117_74#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_73/a_735_102# prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_21/a_112_119#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_23/a_1141_508# prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_25/a_293_74#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_7/Q prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_3/a_112_119#
+ prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_35/B prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_51/X
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_53/a_1178_124# prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_23/a_132_392#
+ prbs_generator_syn_23/sky130_fd_sc_hs__nand2_1_3/B prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_15/a_206_368#
+ prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_63/a_132_392# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_55/a_27_74#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_25/a_437_503# prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_41/a_52_123#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_47/a_651_503# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_73/a_1141_508#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_19/a_696_458# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_57/a_696_458#
+ prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_7/X prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_43/a_1034_424#
+ prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_55/A prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_11/a_112_119#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_21/a_1141_508# prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_35/a_222_392#
+ prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_49/a_230_79# prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_67/Y
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_71/a_27_74# prbs_generator_syn_23/sky130_fd_sc_hs__nand2_1_33/B
+ prbs_generator_syn_23/sky130_fd_sc_hs__conb_1_1/LO prbs_generator_syn_23/sky130_fd_sc_hs__nand2_1_19/a_117_74#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_51/a_1178_124# prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_33/X
+ prbs_generator_syn_23/sky130_fd_sc_hs__nand2_1_29/B prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_41/Y
+ prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_53/a_132_392# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_45/a_206_368#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_15/a_437_503# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_37/a_651_503#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_39/a_544_485# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_53/a_735_102#
+ prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_45/a_52_123# prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_1/B
+ prbs_generator_syn_23/sky130_fd_sc_hs__nand2_2_3/B prbs_generator_syn_23/sky130_fd_sc_hs__clkbuf_16_1/A
+ prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_21/X prbs_generator_syn_23/sky130_fd_sc_hs__nand2_1_25/B
+ prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_39/a_376_368# prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_63/X
+ prbs_generator_syn_23/m3_13600_3481# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_69/a_1178_124#
+ prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_21/a_138_385# prbs_generator_syn_23/sky130_fd_sc_hs__nor2b_1_8/Y
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_19/a_1178_124# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_49/a_27_74#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_45/a_437_503# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_27/a_651_503#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_71/a_1141_508# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_65/a_651_503#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_29/a_544_485# prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_3/a_138_385#
+ prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_55/X prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_43/a_735_102#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_41/a_1034_424# prbs_generator_syn_23/sky130_fd_sc_hs__nand2_1_9/B
+ prbs_generator_syn_23/sky130_fd_sc_hs__nor2b_1_9/Y prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_59/a_1034_424#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_39/a_1141_508# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_33/a_1226_296#
+ prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_49/a_52_123# prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_47/Y
+ prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_43/Y prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_4/a_651_503#
+ prbs_generator_syn_23/sky130_fd_sc_hs__nand2_1_49/B prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_19/A
+ prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_11/a_138_385# prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_5/X
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_63/a_206_368# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_17/a_651_503#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_19/a_544_485# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_55/a_651_503#
+ prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_9/Y prbs_generator_syn_23/sky130_fd_sc_hs__nand2_1_17/B
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_57/a_544_485# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_67/a_696_458#
+ prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_35/X prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_19/a_27_74#
+ prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_45/a_222_392# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_32/a_1226_296#
+ prbs_generator_syn_23/sky130_fd_sc_hs__nand2_1_43/B prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_25/A
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_1/a_206_368# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_49/a_1226_296#
+ prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_1/a_112_119# prbs_generator_syn_23/sky130_fd_sc_hs__or2_1_1/X
+ prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_59/a_376_368# prbs_generator_syn_23/sky130_fd_sc_hs__nand2_1_19/B
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_5/a_696_458# prbs_generator_syn_23/sky130_fd_sc_hs__nor2b_1_1/Y
+ prbs_generator_syn_23/sky130_fd_sc_hs__nor2b_1_5/a_278_368# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_17/a_1178_124#
+ prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_39/X prbs_generator_syn_23/m3_13600_5433#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_63/a_437_503# prbs_generator_syn_23/sky130_fd_sc_hs__nand2_2_5/B
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_23/a_735_102# prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_53/A
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_61/a_735_102# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_57/a_1034_424#
+ prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_63/B prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_37/a_1141_508#
+ prbs_generator_syn_23/sky130_fd_sc_hs__nand2_1_47/B prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_29/X
+ prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_65/Y prbs_generator_syn_23/m3_13600_4701#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_1/a_437_503# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_67/a_1178_124#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_9/a_735_102# prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_13/a_132_392#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_15/a_1178_124# prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_15/A
+ prbs_generator_syn_23/sky130_fd_sc_hs__nand2_1_1/B prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_43/B
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_35/a_651_503# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_8/D
+ prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_29/A prbs_generator_syn_23/sky130_fd_sc_hs__nand2_1_7/B
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_13/a_735_102# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_47/a_696_458#
+ prbs_generator_syn_23/sky130_fd_sc_hs__nand2_1_31/B prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_51/a_735_102#
+ prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_59/X prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_35/a_1141_508#
+ prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_25/a_222_392# prbs_generator_syn_23/sky130_fd_sc_hs__sdlclkp_2_1/a_288_48#
+ prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_55/B prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_17/B
+ prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_43/A prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_7/A
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_65/a_1178_124# prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_59/Y
+ prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_41/X prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_21/a_230_79#
+ prbs_generator_syn_23/sky130_fd_sc_hs__nand2_1_57/a_117_74# prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_1/a_222_392#
+ prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_19/B prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_35/a_293_74#
+ prbs_generator_syn_23/sky130_fd_sc_hs__nand2_1_23/a_117_74# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_73/a_206_368#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_25/a_651_503# prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_1/a_138_385#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_37/a_696_458# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_67/a_544_485#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_43/a_27_74# prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_9/X
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_55/a_1034_424# prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_39/a_112_119#
+ prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_15/a_222_392# prbs_generator_syn_23/sky130_fd_sc_hs__conb_1_1/HI
+ prbs_generator_syn_23/sky130_fd_sc_hs__nand2_1_23/B prbs_generator_syn_23/sky130_fd_sc_hs__nand2_1_53/B
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_9/a_1178_124# prbs_generator_syn_23/sky130_fd_sc_hs__nor2b_1_4/A
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_47/a_1226_296# prbs_generator_syn_23/m3_13600_11045#
+ prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_17/X prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_29/a_376_368#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_5/a_544_485# prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_3/X
+ prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_31/a_132_392# prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_61/A
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_15/a_651_503# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_73/a_437_503#
+ prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_25/a_230_79# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_27/a_696_458#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_65/a_696_458# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_33/a_735_102#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_71/a_735_102# prbs_generator_syn_23/m3_13600_7263#
+ prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_43/a_222_392# prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_50/Y
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_8/a_1178_124# prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_53/B
+ prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_19/a_376_368# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_63/a_1178_124#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_4/a_696_458# prbs_generator_syn_23/sky130_fd_sc_hs__nor2b_1_4/a_278_368#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_13/a_1178_124# prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_61/a_132_392#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_53/a_206_368# prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_21/a_52_123#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_45/a_651_503# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_17/a_696_458#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_47/a_544_485# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_55/a_696_458#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_21/a_735_102# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_37/a_27_74#
+ prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_61/B prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_61/X
+ prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_59/a_112_119# prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_31/A
+ prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_33/a_222_392# prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_29/a_230_79#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_45/a_1226_296# prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_9/a_132_392#
+ prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_5/A prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_57/Y
+ prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_31/X prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_51/a_27_74#
+ prbs_generator_syn_23/sky130_fd_sc_hs__nor2b_1_8/a_27_112# prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_47/a_376_368#
+ prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_53/a_293_74# prbs_generator_syn_23/sky130_fd_sc_hs__nand2_1_43/a_117_74#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_8/a_735_102# prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_21/a_293_74#
+ prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_39/a_138_385# prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_63/Y
+ prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_51/a_132_392# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_43/a_206_368#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_53/a_437_503# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_37/a_544_485#
+ prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_57/X prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_53/a_1034_424#
+ prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_25/a_52_123# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_33/a_1141_508#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_63/Q prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_23/a_222_392#
+ prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_63/a_222_392# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_7/a_1178_124#
+ prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_53/X prbs_generator_syn_23/sky130_fd_sc_hs__nand2_2_5/Y
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_61/a_1178_124# prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_1/a_230_79#
+ prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_43/a_230_79# prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_11/a_230_79#
+ prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_41/a_132_392# prbs_generator_syn_23/sky130_fd_sc_hs__nand2_1_13/a_117_74#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_43/a_437_503# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_27/a_544_485#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_63/a_651_503# prbs_generator_syn_23/sky130_fd_sc_hs__nand2_1_7/a_117_74#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_35/a_696_458# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_65/a_544_485#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_51/a_1034_424# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_41/a_735_102#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_32/a_1141_508# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_49/a_1141_508#
+ prbs_generator_syn_23/sky130_fd_sc_hs__nand2_1_55/B prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_53/a_222_392#
+ prbs_generator_syn_23/sky130_fd_sc_hs__sdlclkp_2_1/a_114_112# prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_9/a_293_74#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_43/a_1226_296# prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_29/a_52_123#
+ prbs_generator_syn_23/sky130_fd_sc_hs__nand2_1_37/B prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_1/a_651_503#
+ prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_27/a_376_368# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_4/a_544_485#
+ prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_67/a_376_368# prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_27/X
+ prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_1/X prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_59/a_138_385#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_29/a_1178_124# prbs_generator_syn_23/m3_13600_2871#
+ prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_5/a_230_79# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_23/a_206_368#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_61/a_206_368# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_17/a_544_485#
+ prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_15/a_230_79# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_25/a_696_458#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_55/a_544_485# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_32/a_735_102#
+ prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_29/a_293_74# prbs_generator_syn_23/sky130_fd_sc_hs__nand2_1_17/a_117_74#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_69/a_1034_424# prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_29/a_112_119#
+ prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_37/X prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_31/B
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_19/a_1034_424# prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_33/A
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_9/a_206_368# prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_57/a_376_368#
+ prbs_generator_syn_23/sky130_fd_sc_hs__sdlclkp_2_1/a_706_317# prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_11/B
+ prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_1/a_52_123# prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_39/B
+ prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_21/a_132_392# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_13/a_206_368#
+ prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_43/a_52_123# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_51/a_206_368#
+ prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_47/X prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_23/a_437_503#
+ prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_11/a_52_123# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_61/a_437_503#
+ prbs_generator_syn_23/sky130_fd_sc_hs__nor2b_1_7/Y prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_51/A
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_15/a_696_458# prbs_generator_syn_23/sky130_fd_sc_hs__nor2b_1_5/Y
+ prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_9/a_230_79# prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_25/X
+ prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_19/a_112_119# prbs_generator_syn_23/sky130_fd_sc_hs__nand2_1_45/B
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_5/a_1178_124# prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_19/a_230_79#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_41/a_1226_296# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_59/a_1226_296#
+ prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_63/a_230_79# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_51/Q
+ prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_7/a_132_392# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_9/a_437_503#
+ prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_46/a_376_368# prbs_generator_syn_23/sky130_fd_sc_hs__nand2_1_33/a_117_74#
+ prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_11/a_293_74# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_27/a_1178_124#
+ prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_11/a_132_392# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_13/a_437_503#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_51/a_437_503# prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_5/a_52_123#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_35/a_544_485# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_73/a_651_503#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_45/a_696_458# prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_15/a_52_123#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_47/a_1141_508# prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_47/a_112_119#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_4/a_1178_124# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_17/a_1034_424#
+ prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_23/B prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_37/a_376_368#
+ prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_15/B prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_7/Y
+ prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_29/a_138_385# prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_33/a_230_79#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_25/a_1178_124# prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_47/a_293_74#
+ prbs_generator_syn_23/sky130_fd_sc_hs__nand2_1_37/a_117_74# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_33/a_206_368#
+ prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_15/a_293_74# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_71/a_206_368#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_25/a_544_485# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_67/a_1034_424#
+ prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_13/a_222_392# prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_9/a_52_123#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_15/a_1034_424# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_57/a_1226_296#
+ prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_19/a_52_123# prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_23/X
+ prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_63/a_52_123# prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_19/a_138_385#
+ prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_9/a_376_368# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_21/a_206_368#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_33/a_437_503# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_71/a_437_503#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_53/a_651_503# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_15/a_544_485#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_63/a_696_458# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_65/a_1034_424#
+ prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_19/a_293_74# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_45/a_1141_508#
+ prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_27/a_112_119# prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_67/a_112_119#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_1/a_1178_124# prbs_generator_syn_23/sky130_fd_sc_hs__conb_1_1/a_21_290#
+ prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_63/a_293_74# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_8/a_206_368#
+ prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_17/a_376_368# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_63/a_27_74#
+ prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_21/A prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_55/a_376_368#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_1/a_696_458# prbs_generator_syn_23/sky130_fd_sc_hs__nor2b_1_1/a_278_368#
+ prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_47/a_138_385# prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_33/a_52_123#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_9/a_1034_424# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_21/a_437_503#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_1/a_27_74# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_43/a_651_503#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_1/Q prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_45/a_544_485#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_69/a_735_102# prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_57/a_112_119#
+ prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_31/a_222_392# prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_13/A
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_55/a_1226_296# prbs_generator_syn_23/sky130_fd_sc_hs__nand2_2_5/a_27_74#
+ prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_53/a_230_79# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_8/a_437_503#
+ prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_67/a_293_74# prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_33/a_293_74#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_7/a_735_102# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_23/a_1178_124#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_41/a_206_368# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_8/a_1034_424#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_63/a_1034_424# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_59/a_735_102#
+ prbs_generator_syn_23/sky130_fd_sc_hs__nand2_1_5/B prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_43/a_1141_508#
+ prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_46/a_112_119# prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_61/a_222_392#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_13/a_1034_424# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_73/a_1178_124#
+ prbs_generator_syn_23/sky130_fd_sc_hs__nand2_1_27/B prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_13/B
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_57/a_27_74# prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_57/a_230_79#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_21/a_1178_124# prbs_generator_syn_23/sky130_fd_sc_hs__nor2b_1_1/a_27_112#
+ prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_27/a_138_385# prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_23/a_230_79#
+ prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_67/a_138_385# prbs_generator_syn_23/sky130_fd_sc_hs__nand2_1_41/B
+ prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_9/a_222_392# prbs_generator_syn_23/sky130_fd_sc_hs__nand2_1_27/a_117_74#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_32/a_206_368# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_23/a_651_503#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_41/a_437_503# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_73/a_27_74#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_61/a_651_503# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_63/a_544_485#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_49/a_735_102# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_73/a_696_458#
+ prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_37/a_112_119# prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_51/a_222_392#
+ prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_43/X prbs_generator_syn_23/sky130_fd_sc_hs__nand2_2_1/B
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_9/a_651_503# prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_53/a_52_123#
+ prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_49/X prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_25/a_376_368#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_1/a_544_485# prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_65/a_376_368#
+ prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_57/a_138_385# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_27/a_27_74#
+ prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_39/a_132_392# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_7/a_1034_424#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_13/a_651_503# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_32/a_437_503#
+ prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_27/a_230_79# prbs_generator_syn_23/m3_13600_12265#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_51/a_651_503# prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_59/B
+ prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_47/A prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_61/a_1034_424#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_41/a_1141_508# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_59/a_1141_508#
+ prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_41/a_222_392# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_53/a_1226_296#
+ prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_3/A prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_71/a_1178_124#
+ prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_9/a_112_119# prbs_generator_syn_23/sky130_fd_sc_hs__nand2_1_3/a_117_74#
+ prbs_generator_syn_23/m3_13600_8483# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_39/a_1178_124#
+ prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_57/a_52_123# prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_46/a_138_385#
+ prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_23/a_52_123# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_67/a_27_74#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_53/a_696_458# prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_17/a_112_119#
+ prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_11/A prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_55/a_112_119#
+ prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_1/A prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_51/a_1226_296#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_29/a_1034_424# prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_59/A
+ prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_23/A prbs_generator_syn_23/sky130_fd_sc_hs__nand2_1_39/B
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_5/a_27_74# prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_57/a_293_74#
+ prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_37/a_138_385# prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_59/a_132_392#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_33/a_651_503# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_71/a_651_503#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_43/a_696_458# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_73/a_544_485#
+ prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_27/a_52_123# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_57/a_1141_508#
+ prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_21/a_222_392# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_35/a_27_74#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_69/a_1226_296# prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_37/B
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_19/a_1226_296# prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_35/a_376_368#
+ prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_47/a_230_79# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_37/a_1178_124#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_5/a_1034_424# prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_49/a_132_392#
+ prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_7/a_222_392# prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_27/a_293_74#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_21/a_651_503# prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_9/a_138_385#
+ prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_11/a_222_392# prbs_generator_syn_23/m3_13600_14095#
+ prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_50/A prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_27/a_1034_424#
+ prbs_generator_syn_23/sky130_fd_sc_hs__nand2_1_13/B prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_8/a_651_503#
+ prbs_generator_syn_23/m3_13600_9703# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_35/a_1178_124#
+ prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_17/a_138_385# prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_55/a_138_385#
+ prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_7/a_230_79# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_4/a_1034_424#
+ prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_7/a_376_368# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_69/a_206_368#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_23/a_696_458# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_53/a_544_485#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_39/a_735_102# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_61/a_696_458#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_55/a_1141_508# prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_25/a_112_119#
+ prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_65/a_112_119# prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_43/a_293_74#
+ prbs_generator_syn_23/sky130_fd_sc_hs__nand2_1_57/B prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_25/a_1034_424#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_7/a_206_368# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_17/a_1226_296#
+ prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_15/a_376_368# prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_53/a_376_368#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_9/a_696_458# prbs_generator_syn_23/m3_13600_431#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_45/a_27_74# prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_47/a_52_123#
+ prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_29/a_132_392# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_59/a_206_368#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_69/a_437_503# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_41/a_651_503#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_43/a_544_485# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_13/a_696_458#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_29/a_735_102# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_51/a_696_458#
+ prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_61/Y prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_67/a_1226_296#
+ prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_5/a_132_392# prbs_generator_syn_23/sky130_fd_sc_hs__and2b_2_1/a_198_48#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_7/a_437_503# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_15/a_1226_296#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_69/a_27_74# prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_46/a_293_74#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_1/a_1034_424# prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_19/a_132_392#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_49/a_206_368# prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_7/a_52_123#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_59/a_437_503# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_32/a_651_503#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_7/a_27_74# prbs_generator_syn_23/sky130_fd_sc_hs__nand2_2_1/a_27_74#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_19/a_735_102# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_57/a_735_102#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_65/a_1226_296# prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_37/A
+ prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_33/a_376_368# prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_37/a_230_79#
+ prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_25/a_138_385# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_39/a_27_74#
+ prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_65/a_138_385# prbs_generator_syn_23/sky130_fd_sc_hs__nor2b_1_9/a_278_368#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_49/a_437_503# prbs_generator_syn_23/sky130_fd_sc_hs__and2b_2_1/a_505_74#
+ prbs_generator_syn_23/sky130_fd_sc_hs__nand2_1_51/a_117_74# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_23/a_544_485#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_33/a_696_458# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_61/a_544_485#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_9/a_1226_296# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_53/a_1141_508#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_71/a_696_458# prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_35/a_112_119#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_23/a_1034_424# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_9/a_544_485#
+ prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_63/a_376_368# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_33/a_1178_124#
+ prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_5/a_376_368# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_13/a_544_485#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_73/a_1034_424# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_21/a_696_458#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_51/a_544_485# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_8/a_1226_296#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_51/a_1141_508# prbs_generator_syn_23/sky130_fd_sc_hs__nand2_1_55/a_117_74#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_21/a_1034_424# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_63/a_1226_296#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_23/a_27_74# prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_7/a_112_119#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_13/a_1226_296# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_8/a_696_458#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_32/a_1178_124# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_49/a_1178_124#
+ prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_37/a_52_123# prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_27/a_132_392#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_71/Q prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_67/a_735_102#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_69/a_1141_508# prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_15/a_112_119#
+ prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_53/a_112_119# prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_39/a_222_392#
+ prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_55/a_230_79# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_19/a_1141_508#
+ prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_37/a_293_74# prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_43/a_376_368#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_5/a_735_102# prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_35/a_138_385#
+ prbs_generator_syn_23/sky130_fd_sc_hs__sdlclkp_2_1/a_114_424# prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_57/a_132_392#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_71/a_1034_424# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_7/a_1226_296#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_33/a_544_485# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_41/a_696_458#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_71/a_544_485# prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_21/B
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_61/a_1226_296# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_39/a_1034_424#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_17/a_27_74# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_9/a_27_74#
+ prbs_generator_syn_23/sky130_fd_sc_hs__nor2b_1_5/a_27_112# prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_47/a_132_392#
+ prbs_generator_syn_23/sky130_fd_sc_hs__nor2b_1_8/a_278_368# prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_9/B
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_39/a_206_368# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_33/a_27_74#
+ prbs_generator_syn_23/sky130_fd_sc_hs__nand2_1_41/a_117_74# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_69/a_651_503#
+ prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_51/a_293_74# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_21/a_544_485#
+ prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_7/a_138_385# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_32/a_696_458#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_47/a_735_102# prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_33/a_112_119#
+ prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_59/a_222_392# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_17/a_1141_508#
+ prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_55/a_52_123# prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_3/a_293_74#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_7/a_651_503# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_29/a_1226_296#
+ prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_23/a_376_368# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_8/a_544_485#
+ prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_47/B prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_47/a_1178_124#
+ prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_15/a_138_385# prbs_generator_syn_23/sky130_fd_sc_hs__sdlclkp_2_1/a_1195_374#
+ prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_53/a_138_385# prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_37/a_132_392#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_29/a_206_368# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_39/a_437_503#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_59/a_651_503# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_37/a_735_102#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_67/a_1141_508# prbs_generator_syn_23/sky130_fd_sc_hs__and2b_2_1/a_27_74#
+ prbs_generator_syn_23/sky130_fd_sc_hs__conb_1_1/a_165_290# prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_55/a_293_74#
+ prbs_generator_syn_23/sky130_fd_sc_hs__nand2_1_45/a_117_74# prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_63/a_112_119#
+ prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_49/a_222_392# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_37/a_1034_424#
+ prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_23/a_293_74# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_15/a_1141_508#
+ prbs_generator_syn_23/sky130_fd_sc_hs__nand2_1_5/a_117_74# prbs_generator_syn_23/m3_13600_13485#
+ prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_5/a_112_119# prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_13/a_376_368#
+ prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_51/a_376_368# prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_7/a_293_74#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_19/a_206_368# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_57/a_206_368#
+ prbs_generator_syn_23/sky130_fd_sc_hs__sdlclkp_2_1/a_318_74# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_29/a_437_503#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_49/a_651_503# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_25/a_27_74#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_5/a_1226_296# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_41/a_544_485#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_27/a_735_102# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_65/a_1141_508#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_65/a_735_102# prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_3/a_230_79#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_35/a_1034_424# prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_13/a_230_79#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_41/a_27_74# prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_3/a_132_392#
+ prbs_generator_syn_23/sky130_fd_sc_hs__nand2_1_49/a_117_74# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_27/a_1226_296#
+ prbs_generator_syn_23/sky130_fd_sc_hs__nand2_1_15/a_117_74# prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_41/a_376_368#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_45/a_1178_124# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_4/a_735_102#
+ prbs_generator_syn_23/sky130_fd_sc_hs__nand2_1_9/a_117_74# prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_33/a_138_385#
+ prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_17/a_132_392# prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_55/a_132_392#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_9/a_1141_508# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_19/a_437_503#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_57/a_437_503# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_4/a_1226_296#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_32/a_544_485# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_17/a_735_102#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_55/a_735_102# prbs_generator_syn_23/m3_13600_2261#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_65/a_27_74# prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_29/a_222_392#
+ prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_43/a_112_119# prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_19/X
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_25/a_1226_296# prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_31/a_376_368#
+ prbs_generator_syn_23/sky130_fd_sc_hs__or2_1_1/a_63_368# prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_17/a_230_79#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_4/a_27_74# prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_61/a_230_79#
+ prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_63/a_138_385# prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_5/a_222_392#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_8/a_1141_508# prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_41/a_293_74#
+ prbs_generator_syn_23/sky130_fd_sc_hs__nand2_1_31/a_117_74# prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_5/a_138_385#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_63/a_1141_508# prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_19/a_222_392#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_13/a_1141_508# prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_3/a_52_123#
+ prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_13/a_52_123# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_43/a_1178_124#
+ prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_61/a_376_368# prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_35/a_132_392#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_67/a_206_368# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_1/a_1226_296#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_69/a_696_458# prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_31/a_230_79#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_35/a_735_102# prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_23/a_112_119#
+ prbs_generator_syn_23/sky130_fd_sc_hs__nand2_1_35/a_117_74# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_59/a_27_74#
+ prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_13/a_293_74# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_5/a_206_368#
+ prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_50/a_376_368# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_7/a_696_458#
+ prbs_generator_syn_23/sky130_fd_sc_hs__nor2b_1_7/a_278_368# prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_17/a_52_123#
+ prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_43/a_138_385# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_7/a_1141_508#
+ prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_61/a_52_123# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_67/a_437_503#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_61/a_1141_508# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_25/a_735_102#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_59/a_696_458# prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_13/a_112_119#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_33/a_1034_424# prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_51/a_112_119#
+ prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_35/a_230_79# prbs_generator_syn_23/m3_13600_4091#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_23/a_1226_296# prbs_generator_syn_23/sky130_fd_sc_hs__nand2_1_39/a_117_74#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_29/a_27_74# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_5/a_437_503#
+ prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_17/a_293_74# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_41/a_1178_124#
+ prbs_generator_syn_23/sky130_fd_sc_hs__or2_1_1/a_152_368# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_59/a_1178_124#
+ prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_61/a_293_74# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_47/a_206_368#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_39/a_651_503# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_49/a_696_458#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_15/a_735_102# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_32/a_1034_424#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_73/a_1226_296# prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_27/a_222_392#
+ prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_41/a_112_119# prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_31/a_52_123#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_49/a_1034_424# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_29/a_1141_508#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_21/a_1226_296# prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_39/a_230_79#
+ prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_23/a_138_385# prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_51/a_230_79#
+ prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_45/a_132_392# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_37/a_206_368#
+ prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_65/a_293_74# prbs_generator_syn_23/sky130_fd_sc_hs__nand2_1_53/a_117_74#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_47/a_437_503# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_29/a_651_503#
+ prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_31/a_293_74# prbs_generator_syn_23/sky130_fd_sc_hs__nand2_1_21/a_117_74#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_69/a_544_485# prbs_generator_syn_23/sky130_fd_sc_hs__clkbuf_16_1/a_114_74#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_45/a_735_102# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_13/a_27_74#
+ prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_31/a_112_119# prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_57/a_222_392#
+ prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_35/a_52_123# prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_21/a_376_368#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_7/a_544_485# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_57/a_1178_124#
+ prbs_generator_syn_23/m3_13600_6043# prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_13/a_138_385#
+ prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_51/a_138_385# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_5/a_1141_508#
+ prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_3/a_376_368# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_27/a_206_368#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_65/a_206_368# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_37/a_437_503#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_19/a_651_503# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_57/a_651_503#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_59/a_544_485# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_71/a_1226_296#
+ prbs_generator_syn_23/sky130_fd_sc_hs__nand2_1_25/a_117_74# prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_61/a_112_119#
+ prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_47/a_222_392# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_27/a_1141_508#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_53/a_27_74# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_4/a_206_368#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_39/a_1226_296# prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_11/a_376_368#
+ prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_39/a_52_123# prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_41/a_138_385#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_4/a_1141_508# prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_25/a_132_392#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_17/a_206_368# prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_41/A
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_55/a_206_368# prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_51/a_52_123#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_27/a_437_503# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_65/a_437_503#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_49/a_544_485# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_63/a_735_102#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_47/a_1034_424# prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_50/a_112_119#
+ prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_37/a_222_392# prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_59/a_230_79#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_25/a_1141_508# prbs_generator_syn_23/sky130_fd_sc_hs__nor2b_1_4/a_27_112#
+ prbs_generator_syn_23/sky130_fd_sc_hs__sdlclkp_2_1/a_685_81# prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_1/a_132_392#
+ prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_39/a_293_74# prbs_generator_syn_23/sky130_fd_sc_hs__nand2_1_29/a_117_74#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_4/a_437_503# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_55/a_1178_124#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_21/a_27_74# prbs_generator_syn_23/m3_13600_12875#
+ prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_50/a_293_74# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_1/a_735_102#
+ prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_31/a_138_385# prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_15/a_132_392#
+ prbs_generator_syn_23/sky130_fd_sc_hs__nand2_1_1/a_117_74# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_17/a_437_503#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_55/a_437_503# prbs_generator_syn
Xsky130_fd_sc_hs__conb_1_2 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__conb_1_3/LO sky130_fd_sc_hs__conb_1_3/HI
+ sky130_fd_sc_hs__conb_1_3/a_165_290# sky130_fd_sc_hs__conb_1_3/a_21_290# sky130_fd_sc_hs__conb_1
Xsky130_fd_sc_hs__buf_2_120 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__buf_2_121/A sky130_fd_sc_hs__buf_2_121/X
+ sky130_fd_sc_hs__buf_2_121/a_21_260# sky130_fd_sc_hs__buf_2
Xsky130_fd_sc_hs__buf_2_131 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__buf_2_131/A sky130_fd_sc_hs__buf_2_131/X
+ sky130_fd_sc_hs__buf_2_131/a_21_260# sky130_fd_sc_hs__buf_2
Xsky130_fd_sc_hs__buf_2_142 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__buf_2_143/A sky130_fd_sc_hs__buf_2_143/X
+ sky130_fd_sc_hs__buf_2_143/a_21_260# sky130_fd_sc_hs__buf_2
Xsky130_fd_sc_hs__buf_2_153 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__buf_2_153/A sky130_fd_sc_hs__buf_2_153/X
+ sky130_fd_sc_hs__buf_2_153/a_21_260# sky130_fd_sc_hs__buf_2
Xsky130_fd_sc_hs__einvp_2_10 DVSS: DVDD: DVDD: DVSS: dout_n sky130_fd_sc_hs__einvp_2_9/A
+ sky130_fd_sc_hs__dlrtp_1_8/Q sky130_fd_sc_hs__einvp_2_11/a_263_323# sky130_fd_sc_hs__einvp_2_11/a_36_74#
+ sky130_fd_sc_hs__einvp_2_11/a_27_368# sky130_fd_sc_hs__einvp_2
Xsky130_fd_sc_hs__einvp_2_21 DVSS: DVDD: DVDD: DVSS: dout_n sky130_fd_sc_hs__buf_8_1/A
+ sky130_fd_sc_hs__dlrtp_1_21/Q sky130_fd_sc_hs__einvp_2_21/a_263_323# sky130_fd_sc_hs__einvp_2_21/a_36_74#
+ sky130_fd_sc_hs__einvp_2_21/a_27_368# sky130_fd_sc_hs__einvp_2
Xsky130_fd_sc_hs__einvp_2_32 DVSS: DVDD: DVDD: DVSS: dout_n sky130_fd_sc_hs__buf_8_1/A
+ sky130_fd_sc_hs__buf_2_125/X sky130_fd_sc_hs__einvp_2_33/a_263_323# sky130_fd_sc_hs__einvp_2_33/a_36_74#
+ sky130_fd_sc_hs__einvp_2_33/a_27_368# sky130_fd_sc_hs__einvp_2
Xsky130_fd_sc_hs__einvp_2_43 DVSS: DVDD: DVDD: DVSS: dout_n sky130_fd_sc_hs__buf_8_1/X
+ sky130_fd_sc_hs__dlrtp_1_31/Q sky130_fd_sc_hs__einvp_2_43/a_263_323# sky130_fd_sc_hs__einvp_2_43/a_36_74#
+ sky130_fd_sc_hs__einvp_2_43/a_27_368# sky130_fd_sc_hs__einvp_2
Xsky130_fd_sc_hs__einvp_2_54 DVSS: DVDD: DVDD: DVSS: dout_p sky130_fd_sc_hs__inv_4_9/Y
+ sky130_fd_sc_hs__dlrtp_1_39/Q sky130_fd_sc_hs__einvp_2_55/a_263_323# sky130_fd_sc_hs__einvp_2_55/a_36_74#
+ sky130_fd_sc_hs__einvp_2_55/a_27_368# sky130_fd_sc_hs__einvp_2
Xsky130_fd_sc_hs__einvp_2_65 DVSS: DVDD: DVDD: DVSS: dout_p sky130_fd_sc_hs__einvp_2_65/A
+ sky130_fd_sc_hs__dlrtp_1_53/Q sky130_fd_sc_hs__einvp_2_65/a_263_323# sky130_fd_sc_hs__einvp_2_65/a_36_74#
+ sky130_fd_sc_hs__einvp_2_65/a_27_368# sky130_fd_sc_hs__einvp_2
Xsky130_fd_sc_hs__einvp_2_76 DVSS: DVDD: DVDD: DVSS: dout_p sky130_fd_sc_hs__einvp_2_97/A
+ sky130_fd_sc_hs__dlrtp_1_65/Q sky130_fd_sc_hs__einvp_2_77/a_263_323# sky130_fd_sc_hs__einvp_2_77/a_36_74#
+ sky130_fd_sc_hs__einvp_2_77/a_27_368# sky130_fd_sc_hs__einvp_2
Xsky130_fd_sc_hs__einvp_2_87 DVSS: DVDD: DVDD: DVSS: dout_p sky130_fd_sc_hs__einvp_2_97/A
+ sky130_fd_sc_hs__dlrtp_1_63/Q sky130_fd_sc_hs__einvp_2_87/a_263_323# sky130_fd_sc_hs__einvp_2_87/a_36_74#
+ sky130_fd_sc_hs__einvp_2_87/a_27_368# sky130_fd_sc_hs__einvp_2
Xsky130_fd_sc_hs__einvp_2_98 DVSS: DVDD: DVDD: DVSS: dout_p sky130_fd_sc_hs__einvp_2_99/A
+ sky130_fd_sc_hs__dlrtp_1_81/Q sky130_fd_sc_hs__einvp_2_99/a_263_323# sky130_fd_sc_hs__einvp_2_99/a_36_74#
+ sky130_fd_sc_hs__einvp_2_99/a_27_368# sky130_fd_sc_hs__einvp_2
Xsky130_fd_sc_hs__or2b_2_2 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__or2b_2_3/X sky130_fd_sc_hs__or2b_2_1/A
+ sky130_fd_sc_hs__or2b_2_3/A sky130_fd_sc_hs__or2b_2_3/a_470_368# sky130_fd_sc_hs__or2b_2_3/a_27_368#
+ sky130_fd_sc_hs__or2b_2_3/a_187_48# sky130_fd_sc_hs__or2b_2
Xsky130_fd_sc_hs__conb_1_20 DVSS: DVDD: DVDD: DVSS: prbs_generator_syn_9/eqn[2] prbs_generator_syn_9/eqn[1]
+ sky130_fd_sc_hs__conb_1_21/a_165_290# sky130_fd_sc_hs__conb_1_21/a_21_290# sky130_fd_sc_hs__conb_1
Xsky130_fd_sc_hs__conb_1_31 DVSS: DVDD: DVDD: DVSS: prbs_generator_syn_5/eqn[23] prbs_generator_syn_5/eqn[20]
+ sky130_fd_sc_hs__conb_1_31/a_165_290# sky130_fd_sc_hs__conb_1_31/a_21_290# sky130_fd_sc_hs__conb_1
Xsky130_fd_sc_hs__conb_1_42 DVSS: DVDD: DVDD: DVSS: prbs_generator_syn_5/eqn[5] prbs_generator_syn_5/eqn[1]
+ sky130_fd_sc_hs__conb_1_43/a_165_290# sky130_fd_sc_hs__conb_1_43/a_21_290# sky130_fd_sc_hs__conb_1
Xsky130_fd_sc_hs__conb_1_53 DVSS: DVDD: DVDD: DVSS: prbs_generator_syn_7/eqn[21] prbs_generator_syn_7/eqn[20]
+ sky130_fd_sc_hs__conb_1_53/a_165_290# sky130_fd_sc_hs__conb_1_53/a_21_290# sky130_fd_sc_hs__conb_1
Xsky130_fd_sc_hs__conb_1_64 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__conb_1_65/LO
+ sky130_fd_sc_hs__conb_1_65/HI sky130_fd_sc_hs__conb_1_65/a_165_290# sky130_fd_sc_hs__conb_1_65/a_21_290#
+ sky130_fd_sc_hs__conb_1
Xsky130_fd_sc_hs__conb_1_75 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__conb_1_75/LO
+ sky130_fd_sc_hs__conb_1_75/HI sky130_fd_sc_hs__conb_1_75/a_165_290# sky130_fd_sc_hs__conb_1_75/a_21_290#
+ sky130_fd_sc_hs__conb_1
Xsky130_fd_sc_hs__conb_1_86 DVSS: DVDD: DVDD: DVSS: prbs_generator_syn_11/eqn[2] prbs_generator_syn_11/eqn[1]
+ sky130_fd_sc_hs__conb_1_87/a_165_290# sky130_fd_sc_hs__conb_1_87/a_21_290# sky130_fd_sc_hs__conb_1
Xsky130_fd_sc_hs__conb_1_97 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__conb_1_97/LO
+ sky130_fd_sc_hs__conb_1_97/HI sky130_fd_sc_hs__conb_1_97/a_165_290# sky130_fd_sc_hs__conb_1_97/a_21_290#
+ sky130_fd_sc_hs__conb_1
Xsky130_fd_sc_hs__inv_4_60 DVSS: DVDD: DVDD: DVSS: hr_16t4_mux_top_3/din[14] prbs_generator_syn_17/out
+ sky130_fd_sc_hs__inv_4
Xsky130_fd_sc_hs__inv_4_71 DVSS: DVDD: DVDD: DVSS: osc_core_1/pi5_r[0] osc_core_1/pi5_l[0]
+ sky130_fd_sc_hs__inv_4
Xsky130_fd_sc_hs__inv_4_82 DVSS: DVDD: DVDD: DVSS: hr_16t4_mux_top_3/din[6] hr_16t4_mux_top_1/din[6]
+ sky130_fd_sc_hs__inv_4
Xsky130_fd_sc_hs__dlrtp_1_109 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__buf_2_115/A
+ sky130_fd_sc_hs__dlrtp_1_9/GATE sky130_fd_sc_hs__conb_1_133/HI sky130_fd_sc_hs__inv_4_23/A
+ sky130_fd_sc_hs__dlrtp_1_109/a_216_424# sky130_fd_sc_hs__dlrtp_1_109/a_759_508#
+ sky130_fd_sc_hs__dlrtp_1_109/a_565_74# sky130_fd_sc_hs__dlrtp_1_109/a_27_424# sky130_fd_sc_hs__dlrtp_1_109/a_1045_74#
+ sky130_fd_sc_hs__dlrtp_1_109/a_643_74# sky130_fd_sc_hs__dlrtp_1_109/a_817_48# sky130_fd_sc_hs__dlrtp_1_109/a_568_392#
+ sky130_fd_sc_hs__dlrtp_1_109/a_363_74# sky130_fd_sc_hs__dlrtp_1_109/a_769_74# sky130_fd_sc_hs__dlrtp_1
Xsky130_fd_sc_hs__dlrtp_1_11 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__dlrtp_1_9/Q
+ sky130_fd_sc_hs__dlrtp_1_9/GATE sky130_fd_sc_hs__conb_1_117/HI sky130_fd_sc_hs__dlrtp_1_9/D
+ sky130_fd_sc_hs__dlrtp_1_9/a_216_424# sky130_fd_sc_hs__dlrtp_1_9/a_759_508# sky130_fd_sc_hs__dlrtp_1_9/a_565_74#
+ sky130_fd_sc_hs__dlrtp_1_9/a_27_424# sky130_fd_sc_hs__dlrtp_1_9/a_1045_74# sky130_fd_sc_hs__dlrtp_1_9/a_643_74#
+ sky130_fd_sc_hs__dlrtp_1_9/a_817_48# sky130_fd_sc_hs__dlrtp_1_9/a_568_392# sky130_fd_sc_hs__dlrtp_1_9/a_363_74#
+ sky130_fd_sc_hs__dlrtp_1_9/a_769_74# sky130_fd_sc_hs__dlrtp_1
Xsky130_fd_sc_hs__dlrtp_1_22 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__dlrtp_1_24/Q
+ sky130_fd_sc_hs__clkbuf_2_3/X sky130_fd_sc_hs__conb_1_119/HI sky130_fd_sc_hs__dlrtp_1_24/D
+ sky130_fd_sc_hs__dlrtp_1_24/a_216_424# sky130_fd_sc_hs__dlrtp_1_24/a_759_508# sky130_fd_sc_hs__dlrtp_1_24/a_565_74#
+ sky130_fd_sc_hs__dlrtp_1_24/a_27_424# sky130_fd_sc_hs__dlrtp_1_24/a_1045_74# sky130_fd_sc_hs__dlrtp_1_24/a_643_74#
+ sky130_fd_sc_hs__dlrtp_1_24/a_817_48# sky130_fd_sc_hs__dlrtp_1_24/a_568_392# sky130_fd_sc_hs__dlrtp_1_24/a_363_74#
+ sky130_fd_sc_hs__dlrtp_1_24/a_769_74# sky130_fd_sc_hs__dlrtp_1
Xsky130_fd_sc_hs__dlrtp_1_33 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__dlrtp_1_33/Q
+ sky130_fd_sc_hs__clkbuf_2_3/A sky130_fd_sc_hs__conb_1_123/HI sky130_fd_sc_hs__buf_2_15/X
+ sky130_fd_sc_hs__dlrtp_1_33/a_216_424# sky130_fd_sc_hs__dlrtp_1_33/a_759_508# sky130_fd_sc_hs__dlrtp_1_33/a_565_74#
+ sky130_fd_sc_hs__dlrtp_1_33/a_27_424# sky130_fd_sc_hs__dlrtp_1_33/a_1045_74# sky130_fd_sc_hs__dlrtp_1_33/a_643_74#
+ sky130_fd_sc_hs__dlrtp_1_33/a_817_48# sky130_fd_sc_hs__dlrtp_1_33/a_568_392# sky130_fd_sc_hs__dlrtp_1_33/a_363_74#
+ sky130_fd_sc_hs__dlrtp_1_33/a_769_74# sky130_fd_sc_hs__dlrtp_1
Xsky130_fd_sc_hs__dlrtp_1_44 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__dlrtp_1_45/Q
+ sky130_fd_sc_hs__clkbuf_16_53/A sky130_fd_sc_hs__conb_1_123/HI sky130_fd_sc_hs__buf_2_49/X
+ sky130_fd_sc_hs__dlrtp_1_45/a_216_424# sky130_fd_sc_hs__dlrtp_1_45/a_759_508# sky130_fd_sc_hs__dlrtp_1_45/a_565_74#
+ sky130_fd_sc_hs__dlrtp_1_45/a_27_424# sky130_fd_sc_hs__dlrtp_1_45/a_1045_74# sky130_fd_sc_hs__dlrtp_1_45/a_643_74#
+ sky130_fd_sc_hs__dlrtp_1_45/a_817_48# sky130_fd_sc_hs__dlrtp_1_45/a_568_392# sky130_fd_sc_hs__dlrtp_1_45/a_363_74#
+ sky130_fd_sc_hs__dlrtp_1_45/a_769_74# sky130_fd_sc_hs__dlrtp_1
Xsky130_fd_sc_hs__dlrtp_1_55 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__dlrtp_1_55/Q
+ sky130_fd_sc_hs__clkbuf_16_53/A sky130_fd_sc_hs__conb_1_135/HI sky130_fd_sc_hs__dlrtp_1_55/D
+ sky130_fd_sc_hs__dlrtp_1_55/a_216_424# sky130_fd_sc_hs__dlrtp_1_55/a_759_508# sky130_fd_sc_hs__dlrtp_1_55/a_565_74#
+ sky130_fd_sc_hs__dlrtp_1_55/a_27_424# sky130_fd_sc_hs__dlrtp_1_55/a_1045_74# sky130_fd_sc_hs__dlrtp_1_55/a_643_74#
+ sky130_fd_sc_hs__dlrtp_1_55/a_817_48# sky130_fd_sc_hs__dlrtp_1_55/a_568_392# sky130_fd_sc_hs__dlrtp_1_55/a_363_74#
+ sky130_fd_sc_hs__dlrtp_1_55/a_769_74# sky130_fd_sc_hs__dlrtp_1
Xsky130_fd_sc_hs__dlrtp_1_66 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__dlrtp_1_67/Q
+ sky130_fd_sc_hs__clkbuf_16_53/A sky130_fd_sc_hs__conb_1_129/HI sky130_fd_sc_hs__buf_2_57/X
+ sky130_fd_sc_hs__dlrtp_1_67/a_216_424# sky130_fd_sc_hs__dlrtp_1_67/a_759_508# sky130_fd_sc_hs__dlrtp_1_67/a_565_74#
+ sky130_fd_sc_hs__dlrtp_1_67/a_27_424# sky130_fd_sc_hs__dlrtp_1_67/a_1045_74# sky130_fd_sc_hs__dlrtp_1_67/a_643_74#
+ sky130_fd_sc_hs__dlrtp_1_67/a_817_48# sky130_fd_sc_hs__dlrtp_1_67/a_568_392# sky130_fd_sc_hs__dlrtp_1_67/a_363_74#
+ sky130_fd_sc_hs__dlrtp_1_67/a_769_74# sky130_fd_sc_hs__dlrtp_1
Xsky130_fd_sc_hs__dlrtp_1_77 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__dlrtp_1_77/Q
+ sky130_fd_sc_hs__clkbuf_16_53/A sky130_fd_sc_hs__conb_1_129/HI sky130_fd_sc_hs__inv_4_15/A
+ sky130_fd_sc_hs__dlrtp_1_77/a_216_424# sky130_fd_sc_hs__dlrtp_1_77/a_759_508# sky130_fd_sc_hs__dlrtp_1_77/a_565_74#
+ sky130_fd_sc_hs__dlrtp_1_77/a_27_424# sky130_fd_sc_hs__dlrtp_1_77/a_1045_74# sky130_fd_sc_hs__dlrtp_1_77/a_643_74#
+ sky130_fd_sc_hs__dlrtp_1_77/a_817_48# sky130_fd_sc_hs__dlrtp_1_77/a_568_392# sky130_fd_sc_hs__dlrtp_1_77/a_363_74#
+ sky130_fd_sc_hs__dlrtp_1_77/a_769_74# sky130_fd_sc_hs__dlrtp_1
Xsky130_fd_sc_hs__dlrtp_1_88 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__buf_2_71/A sky130_fd_sc_hs__clkbuf_16_53/A
+ sky130_fd_sc_hs__conb_1_137/HI sky130_fd_sc_hs__dlrtp_1_89/D sky130_fd_sc_hs__dlrtp_1_89/a_216_424#
+ sky130_fd_sc_hs__dlrtp_1_89/a_759_508# sky130_fd_sc_hs__dlrtp_1_89/a_565_74# sky130_fd_sc_hs__dlrtp_1_89/a_27_424#
+ sky130_fd_sc_hs__dlrtp_1_89/a_1045_74# sky130_fd_sc_hs__dlrtp_1_89/a_643_74# sky130_fd_sc_hs__dlrtp_1_89/a_817_48#
+ sky130_fd_sc_hs__dlrtp_1_89/a_568_392# sky130_fd_sc_hs__dlrtp_1_89/a_363_74# sky130_fd_sc_hs__dlrtp_1_89/a_769_74#
+ sky130_fd_sc_hs__dlrtp_1
Xsky130_fd_sc_hs__dlrtp_1_99 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__buf_2_99/A sky130_fd_sc_hs__dlrtp_1_9/GATE
+ sky130_fd_sc_hs__conb_1_131/HI sky130_fd_sc_hs__dlrtp_1_99/D sky130_fd_sc_hs__dlrtp_1_99/a_216_424#
+ sky130_fd_sc_hs__dlrtp_1_99/a_759_508# sky130_fd_sc_hs__dlrtp_1_99/a_565_74# sky130_fd_sc_hs__dlrtp_1_99/a_27_424#
+ sky130_fd_sc_hs__dlrtp_1_99/a_1045_74# sky130_fd_sc_hs__dlrtp_1_99/a_643_74# sky130_fd_sc_hs__dlrtp_1_99/a_817_48#
+ sky130_fd_sc_hs__dlrtp_1_99/a_568_392# sky130_fd_sc_hs__dlrtp_1_99/a_363_74# sky130_fd_sc_hs__dlrtp_1_99/a_769_74#
+ sky130_fd_sc_hs__dlrtp_1
Xsky130_fd_sc_hs__einvp_2_4 DVSS: DVDD: DVDD: DVSS: dout_n sky130_fd_sc_hs__buf_8_1/A
+ sky130_fd_sc_hs__dlrtp_1_7/Q sky130_fd_sc_hs__einvp_2_5/a_263_323# sky130_fd_sc_hs__einvp_2_5/a_36_74#
+ sky130_fd_sc_hs__einvp_2_5/a_27_368# sky130_fd_sc_hs__einvp_2
Xsky130_fd_sc_hs__clkbuf_2_7 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__clkbuf_2_7/X
+ sky130_fd_sc_hs__o21ai_2_5/Y sky130_fd_sc_hs__clkbuf_2_7/a_43_192# sky130_fd_sc_hs__clkbuf_2
Xsky130_fd_sc_hs__clkbuf_2_18 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__dlrtp_1_65/D
+ sky130_fd_sc_hs__o21ai_2_15/Y sky130_fd_sc_hs__clkbuf_2_19/a_43_192# sky130_fd_sc_hs__clkbuf_2
Xsky130_fd_sc_hs__clkbuf_2_29 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__o21ai_2_23/A2
+ sky130_fd_sc_hs__or2b_4_5/A sky130_fd_sc_hs__clkbuf_2_29/a_43_192# sky130_fd_sc_hs__clkbuf_2
Xsky130_fd_sc_hs__buf_2_9 DVSS: DVDD: DVDD: DVSS: manual_control_osc[11] sky130_fd_sc_hs__buf_2_9/X
+ sky130_fd_sc_hs__buf_2_9/a_21_260# sky130_fd_sc_hs__buf_2
Xsky130_fd_sc_hs__buf_2_14 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__buf_2_15/A sky130_fd_sc_hs__buf_2_15/X
+ sky130_fd_sc_hs__buf_2_15/a_21_260# sky130_fd_sc_hs__buf_2
Xsky130_fd_sc_hs__buf_2_25 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__buf_2_25/A sky130_fd_sc_hs__buf_2_25/X
+ sky130_fd_sc_hs__buf_2_25/a_21_260# sky130_fd_sc_hs__buf_2
Xsky130_fd_sc_hs__buf_2_36 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__buf_2_37/A sky130_fd_sc_hs__buf_2_37/X
+ sky130_fd_sc_hs__buf_2_37/a_21_260# sky130_fd_sc_hs__buf_2
Xsky130_fd_sc_hs__buf_2_47 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__buf_2_47/A sky130_fd_sc_hs__buf_2_47/X
+ sky130_fd_sc_hs__buf_2_47/a_21_260# sky130_fd_sc_hs__buf_2
Xsky130_fd_sc_hs__buf_2_58 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__buf_2_59/A sky130_fd_sc_hs__buf_2_59/X
+ sky130_fd_sc_hs__buf_2_59/a_21_260# sky130_fd_sc_hs__buf_2
Xsky130_fd_sc_hs__buf_2_69 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__buf_2_69/A sky130_fd_sc_hs__buf_2_69/X
+ sky130_fd_sc_hs__buf_2_69/a_21_260# sky130_fd_sc_hs__buf_2
Xsky130_fd_sc_hs__o21bai_2_16 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__o21bai_2_5/A1
+ sky130_fd_sc_hs__nand2_2_11/B sky130_fd_sc_hs__dlrtp_1_157/D sky130_fd_sc_hs__buf_2_69/A
+ sky130_fd_sc_hs__o21bai_2_17/a_27_74# sky130_fd_sc_hs__o21bai_2_17/a_225_74# sky130_fd_sc_hs__o21bai_2_17/a_507_368#
+ sky130_fd_sc_hs__o21bai_2
Xsky130_fd_sc_hs__o21bai_2_27 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__or2b_2_3/A
+ sky130_fd_sc_hs__clkbuf_4_81/X sky130_fd_sc_hs__dlrtp_1_99/D sky130_fd_sc_hs__buf_2_105/A
+ sky130_fd_sc_hs__o21bai_2_27/a_27_74# sky130_fd_sc_hs__o21bai_2_27/a_225_74# sky130_fd_sc_hs__o21bai_2_27/a_507_368#
+ sky130_fd_sc_hs__o21bai_2
Xsky130_fd_sc_hs__o21bai_2_38 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__o21ai_4_1/A1
+ sky130_fd_sc_hs__clkinv_4_5/Y sky130_fd_sc_hs__dlrtp_1_19/D sky130_fd_sc_hs__buf_2_113/A
+ sky130_fd_sc_hs__o21bai_2_39/a_27_74# sky130_fd_sc_hs__o21bai_2_39/a_225_74# sky130_fd_sc_hs__o21bai_2_39/a_507_368#
+ sky130_fd_sc_hs__o21bai_2
Xsky130_fd_sc_hs__o21bai_2_49 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__nand2_8_1/Y
+ sky130_fd_sc_hs__nand2_2_21/B sky130_fd_sc_hs__dlrtp_1_121/D sky130_fd_sc_hs__o21bai_2_49/Y
+ sky130_fd_sc_hs__o21bai_2_49/a_27_74# sky130_fd_sc_hs__o21bai_2_49/a_225_74# sky130_fd_sc_hs__o21bai_2_49/a_507_368#
+ sky130_fd_sc_hs__o21bai_2
Xsky130_fd_sc_hs__o21bai_4_5 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__buf_2_143/A
+ sky130_fd_sc_hs__nand2_2_5/B sky130_fd_sc_hs__o21bai_4_7/A1 sky130_fd_sc_hs__buf_2_153/X
+ sky130_fd_sc_hs__o21bai_4_5/a_28_368# sky130_fd_sc_hs__o21bai_4_5/a_27_74# sky130_fd_sc_hs__o21bai_4_5/a_828_48#
+ sky130_fd_sc_hs__o21bai_4
Xsky130_fd_sc_hs__conb_1_203 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__conb_1_203/LO
+ sky130_fd_sc_hs__conb_1_203/HI sky130_fd_sc_hs__conb_1_203/a_165_290# sky130_fd_sc_hs__conb_1_203/a_21_290#
+ sky130_fd_sc_hs__conb_1
Xsky130_fd_sc_hs__conb_1_214 DVSS: DVDD: DVDD: DVSS: prbs_generator_syn_25/eqn[9]
+ sky130_fd_sc_hs__conb_1_215/HI sky130_fd_sc_hs__conb_1_215/a_165_290# sky130_fd_sc_hs__conb_1_215/a_21_290#
+ sky130_fd_sc_hs__conb_1
Xsky130_fd_sc_hs__conb_1_225 DVSS: DVDD: DVDD: DVSS: prbs_generator_syn_25/eqn[8]
+ prbs_generator_syn_25/eqn[1] sky130_fd_sc_hs__conb_1_225/a_165_290# sky130_fd_sc_hs__conb_1_225/a_21_290#
+ sky130_fd_sc_hs__conb_1
Xsky130_fd_sc_hs__conb_1_236 DVSS: DVDD: DVDD: DVSS: prbs_generator_syn_27/eqn[22]
+ prbs_generator_syn_27/eqn[20] sky130_fd_sc_hs__conb_1_237/a_165_290# sky130_fd_sc_hs__conb_1_237/a_21_290#
+ sky130_fd_sc_hs__conb_1
Xsky130_fd_sc_hs__conb_1_247 DVSS: DVDD: DVDD: DVSS: prbs_generator_syn_31/eqn[28]
+ sky130_fd_sc_hs__conb_1_247/HI sky130_fd_sc_hs__conb_1_247/a_165_290# sky130_fd_sc_hs__conb_1_247/a_21_290#
+ sky130_fd_sc_hs__conb_1
Xsky130_fd_sc_hs__conb_1_258 DVSS: DVDD: DVDD: DVSS: prbs_generator_syn_31/eqn[30]
+ sky130_fd_sc_hs__conb_1_259/HI sky130_fd_sc_hs__conb_1_259/a_165_290# sky130_fd_sc_hs__conb_1_259/a_21_290#
+ sky130_fd_sc_hs__conb_1
Xsky130_fd_sc_hs__conb_1_269 DVSS: DVDD: DVDD: DVSS: prbs_generator_syn_31/eqn[2]
+ prbs_generator_syn_31/eqn[1] sky130_fd_sc_hs__conb_1_269/a_165_290# sky130_fd_sc_hs__conb_1_269/a_21_290#
+ sky130_fd_sc_hs__conb_1
Xsky130_fd_sc_hs__clkbuf_8_17 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__clkbuf_8_17/X
+ sky130_fd_sc_hs__buf_2_9/X sky130_fd_sc_hs__clkbuf_8_17/a_125_368# sky130_fd_sc_hs__clkbuf_8
Xsky130_fd_sc_hs__clkbuf_8_28 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__clkbuf_8_29/X
+ sky130_fd_sc_hs__clkbuf_8_29/A sky130_fd_sc_hs__clkbuf_8_29/a_125_368# sky130_fd_sc_hs__clkbuf_8
Xsky130_fd_sc_hs__clkbuf_8_39 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__nand2_2_21/B
+ sky130_fd_sc_hs__or2b_2_3/X sky130_fd_sc_hs__clkbuf_8_39/a_125_368# sky130_fd_sc_hs__clkbuf_8
Xsky130_fd_sc_hs__o21bai_2_2 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__nand2_2_5/B
+ sky130_fd_sc_hs__o21bai_2_3/A2 sky130_fd_sc_hs__buf_2_55/X sky130_fd_sc_hs__o21bai_2_3/Y
+ sky130_fd_sc_hs__o21bai_2_3/a_27_74# sky130_fd_sc_hs__o21bai_2_3/a_225_74# sky130_fd_sc_hs__o21bai_2_3/a_507_368#
+ sky130_fd_sc_hs__o21bai_2
Xsky130_fd_sc_hs__o21ai_2_40 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__inv_4_23/Y sky130_fd_sc_hs__nand2_2_15/B
+ sky130_fd_sc_hs__clkinv_4_7/Y sky130_fd_sc_hs__o21ai_2_41/Y sky130_fd_sc_hs__o21ai_2_41/a_116_368#
+ sky130_fd_sc_hs__o21ai_2_41/a_27_74# sky130_fd_sc_hs__o21ai_2
Xsky130_fd_sc_hs__o21ai_2_51 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__inv_4_25/Y sky130_fd_sc_hs__or2b_4_1/A
+ sky130_fd_sc_hs__o21ai_2_51/A1 sky130_fd_sc_hs__o21ai_2_51/Y sky130_fd_sc_hs__o21ai_2_51/a_116_368#
+ sky130_fd_sc_hs__o21ai_2_51/a_27_74# sky130_fd_sc_hs__o21ai_2
Xsky130_fd_sc_hs__clkinv_4_10 DVSS: DVDD: DVDD: DVSS: osc_core_1/pi2_r[3] osc_core_1/pi2_l[3]
+ sky130_fd_sc_hs__clkinv_4
Xprbs_generator_syn_12 prbs_generator_syn_19/clk prbs_generator_syn_13/rst prbs_generator_syn_13/cke
+ sky130_fd_sc_hs__conb_1_109/LO sky130_fd_sc_hs__conb_1_109/LO sky130_fd_sc_hs__conb_1_109/LO
+ sky130_fd_sc_hs__conb_1_109/LO sky130_fd_sc_hs__conb_1_109/LO sky130_fd_sc_hs__conb_1_109/LO
+ sky130_fd_sc_hs__conb_1_109/HI sky130_fd_sc_hs__conb_1_109/HI sky130_fd_sc_hs__conb_1_109/HI
+ sky130_fd_sc_hs__conb_1_109/HI sky130_fd_sc_hs__conb_1_109/HI prbs_generator_syn_13/cke
+ sky130_fd_sc_hs__conb_1_111/HI sky130_fd_sc_hs__conb_1_111/HI sky130_fd_sc_hs__conb_1_111/HI
+ sky130_fd_sc_hs__conb_1_111/HI prbs_generator_syn_15/eqn[13] sky130_fd_sc_hs__conb_1_111/HI
+ prbs_generator_syn_13/eqn[2] prbs_generator_syn_13/eqn[1] prbs_generator_syn_13/eqn[2]
+ prbs_generator_syn_13/eqn[1] prbs_generator_syn_13/eqn[2] prbs_generator_syn_13/eqn[1]
+ sky130_fd_sc_hs__conb_1_115/LO sky130_fd_sc_hs__conb_1_115/HI sky130_fd_sc_hs__conb_1_115/LO
+ sky130_fd_sc_hs__conb_1_115/LO sky130_fd_sc_hs__conb_1_115/HI sky130_fd_sc_hs__conb_1_115/HI
+ sky130_fd_sc_hs__conb_1_115/LO sky130_fd_sc_hs__conb_1_115/LO prbs_generator_syn_13/eqn[31]
+ prbs_generator_syn_13/eqn[30] prbs_generator_syn_13/eqn[30] prbs_generator_syn_13/eqn[30]
+ prbs_generator_syn_13/eqn[30] prbs_generator_syn_13/eqn[30] prbs_generator_syn_13/eqn[30]
+ prbs_generator_syn_13/eqn[30] prbs_generator_syn_13/eqn[30] prbs_generator_syn_13/eqn[22]
+ prbs_generator_syn_13/eqn[22] prbs_generator_syn_13/eqn[20] prbs_generator_syn_13/eqn[22]
+ prbs_generator_syn_13/eqn[22] prbs_generator_syn_13/eqn[22] prbs_generator_syn_13/eqn[22]
+ prbs_generator_syn_13/eqn[22] prbs_generator_syn_13/eqn[22] sky130_fd_sc_hs__conb_1_97/LO
+ sky130_fd_sc_hs__conb_1_97/LO sky130_fd_sc_hs__conb_1_97/LO prbs_generator_syn_13/eqn[9]
+ prbs_generator_syn_13/eqn[9] prbs_generator_syn_13/eqn[9] prbs_generator_syn_13/eqn[9]
+ prbs_generator_syn_13/eqn[9] prbs_generator_syn_13/eqn[9] prbs_generator_syn_13/eqn[9]
+ prbs_generator_syn_13/eqn[9] prbs_generator_syn_13/eqn[2] prbs_generator_syn_13/eqn[1]
+ prbs_generator_syn_13/eqn[2] prbs_generator_syn_19/inj_err prbs_generator_syn_13/eqn[31]
+ prbs_generator_syn_13/eqn[31] hr_16t4_mux_top_1/din[5] DVSS: DVDD: prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_1/a_293_74#
+ prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_15/X prbs_generator_syn_13/sky130_fd_sc_hs__nand2_1_35/B
+ prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_51/Y prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_9/A
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_9/CLK prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_47/a_27_74#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_37/a_1226_296# prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_3/B
+ prbs_generator_syn_13/sky130_fd_sc_hs__nor2b_1_7/a_27_112# prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_29/B
+ prbs_generator_syn_13/sky130_fd_sc_hs__sdlclkp_2_1/a_580_74# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_1/a_1141_508#
+ prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_5/Y prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_41/a_230_79#
+ prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_61/a_138_385# prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_43/a_132_392#
+ prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_3/a_222_392# prbs_generator_syn_13/sky130_fd_sc_hs__nor2b_1_9/a_27_112#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_61/a_27_74# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_35/a_206_368#
+ prbs_generator_syn_13/sky130_fd_sc_hs__nand2_2_3/Y prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_25/B
+ prbs_generator_syn_13/sky130_fd_sc_hs__nand2_1_11/a_117_74# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_67/a_651_503#
+ prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_45/X prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_39/a_696_458#
+ prbs_generator_syn_13/sky130_fd_sc_hs__sdlclkp_2_1/a_1198_74# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_45/a_1034_424#
+ prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_17/a_222_392# prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_55/a_222_392#
+ prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_53/Y prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_35/A
+ prbs_generator_syn_13/m3_13600_1651# prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_59/a_52_123#
+ prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_5/a_293_74# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_35/a_1226_296#
+ prbs_generator_syn_13/sky130_fd_sc_hs__nand2_1_51/B prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_5/a_651_503#
+ prbs_generator_syn_13/sky130_fd_sc_hs__nand2_1_21/B prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_8/a_27_74#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_15/a_27_74# prbs_generator_syn_13/sky130_fd_sc_hs__and2b_2_1/X
+ prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_13/X prbs_generator_syn_13/sky130_fd_sc_hs__nand2_2_3/a_27_74#
+ prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_50/a_138_385# prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_33/a_132_392#
+ prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_1/a_376_368# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_25/a_206_368#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_35/a_437_503# prbs_generator_syn_13/sky130_fd_sc_hs__sdlclkp_2_1/a_708_451#
+ prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_45/a_230_79# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_29/a_696_458#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_32/a_27_74# prbs_generator_syn_13/sky130_fd_sc_hs__nor2b_1_4/Y
+ prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_59/a_293_74# prbs_generator_syn_13/sky130_fd_sc_hs__nand2_1_47/a_117_74#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_73/a_735_102# prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_21/a_112_119#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_23/a_1141_508# prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_25/a_293_74#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_7/Q prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_3/a_112_119#
+ prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_35/B prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_51/X
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_53/a_1178_124# prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_23/a_132_392#
+ prbs_generator_syn_13/sky130_fd_sc_hs__nand2_1_3/B prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_15/a_206_368#
+ prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_63/a_132_392# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_55/a_27_74#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_25/a_437_503# prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_41/a_52_123#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_47/a_651_503# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_73/a_1141_508#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_19/a_696_458# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_57/a_696_458#
+ prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_7/X prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_43/a_1034_424#
+ prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_55/A prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_11/a_112_119#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_21/a_1141_508# prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_35/a_222_392#
+ prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_49/a_230_79# prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_67/Y
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_71/a_27_74# prbs_generator_syn_13/sky130_fd_sc_hs__nand2_1_33/B
+ prbs_generator_syn_13/sky130_fd_sc_hs__conb_1_1/LO prbs_generator_syn_13/sky130_fd_sc_hs__nand2_1_19/a_117_74#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_51/a_1178_124# prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_33/X
+ prbs_generator_syn_13/sky130_fd_sc_hs__nand2_1_29/B prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_41/Y
+ prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_53/a_132_392# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_45/a_206_368#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_15/a_437_503# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_37/a_651_503#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_39/a_544_485# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_53/a_735_102#
+ prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_45/a_52_123# prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_1/B
+ prbs_generator_syn_13/sky130_fd_sc_hs__nand2_2_3/B prbs_generator_syn_13/sky130_fd_sc_hs__clkbuf_16_1/A
+ prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_21/X prbs_generator_syn_13/sky130_fd_sc_hs__nand2_1_25/B
+ prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_39/a_376_368# prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_63/X
+ prbs_generator_syn_13/m3_13600_3481# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_69/a_1178_124#
+ prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_21/a_138_385# prbs_generator_syn_13/sky130_fd_sc_hs__nor2b_1_8/Y
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_19/a_1178_124# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_49/a_27_74#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_45/a_437_503# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_27/a_651_503#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_71/a_1141_508# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_65/a_651_503#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_29/a_544_485# prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_3/a_138_385#
+ prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_55/X prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_43/a_735_102#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_41/a_1034_424# prbs_generator_syn_13/sky130_fd_sc_hs__nand2_1_9/B
+ prbs_generator_syn_13/sky130_fd_sc_hs__nor2b_1_9/Y prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_59/a_1034_424#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_39/a_1141_508# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_33/a_1226_296#
+ prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_49/a_52_123# prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_47/Y
+ prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_43/Y prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_4/a_651_503#
+ prbs_generator_syn_13/sky130_fd_sc_hs__nand2_1_49/B prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_19/A
+ prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_11/a_138_385# prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_5/X
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_63/a_206_368# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_17/a_651_503#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_19/a_544_485# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_55/a_651_503#
+ prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_9/Y prbs_generator_syn_13/sky130_fd_sc_hs__nand2_1_17/B
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_57/a_544_485# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_67/a_696_458#
+ prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_35/X prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_19/a_27_74#
+ prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_45/a_222_392# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_32/a_1226_296#
+ prbs_generator_syn_13/sky130_fd_sc_hs__nand2_1_43/B prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_25/A
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_1/a_206_368# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_49/a_1226_296#
+ prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_1/a_112_119# prbs_generator_syn_13/sky130_fd_sc_hs__or2_1_1/X
+ prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_59/a_376_368# prbs_generator_syn_13/sky130_fd_sc_hs__nand2_1_19/B
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_5/a_696_458# prbs_generator_syn_13/sky130_fd_sc_hs__nor2b_1_1/Y
+ prbs_generator_syn_13/sky130_fd_sc_hs__nor2b_1_5/a_278_368# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_17/a_1178_124#
+ prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_39/X prbs_generator_syn_13/m3_13600_5433#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_63/a_437_503# prbs_generator_syn_13/sky130_fd_sc_hs__nand2_2_5/B
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_23/a_735_102# prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_53/A
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_61/a_735_102# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_57/a_1034_424#
+ prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_63/B prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_37/a_1141_508#
+ prbs_generator_syn_13/sky130_fd_sc_hs__nand2_1_47/B prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_29/X
+ prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_65/Y prbs_generator_syn_13/m3_13600_4701#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_1/a_437_503# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_67/a_1178_124#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_9/a_735_102# prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_13/a_132_392#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_15/a_1178_124# prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_15/A
+ prbs_generator_syn_13/sky130_fd_sc_hs__nand2_1_1/B prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_43/B
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_35/a_651_503# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_8/D
+ prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_29/A prbs_generator_syn_13/sky130_fd_sc_hs__nand2_1_7/B
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_13/a_735_102# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_47/a_696_458#
+ prbs_generator_syn_13/sky130_fd_sc_hs__nand2_1_31/B prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_51/a_735_102#
+ prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_59/X prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_35/a_1141_508#
+ prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_25/a_222_392# prbs_generator_syn_13/sky130_fd_sc_hs__sdlclkp_2_1/a_288_48#
+ prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_55/B prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_17/B
+ prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_43/A prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_7/A
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_65/a_1178_124# prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_59/Y
+ prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_41/X prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_21/a_230_79#
+ prbs_generator_syn_13/sky130_fd_sc_hs__nand2_1_57/a_117_74# prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_1/a_222_392#
+ prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_19/B prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_35/a_293_74#
+ prbs_generator_syn_13/sky130_fd_sc_hs__nand2_1_23/a_117_74# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_73/a_206_368#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_25/a_651_503# prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_1/a_138_385#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_37/a_696_458# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_67/a_544_485#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_43/a_27_74# prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_9/X
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_55/a_1034_424# prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_39/a_112_119#
+ prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_15/a_222_392# prbs_generator_syn_13/sky130_fd_sc_hs__conb_1_1/HI
+ prbs_generator_syn_13/sky130_fd_sc_hs__nand2_1_23/B prbs_generator_syn_13/sky130_fd_sc_hs__nand2_1_53/B
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_9/a_1178_124# prbs_generator_syn_13/sky130_fd_sc_hs__nor2b_1_4/A
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_47/a_1226_296# prbs_generator_syn_13/m3_13600_11045#
+ prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_17/X prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_29/a_376_368#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_5/a_544_485# prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_3/X
+ prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_31/a_132_392# prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_61/A
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_15/a_651_503# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_73/a_437_503#
+ prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_25/a_230_79# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_27/a_696_458#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_65/a_696_458# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_33/a_735_102#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_71/a_735_102# prbs_generator_syn_13/m3_13600_7263#
+ prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_43/a_222_392# prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_50/Y
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_8/a_1178_124# prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_53/B
+ prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_19/a_376_368# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_63/a_1178_124#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_4/a_696_458# prbs_generator_syn_13/sky130_fd_sc_hs__nor2b_1_4/a_278_368#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_13/a_1178_124# prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_61/a_132_392#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_53/a_206_368# prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_21/a_52_123#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_45/a_651_503# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_17/a_696_458#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_47/a_544_485# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_55/a_696_458#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_21/a_735_102# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_37/a_27_74#
+ prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_61/B prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_61/X
+ prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_59/a_112_119# prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_31/A
+ prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_33/a_222_392# prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_29/a_230_79#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_45/a_1226_296# prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_9/a_132_392#
+ prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_5/A prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_57/Y
+ prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_31/X prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_51/a_27_74#
+ prbs_generator_syn_13/sky130_fd_sc_hs__nor2b_1_8/a_27_112# prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_47/a_376_368#
+ prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_53/a_293_74# prbs_generator_syn_13/sky130_fd_sc_hs__nand2_1_43/a_117_74#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_8/a_735_102# prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_21/a_293_74#
+ prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_39/a_138_385# prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_63/Y
+ prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_51/a_132_392# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_43/a_206_368#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_53/a_437_503# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_37/a_544_485#
+ prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_57/X prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_53/a_1034_424#
+ prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_25/a_52_123# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_33/a_1141_508#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_63/Q prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_23/a_222_392#
+ prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_63/a_222_392# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_7/a_1178_124#
+ prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_53/X prbs_generator_syn_13/sky130_fd_sc_hs__nand2_2_5/Y
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_61/a_1178_124# prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_1/a_230_79#
+ prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_43/a_230_79# prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_11/a_230_79#
+ prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_41/a_132_392# prbs_generator_syn_13/sky130_fd_sc_hs__nand2_1_13/a_117_74#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_43/a_437_503# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_27/a_544_485#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_63/a_651_503# prbs_generator_syn_13/sky130_fd_sc_hs__nand2_1_7/a_117_74#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_35/a_696_458# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_65/a_544_485#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_51/a_1034_424# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_41/a_735_102#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_32/a_1141_508# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_49/a_1141_508#
+ prbs_generator_syn_13/sky130_fd_sc_hs__nand2_1_55/B prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_53/a_222_392#
+ prbs_generator_syn_13/sky130_fd_sc_hs__sdlclkp_2_1/a_114_112# prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_9/a_293_74#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_43/a_1226_296# prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_29/a_52_123#
+ prbs_generator_syn_13/sky130_fd_sc_hs__nand2_1_37/B prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_1/a_651_503#
+ prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_27/a_376_368# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_4/a_544_485#
+ prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_67/a_376_368# prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_27/X
+ prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_1/X prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_59/a_138_385#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_29/a_1178_124# prbs_generator_syn_13/m3_13600_2871#
+ prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_5/a_230_79# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_23/a_206_368#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_61/a_206_368# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_17/a_544_485#
+ prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_15/a_230_79# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_25/a_696_458#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_55/a_544_485# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_32/a_735_102#
+ prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_29/a_293_74# prbs_generator_syn_13/sky130_fd_sc_hs__nand2_1_17/a_117_74#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_69/a_1034_424# prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_29/a_112_119#
+ prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_37/X prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_31/B
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_19/a_1034_424# prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_33/A
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_9/a_206_368# prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_57/a_376_368#
+ prbs_generator_syn_13/sky130_fd_sc_hs__sdlclkp_2_1/a_706_317# prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_11/B
+ prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_1/a_52_123# prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_39/B
+ prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_21/a_132_392# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_13/a_206_368#
+ prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_43/a_52_123# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_51/a_206_368#
+ prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_47/X prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_23/a_437_503#
+ prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_11/a_52_123# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_61/a_437_503#
+ prbs_generator_syn_13/sky130_fd_sc_hs__nor2b_1_7/Y prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_51/A
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_15/a_696_458# prbs_generator_syn_13/sky130_fd_sc_hs__nor2b_1_5/Y
+ prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_9/a_230_79# prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_25/X
+ prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_19/a_112_119# prbs_generator_syn_13/sky130_fd_sc_hs__nand2_1_45/B
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_5/a_1178_124# prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_19/a_230_79#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_41/a_1226_296# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_59/a_1226_296#
+ prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_63/a_230_79# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_51/Q
+ prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_7/a_132_392# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_9/a_437_503#
+ prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_46/a_376_368# prbs_generator_syn_13/sky130_fd_sc_hs__nand2_1_33/a_117_74#
+ prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_11/a_293_74# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_27/a_1178_124#
+ prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_11/a_132_392# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_13/a_437_503#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_51/a_437_503# prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_5/a_52_123#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_35/a_544_485# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_73/a_651_503#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_45/a_696_458# prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_15/a_52_123#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_47/a_1141_508# prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_47/a_112_119#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_4/a_1178_124# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_17/a_1034_424#
+ prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_23/B prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_37/a_376_368#
+ prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_15/B prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_7/Y
+ prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_29/a_138_385# prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_33/a_230_79#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_25/a_1178_124# prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_47/a_293_74#
+ prbs_generator_syn_13/sky130_fd_sc_hs__nand2_1_37/a_117_74# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_33/a_206_368#
+ prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_15/a_293_74# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_71/a_206_368#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_25/a_544_485# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_67/a_1034_424#
+ prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_13/a_222_392# prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_9/a_52_123#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_15/a_1034_424# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_57/a_1226_296#
+ prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_19/a_52_123# prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_23/X
+ prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_63/a_52_123# prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_19/a_138_385#
+ prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_9/a_376_368# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_21/a_206_368#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_33/a_437_503# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_71/a_437_503#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_53/a_651_503# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_15/a_544_485#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_63/a_696_458# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_65/a_1034_424#
+ prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_19/a_293_74# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_45/a_1141_508#
+ prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_27/a_112_119# prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_67/a_112_119#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_1/a_1178_124# prbs_generator_syn_13/sky130_fd_sc_hs__conb_1_1/a_21_290#
+ prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_63/a_293_74# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_8/a_206_368#
+ prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_17/a_376_368# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_63/a_27_74#
+ prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_21/A prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_55/a_376_368#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_1/a_696_458# prbs_generator_syn_13/sky130_fd_sc_hs__nor2b_1_1/a_278_368#
+ prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_47/a_138_385# prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_33/a_52_123#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_9/a_1034_424# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_21/a_437_503#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_1/a_27_74# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_43/a_651_503#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_1/Q prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_45/a_544_485#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_69/a_735_102# prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_57/a_112_119#
+ prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_31/a_222_392# prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_13/A
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_55/a_1226_296# prbs_generator_syn_13/sky130_fd_sc_hs__nand2_2_5/a_27_74#
+ prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_53/a_230_79# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_8/a_437_503#
+ prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_67/a_293_74# prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_33/a_293_74#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_7/a_735_102# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_23/a_1178_124#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_41/a_206_368# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_8/a_1034_424#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_63/a_1034_424# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_59/a_735_102#
+ prbs_generator_syn_13/sky130_fd_sc_hs__nand2_1_5/B prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_43/a_1141_508#
+ prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_46/a_112_119# prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_61/a_222_392#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_13/a_1034_424# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_73/a_1178_124#
+ prbs_generator_syn_13/sky130_fd_sc_hs__nand2_1_27/B prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_13/B
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_57/a_27_74# prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_57/a_230_79#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_21/a_1178_124# prbs_generator_syn_13/sky130_fd_sc_hs__nor2b_1_1/a_27_112#
+ prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_27/a_138_385# prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_23/a_230_79#
+ prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_67/a_138_385# prbs_generator_syn_13/sky130_fd_sc_hs__nand2_1_41/B
+ prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_9/a_222_392# prbs_generator_syn_13/sky130_fd_sc_hs__nand2_1_27/a_117_74#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_32/a_206_368# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_23/a_651_503#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_41/a_437_503# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_73/a_27_74#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_61/a_651_503# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_63/a_544_485#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_49/a_735_102# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_73/a_696_458#
+ prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_37/a_112_119# prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_51/a_222_392#
+ prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_43/X prbs_generator_syn_13/sky130_fd_sc_hs__nand2_2_1/B
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_9/a_651_503# prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_53/a_52_123#
+ prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_49/X prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_25/a_376_368#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_1/a_544_485# prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_65/a_376_368#
+ prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_57/a_138_385# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_27/a_27_74#
+ prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_39/a_132_392# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_7/a_1034_424#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_13/a_651_503# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_32/a_437_503#
+ prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_27/a_230_79# prbs_generator_syn_13/m3_13600_12265#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_51/a_651_503# prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_59/B
+ prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_47/A prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_61/a_1034_424#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_41/a_1141_508# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_59/a_1141_508#
+ prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_41/a_222_392# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_53/a_1226_296#
+ prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_3/A prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_71/a_1178_124#
+ prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_9/a_112_119# prbs_generator_syn_13/sky130_fd_sc_hs__nand2_1_3/a_117_74#
+ prbs_generator_syn_13/m3_13600_8483# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_39/a_1178_124#
+ prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_57/a_52_123# prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_46/a_138_385#
+ prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_23/a_52_123# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_67/a_27_74#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_53/a_696_458# prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_17/a_112_119#
+ prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_11/A prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_55/a_112_119#
+ prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_1/A prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_51/a_1226_296#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_29/a_1034_424# prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_59/A
+ prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_23/A prbs_generator_syn_13/sky130_fd_sc_hs__nand2_1_39/B
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_5/a_27_74# prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_57/a_293_74#
+ prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_37/a_138_385# prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_59/a_132_392#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_33/a_651_503# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_71/a_651_503#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_43/a_696_458# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_73/a_544_485#
+ prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_27/a_52_123# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_57/a_1141_508#
+ prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_21/a_222_392# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_35/a_27_74#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_69/a_1226_296# prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_37/B
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_19/a_1226_296# prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_35/a_376_368#
+ prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_47/a_230_79# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_37/a_1178_124#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_5/a_1034_424# prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_49/a_132_392#
+ prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_7/a_222_392# prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_27/a_293_74#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_21/a_651_503# prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_9/a_138_385#
+ prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_11/a_222_392# prbs_generator_syn_13/m3_13600_14095#
+ prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_50/A prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_27/a_1034_424#
+ prbs_generator_syn_13/sky130_fd_sc_hs__nand2_1_13/B prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_8/a_651_503#
+ prbs_generator_syn_13/m3_13600_9703# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_35/a_1178_124#
+ prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_17/a_138_385# prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_55/a_138_385#
+ prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_7/a_230_79# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_4/a_1034_424#
+ prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_7/a_376_368# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_69/a_206_368#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_23/a_696_458# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_53/a_544_485#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_39/a_735_102# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_61/a_696_458#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_55/a_1141_508# prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_25/a_112_119#
+ prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_65/a_112_119# prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_43/a_293_74#
+ prbs_generator_syn_13/sky130_fd_sc_hs__nand2_1_57/B prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_25/a_1034_424#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_7/a_206_368# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_17/a_1226_296#
+ prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_15/a_376_368# prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_53/a_376_368#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_9/a_696_458# prbs_generator_syn_13/m3_13600_431#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_45/a_27_74# prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_47/a_52_123#
+ prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_29/a_132_392# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_59/a_206_368#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_69/a_437_503# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_41/a_651_503#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_43/a_544_485# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_13/a_696_458#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_29/a_735_102# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_51/a_696_458#
+ prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_61/Y prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_67/a_1226_296#
+ prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_5/a_132_392# prbs_generator_syn_13/sky130_fd_sc_hs__and2b_2_1/a_198_48#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_7/a_437_503# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_15/a_1226_296#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_69/a_27_74# prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_46/a_293_74#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_1/a_1034_424# prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_19/a_132_392#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_49/a_206_368# prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_7/a_52_123#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_59/a_437_503# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_32/a_651_503#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_7/a_27_74# prbs_generator_syn_13/sky130_fd_sc_hs__nand2_2_1/a_27_74#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_19/a_735_102# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_57/a_735_102#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_65/a_1226_296# prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_37/A
+ prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_33/a_376_368# prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_37/a_230_79#
+ prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_25/a_138_385# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_39/a_27_74#
+ prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_65/a_138_385# prbs_generator_syn_13/sky130_fd_sc_hs__nor2b_1_9/a_278_368#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_49/a_437_503# prbs_generator_syn_13/sky130_fd_sc_hs__and2b_2_1/a_505_74#
+ prbs_generator_syn_13/sky130_fd_sc_hs__nand2_1_51/a_117_74# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_23/a_544_485#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_33/a_696_458# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_61/a_544_485#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_9/a_1226_296# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_53/a_1141_508#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_71/a_696_458# prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_35/a_112_119#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_23/a_1034_424# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_9/a_544_485#
+ prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_63/a_376_368# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_33/a_1178_124#
+ prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_5/a_376_368# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_13/a_544_485#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_73/a_1034_424# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_21/a_696_458#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_51/a_544_485# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_8/a_1226_296#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_51/a_1141_508# prbs_generator_syn_13/sky130_fd_sc_hs__nand2_1_55/a_117_74#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_21/a_1034_424# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_63/a_1226_296#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_23/a_27_74# prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_7/a_112_119#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_13/a_1226_296# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_8/a_696_458#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_32/a_1178_124# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_49/a_1178_124#
+ prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_37/a_52_123# prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_27/a_132_392#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_71/Q prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_67/a_735_102#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_69/a_1141_508# prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_15/a_112_119#
+ prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_53/a_112_119# prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_39/a_222_392#
+ prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_55/a_230_79# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_19/a_1141_508#
+ prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_37/a_293_74# prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_43/a_376_368#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_5/a_735_102# prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_35/a_138_385#
+ prbs_generator_syn_13/sky130_fd_sc_hs__sdlclkp_2_1/a_114_424# prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_57/a_132_392#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_71/a_1034_424# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_7/a_1226_296#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_33/a_544_485# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_41/a_696_458#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_71/a_544_485# prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_21/B
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_61/a_1226_296# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_39/a_1034_424#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_17/a_27_74# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_9/a_27_74#
+ prbs_generator_syn_13/sky130_fd_sc_hs__nor2b_1_5/a_27_112# prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_47/a_132_392#
+ prbs_generator_syn_13/sky130_fd_sc_hs__nor2b_1_8/a_278_368# prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_9/B
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_39/a_206_368# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_33/a_27_74#
+ prbs_generator_syn_13/sky130_fd_sc_hs__nand2_1_41/a_117_74# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_69/a_651_503#
+ prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_51/a_293_74# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_21/a_544_485#
+ prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_7/a_138_385# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_32/a_696_458#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_47/a_735_102# prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_33/a_112_119#
+ prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_59/a_222_392# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_17/a_1141_508#
+ prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_55/a_52_123# prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_3/a_293_74#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_7/a_651_503# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_29/a_1226_296#
+ prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_23/a_376_368# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_8/a_544_485#
+ prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_47/B prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_47/a_1178_124#
+ prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_15/a_138_385# prbs_generator_syn_13/sky130_fd_sc_hs__sdlclkp_2_1/a_1195_374#
+ prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_53/a_138_385# prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_37/a_132_392#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_29/a_206_368# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_39/a_437_503#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_59/a_651_503# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_37/a_735_102#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_67/a_1141_508# prbs_generator_syn_13/sky130_fd_sc_hs__and2b_2_1/a_27_74#
+ prbs_generator_syn_13/sky130_fd_sc_hs__conb_1_1/a_165_290# prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_55/a_293_74#
+ prbs_generator_syn_13/sky130_fd_sc_hs__nand2_1_45/a_117_74# prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_63/a_112_119#
+ prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_49/a_222_392# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_37/a_1034_424#
+ prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_23/a_293_74# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_15/a_1141_508#
+ prbs_generator_syn_13/sky130_fd_sc_hs__nand2_1_5/a_117_74# prbs_generator_syn_13/m3_13600_13485#
+ prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_5/a_112_119# prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_13/a_376_368#
+ prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_51/a_376_368# prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_7/a_293_74#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_19/a_206_368# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_57/a_206_368#
+ prbs_generator_syn_13/sky130_fd_sc_hs__sdlclkp_2_1/a_318_74# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_29/a_437_503#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_49/a_651_503# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_25/a_27_74#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_5/a_1226_296# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_41/a_544_485#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_27/a_735_102# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_65/a_1141_508#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_65/a_735_102# prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_3/a_230_79#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_35/a_1034_424# prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_13/a_230_79#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_41/a_27_74# prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_3/a_132_392#
+ prbs_generator_syn_13/sky130_fd_sc_hs__nand2_1_49/a_117_74# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_27/a_1226_296#
+ prbs_generator_syn_13/sky130_fd_sc_hs__nand2_1_15/a_117_74# prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_41/a_376_368#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_45/a_1178_124# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_4/a_735_102#
+ prbs_generator_syn_13/sky130_fd_sc_hs__nand2_1_9/a_117_74# prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_33/a_138_385#
+ prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_17/a_132_392# prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_55/a_132_392#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_9/a_1141_508# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_19/a_437_503#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_57/a_437_503# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_4/a_1226_296#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_32/a_544_485# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_17/a_735_102#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_55/a_735_102# prbs_generator_syn_13/m3_13600_2261#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_65/a_27_74# prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_29/a_222_392#
+ prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_43/a_112_119# prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_19/X
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_25/a_1226_296# prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_31/a_376_368#
+ prbs_generator_syn_13/sky130_fd_sc_hs__or2_1_1/a_63_368# prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_17/a_230_79#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_4/a_27_74# prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_61/a_230_79#
+ prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_63/a_138_385# prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_5/a_222_392#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_8/a_1141_508# prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_41/a_293_74#
+ prbs_generator_syn_13/sky130_fd_sc_hs__nand2_1_31/a_117_74# prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_5/a_138_385#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_63/a_1141_508# prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_19/a_222_392#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_13/a_1141_508# prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_3/a_52_123#
+ prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_13/a_52_123# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_43/a_1178_124#
+ prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_61/a_376_368# prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_35/a_132_392#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_67/a_206_368# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_1/a_1226_296#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_69/a_696_458# prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_31/a_230_79#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_35/a_735_102# prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_23/a_112_119#
+ prbs_generator_syn_13/sky130_fd_sc_hs__nand2_1_35/a_117_74# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_59/a_27_74#
+ prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_13/a_293_74# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_5/a_206_368#
+ prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_50/a_376_368# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_7/a_696_458#
+ prbs_generator_syn_13/sky130_fd_sc_hs__nor2b_1_7/a_278_368# prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_17/a_52_123#
+ prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_43/a_138_385# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_7/a_1141_508#
+ prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_61/a_52_123# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_67/a_437_503#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_61/a_1141_508# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_25/a_735_102#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_59/a_696_458# prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_13/a_112_119#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_33/a_1034_424# prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_51/a_112_119#
+ prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_35/a_230_79# prbs_generator_syn_13/m3_13600_4091#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_23/a_1226_296# prbs_generator_syn_13/sky130_fd_sc_hs__nand2_1_39/a_117_74#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_29/a_27_74# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_5/a_437_503#
+ prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_17/a_293_74# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_41/a_1178_124#
+ prbs_generator_syn_13/sky130_fd_sc_hs__or2_1_1/a_152_368# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_59/a_1178_124#
+ prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_61/a_293_74# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_47/a_206_368#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_39/a_651_503# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_49/a_696_458#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_15/a_735_102# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_32/a_1034_424#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_73/a_1226_296# prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_27/a_222_392#
+ prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_41/a_112_119# prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_31/a_52_123#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_49/a_1034_424# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_29/a_1141_508#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_21/a_1226_296# prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_39/a_230_79#
+ prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_23/a_138_385# prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_51/a_230_79#
+ prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_45/a_132_392# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_37/a_206_368#
+ prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_65/a_293_74# prbs_generator_syn_13/sky130_fd_sc_hs__nand2_1_53/a_117_74#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_47/a_437_503# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_29/a_651_503#
+ prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_31/a_293_74# prbs_generator_syn_13/sky130_fd_sc_hs__nand2_1_21/a_117_74#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_69/a_544_485# prbs_generator_syn_13/sky130_fd_sc_hs__clkbuf_16_1/a_114_74#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_45/a_735_102# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_13/a_27_74#
+ prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_31/a_112_119# prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_57/a_222_392#
+ prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_35/a_52_123# prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_21/a_376_368#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_7/a_544_485# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_57/a_1178_124#
+ prbs_generator_syn_13/m3_13600_6043# prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_13/a_138_385#
+ prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_51/a_138_385# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_5/a_1141_508#
+ prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_3/a_376_368# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_27/a_206_368#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_65/a_206_368# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_37/a_437_503#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_19/a_651_503# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_57/a_651_503#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_59/a_544_485# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_71/a_1226_296#
+ prbs_generator_syn_13/sky130_fd_sc_hs__nand2_1_25/a_117_74# prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_61/a_112_119#
+ prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_47/a_222_392# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_27/a_1141_508#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_53/a_27_74# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_4/a_206_368#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_39/a_1226_296# prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_11/a_376_368#
+ prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_39/a_52_123# prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_41/a_138_385#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_4/a_1141_508# prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_25/a_132_392#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_17/a_206_368# prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_41/A
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_55/a_206_368# prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_51/a_52_123#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_27/a_437_503# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_65/a_437_503#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_49/a_544_485# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_63/a_735_102#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_47/a_1034_424# prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_50/a_112_119#
+ prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_37/a_222_392# prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_59/a_230_79#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_25/a_1141_508# prbs_generator_syn_13/sky130_fd_sc_hs__nor2b_1_4/a_27_112#
+ prbs_generator_syn_13/sky130_fd_sc_hs__sdlclkp_2_1/a_685_81# prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_1/a_132_392#
+ prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_39/a_293_74# prbs_generator_syn_13/sky130_fd_sc_hs__nand2_1_29/a_117_74#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_4/a_437_503# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_55/a_1178_124#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_21/a_27_74# prbs_generator_syn_13/m3_13600_12875#
+ prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_50/a_293_74# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_1/a_735_102#
+ prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_31/a_138_385# prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_15/a_132_392#
+ prbs_generator_syn_13/sky130_fd_sc_hs__nand2_1_1/a_117_74# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_17/a_437_503#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_55/a_437_503# prbs_generator_syn
Xprbs_generator_syn_23 prbs_generator_syn_31/clk prbs_generator_syn_31/rst prbs_generator_syn_23/cke
+ sky130_fd_sc_hs__conb_1_231/LO sky130_fd_sc_hs__conb_1_231/LO sky130_fd_sc_hs__conb_1_231/HI
+ prbs_generator_syn_27/eqn[1] prbs_generator_syn_27/eqn[8] sky130_fd_sc_hs__conb_1_231/LO
+ sky130_fd_sc_hs__conb_1_231/LO sky130_fd_sc_hs__conb_1_231/LO sky130_fd_sc_hs__conb_1_231/LO
+ sky130_fd_sc_hs__conb_1_231/LO sky130_fd_sc_hs__conb_1_231/LO prbs_generator_syn_23/eqn[31]
+ prbs_generator_syn_23/cke prbs_generator_syn_23/eqn[31] sky130_fd_sc_hs__conb_1_233/HI
+ sky130_fd_sc_hs__conb_1_233/HI sky130_fd_sc_hs__conb_1_233/HI prbs_generator_syn_27/eqn[9]
+ sky130_fd_sc_hs__conb_1_187/HI prbs_generator_syn_29/eqn[22] prbs_generator_syn_29/eqn[20]
+ prbs_generator_syn_29/eqn[22] prbs_generator_syn_29/eqn[20] sky130_fd_sc_hs__conb_1_191/HI
+ prbs_generator_syn_29/eqn[28] sky130_fd_sc_hs__conb_1_191/HI prbs_generator_syn_29/eqn[28]
+ prbs_generator_syn_29/cke prbs_generator_syn_29/eqn[31] prbs_generator_syn_29/cke
+ prbs_generator_syn_29/eqn[31] prbs_generator_syn_29/cke prbs_generator_syn_23/eqn[31]
+ prbs_generator_syn_23/eqn[30] prbs_generator_syn_23/eqn[30] prbs_generator_syn_23/eqn[28]
+ prbs_generator_syn_23/eqn[28] prbs_generator_syn_23/eqn[28] prbs_generator_syn_23/eqn[28]
+ prbs_generator_syn_23/eqn[28] prbs_generator_syn_23/eqn[28] prbs_generator_syn_23/eqn[22]
+ prbs_generator_syn_23/eqn[22] prbs_generator_syn_23/eqn[20] prbs_generator_syn_23/eqn[22]
+ prbs_generator_syn_23/eqn[22] prbs_generator_syn_23/eqn[22] prbs_generator_syn_23/eqn[22]
+ prbs_generator_syn_21/eqn[0] prbs_generator_syn_21/eqn[0] prbs_generator_syn_21/eqn[0]
+ prbs_generator_syn_21/eqn[0] prbs_generator_syn_21/eqn[0] prbs_generator_syn_21/eqn[0]
+ prbs_generator_syn_23/eqn[9] prbs_generator_syn_23/eqn[8] prbs_generator_syn_23/eqn[8]
+ prbs_generator_syn_23/eqn[8] prbs_generator_syn_23/eqn[8] prbs_generator_syn_23/eqn[8]
+ prbs_generator_syn_23/eqn[8] prbs_generator_syn_23/eqn[8] prbs_generator_syn_23/eqn[1]
+ prbs_generator_syn_23/eqn[0] prbs_generator_syn_31/inj_err prbs_generator_syn_23/eqn[31]
+ prbs_generator_syn_23/eqn[31] hr_16t4_mux_top_1/din[2] DVSS: DVDD: prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_1/a_293_74#
+ prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_15/X prbs_generator_syn_23/sky130_fd_sc_hs__nand2_1_35/B
+ prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_51/Y prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_9/A
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_9/CLK prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_47/a_27_74#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_37/a_1226_296# prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_3/B
+ prbs_generator_syn_23/sky130_fd_sc_hs__nor2b_1_7/a_27_112# prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_29/B
+ prbs_generator_syn_23/sky130_fd_sc_hs__sdlclkp_2_1/a_580_74# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_1/a_1141_508#
+ prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_5/Y prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_41/a_230_79#
+ prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_61/a_138_385# prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_43/a_132_392#
+ prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_3/a_222_392# prbs_generator_syn_23/sky130_fd_sc_hs__nor2b_1_9/a_27_112#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_61/a_27_74# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_35/a_206_368#
+ prbs_generator_syn_23/sky130_fd_sc_hs__nand2_2_3/Y prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_25/B
+ prbs_generator_syn_23/sky130_fd_sc_hs__nand2_1_11/a_117_74# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_67/a_651_503#
+ prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_45/X prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_39/a_696_458#
+ prbs_generator_syn_23/sky130_fd_sc_hs__sdlclkp_2_1/a_1198_74# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_45/a_1034_424#
+ prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_17/a_222_392# prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_55/a_222_392#
+ prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_53/Y prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_35/A
+ prbs_generator_syn_23/m3_13600_1651# prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_59/a_52_123#
+ prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_5/a_293_74# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_35/a_1226_296#
+ prbs_generator_syn_23/sky130_fd_sc_hs__nand2_1_51/B prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_5/a_651_503#
+ prbs_generator_syn_23/sky130_fd_sc_hs__nand2_1_21/B prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_8/a_27_74#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_15/a_27_74# prbs_generator_syn_23/sky130_fd_sc_hs__and2b_2_1/X
+ prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_13/X prbs_generator_syn_23/sky130_fd_sc_hs__nand2_2_3/a_27_74#
+ prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_50/a_138_385# prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_33/a_132_392#
+ prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_1/a_376_368# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_25/a_206_368#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_35/a_437_503# prbs_generator_syn_23/sky130_fd_sc_hs__sdlclkp_2_1/a_708_451#
+ prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_45/a_230_79# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_29/a_696_458#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_32/a_27_74# prbs_generator_syn_23/sky130_fd_sc_hs__nor2b_1_4/Y
+ prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_59/a_293_74# prbs_generator_syn_23/sky130_fd_sc_hs__nand2_1_47/a_117_74#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_73/a_735_102# prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_21/a_112_119#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_23/a_1141_508# prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_25/a_293_74#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_7/Q prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_3/a_112_119#
+ prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_35/B prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_51/X
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_53/a_1178_124# prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_23/a_132_392#
+ prbs_generator_syn_23/sky130_fd_sc_hs__nand2_1_3/B prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_15/a_206_368#
+ prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_63/a_132_392# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_55/a_27_74#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_25/a_437_503# prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_41/a_52_123#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_47/a_651_503# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_73/a_1141_508#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_19/a_696_458# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_57/a_696_458#
+ prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_7/X prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_43/a_1034_424#
+ prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_55/A prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_11/a_112_119#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_21/a_1141_508# prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_35/a_222_392#
+ prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_49/a_230_79# prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_67/Y
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_71/a_27_74# prbs_generator_syn_23/sky130_fd_sc_hs__nand2_1_33/B
+ prbs_generator_syn_23/sky130_fd_sc_hs__conb_1_1/LO prbs_generator_syn_23/sky130_fd_sc_hs__nand2_1_19/a_117_74#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_51/a_1178_124# prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_33/X
+ prbs_generator_syn_23/sky130_fd_sc_hs__nand2_1_29/B prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_41/Y
+ prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_53/a_132_392# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_45/a_206_368#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_15/a_437_503# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_37/a_651_503#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_39/a_544_485# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_53/a_735_102#
+ prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_45/a_52_123# prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_1/B
+ prbs_generator_syn_23/sky130_fd_sc_hs__nand2_2_3/B prbs_generator_syn_23/sky130_fd_sc_hs__clkbuf_16_1/A
+ prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_21/X prbs_generator_syn_23/sky130_fd_sc_hs__nand2_1_25/B
+ prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_39/a_376_368# prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_63/X
+ prbs_generator_syn_23/m3_13600_3481# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_69/a_1178_124#
+ prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_21/a_138_385# prbs_generator_syn_23/sky130_fd_sc_hs__nor2b_1_8/Y
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_19/a_1178_124# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_49/a_27_74#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_45/a_437_503# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_27/a_651_503#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_71/a_1141_508# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_65/a_651_503#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_29/a_544_485# prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_3/a_138_385#
+ prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_55/X prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_43/a_735_102#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_41/a_1034_424# prbs_generator_syn_23/sky130_fd_sc_hs__nand2_1_9/B
+ prbs_generator_syn_23/sky130_fd_sc_hs__nor2b_1_9/Y prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_59/a_1034_424#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_39/a_1141_508# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_33/a_1226_296#
+ prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_49/a_52_123# prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_47/Y
+ prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_43/Y prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_4/a_651_503#
+ prbs_generator_syn_23/sky130_fd_sc_hs__nand2_1_49/B prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_19/A
+ prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_11/a_138_385# prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_5/X
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_63/a_206_368# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_17/a_651_503#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_19/a_544_485# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_55/a_651_503#
+ prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_9/Y prbs_generator_syn_23/sky130_fd_sc_hs__nand2_1_17/B
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_57/a_544_485# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_67/a_696_458#
+ prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_35/X prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_19/a_27_74#
+ prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_45/a_222_392# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_32/a_1226_296#
+ prbs_generator_syn_23/sky130_fd_sc_hs__nand2_1_43/B prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_25/A
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_1/a_206_368# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_49/a_1226_296#
+ prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_1/a_112_119# prbs_generator_syn_23/sky130_fd_sc_hs__or2_1_1/X
+ prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_59/a_376_368# prbs_generator_syn_23/sky130_fd_sc_hs__nand2_1_19/B
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_5/a_696_458# prbs_generator_syn_23/sky130_fd_sc_hs__nor2b_1_1/Y
+ prbs_generator_syn_23/sky130_fd_sc_hs__nor2b_1_5/a_278_368# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_17/a_1178_124#
+ prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_39/X prbs_generator_syn_23/m3_13600_5433#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_63/a_437_503# prbs_generator_syn_23/sky130_fd_sc_hs__nand2_2_5/B
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_23/a_735_102# prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_53/A
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_61/a_735_102# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_57/a_1034_424#
+ prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_63/B prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_37/a_1141_508#
+ prbs_generator_syn_23/sky130_fd_sc_hs__nand2_1_47/B prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_29/X
+ prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_65/Y prbs_generator_syn_23/m3_13600_4701#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_1/a_437_503# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_67/a_1178_124#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_9/a_735_102# prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_13/a_132_392#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_15/a_1178_124# prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_15/A
+ prbs_generator_syn_23/sky130_fd_sc_hs__nand2_1_1/B prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_43/B
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_35/a_651_503# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_8/D
+ prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_29/A prbs_generator_syn_23/sky130_fd_sc_hs__nand2_1_7/B
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_13/a_735_102# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_47/a_696_458#
+ prbs_generator_syn_23/sky130_fd_sc_hs__nand2_1_31/B prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_51/a_735_102#
+ prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_59/X prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_35/a_1141_508#
+ prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_25/a_222_392# prbs_generator_syn_23/sky130_fd_sc_hs__sdlclkp_2_1/a_288_48#
+ prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_55/B prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_17/B
+ prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_43/A prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_7/A
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_65/a_1178_124# prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_59/Y
+ prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_41/X prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_21/a_230_79#
+ prbs_generator_syn_23/sky130_fd_sc_hs__nand2_1_57/a_117_74# prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_1/a_222_392#
+ prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_19/B prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_35/a_293_74#
+ prbs_generator_syn_23/sky130_fd_sc_hs__nand2_1_23/a_117_74# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_73/a_206_368#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_25/a_651_503# prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_1/a_138_385#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_37/a_696_458# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_67/a_544_485#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_43/a_27_74# prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_9/X
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_55/a_1034_424# prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_39/a_112_119#
+ prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_15/a_222_392# prbs_generator_syn_23/sky130_fd_sc_hs__conb_1_1/HI
+ prbs_generator_syn_23/sky130_fd_sc_hs__nand2_1_23/B prbs_generator_syn_23/sky130_fd_sc_hs__nand2_1_53/B
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_9/a_1178_124# prbs_generator_syn_23/sky130_fd_sc_hs__nor2b_1_4/A
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_47/a_1226_296# prbs_generator_syn_23/m3_13600_11045#
+ prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_17/X prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_29/a_376_368#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_5/a_544_485# prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_3/X
+ prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_31/a_132_392# prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_61/A
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_15/a_651_503# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_73/a_437_503#
+ prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_25/a_230_79# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_27/a_696_458#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_65/a_696_458# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_33/a_735_102#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_71/a_735_102# prbs_generator_syn_23/m3_13600_7263#
+ prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_43/a_222_392# prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_50/Y
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_8/a_1178_124# prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_53/B
+ prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_19/a_376_368# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_63/a_1178_124#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_4/a_696_458# prbs_generator_syn_23/sky130_fd_sc_hs__nor2b_1_4/a_278_368#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_13/a_1178_124# prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_61/a_132_392#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_53/a_206_368# prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_21/a_52_123#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_45/a_651_503# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_17/a_696_458#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_47/a_544_485# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_55/a_696_458#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_21/a_735_102# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_37/a_27_74#
+ prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_61/B prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_61/X
+ prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_59/a_112_119# prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_31/A
+ prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_33/a_222_392# prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_29/a_230_79#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_45/a_1226_296# prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_9/a_132_392#
+ prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_5/A prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_57/Y
+ prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_31/X prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_51/a_27_74#
+ prbs_generator_syn_23/sky130_fd_sc_hs__nor2b_1_8/a_27_112# prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_47/a_376_368#
+ prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_53/a_293_74# prbs_generator_syn_23/sky130_fd_sc_hs__nand2_1_43/a_117_74#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_8/a_735_102# prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_21/a_293_74#
+ prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_39/a_138_385# prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_63/Y
+ prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_51/a_132_392# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_43/a_206_368#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_53/a_437_503# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_37/a_544_485#
+ prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_57/X prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_53/a_1034_424#
+ prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_25/a_52_123# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_33/a_1141_508#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_63/Q prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_23/a_222_392#
+ prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_63/a_222_392# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_7/a_1178_124#
+ prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_53/X prbs_generator_syn_23/sky130_fd_sc_hs__nand2_2_5/Y
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_61/a_1178_124# prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_1/a_230_79#
+ prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_43/a_230_79# prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_11/a_230_79#
+ prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_41/a_132_392# prbs_generator_syn_23/sky130_fd_sc_hs__nand2_1_13/a_117_74#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_43/a_437_503# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_27/a_544_485#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_63/a_651_503# prbs_generator_syn_23/sky130_fd_sc_hs__nand2_1_7/a_117_74#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_35/a_696_458# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_65/a_544_485#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_51/a_1034_424# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_41/a_735_102#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_32/a_1141_508# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_49/a_1141_508#
+ prbs_generator_syn_23/sky130_fd_sc_hs__nand2_1_55/B prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_53/a_222_392#
+ prbs_generator_syn_23/sky130_fd_sc_hs__sdlclkp_2_1/a_114_112# prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_9/a_293_74#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_43/a_1226_296# prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_29/a_52_123#
+ prbs_generator_syn_23/sky130_fd_sc_hs__nand2_1_37/B prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_1/a_651_503#
+ prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_27/a_376_368# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_4/a_544_485#
+ prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_67/a_376_368# prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_27/X
+ prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_1/X prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_59/a_138_385#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_29/a_1178_124# prbs_generator_syn_23/m3_13600_2871#
+ prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_5/a_230_79# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_23/a_206_368#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_61/a_206_368# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_17/a_544_485#
+ prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_15/a_230_79# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_25/a_696_458#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_55/a_544_485# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_32/a_735_102#
+ prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_29/a_293_74# prbs_generator_syn_23/sky130_fd_sc_hs__nand2_1_17/a_117_74#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_69/a_1034_424# prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_29/a_112_119#
+ prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_37/X prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_31/B
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_19/a_1034_424# prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_33/A
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_9/a_206_368# prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_57/a_376_368#
+ prbs_generator_syn_23/sky130_fd_sc_hs__sdlclkp_2_1/a_706_317# prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_11/B
+ prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_1/a_52_123# prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_39/B
+ prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_21/a_132_392# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_13/a_206_368#
+ prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_43/a_52_123# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_51/a_206_368#
+ prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_47/X prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_23/a_437_503#
+ prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_11/a_52_123# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_61/a_437_503#
+ prbs_generator_syn_23/sky130_fd_sc_hs__nor2b_1_7/Y prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_51/A
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_15/a_696_458# prbs_generator_syn_23/sky130_fd_sc_hs__nor2b_1_5/Y
+ prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_9/a_230_79# prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_25/X
+ prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_19/a_112_119# prbs_generator_syn_23/sky130_fd_sc_hs__nand2_1_45/B
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_5/a_1178_124# prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_19/a_230_79#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_41/a_1226_296# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_59/a_1226_296#
+ prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_63/a_230_79# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_51/Q
+ prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_7/a_132_392# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_9/a_437_503#
+ prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_46/a_376_368# prbs_generator_syn_23/sky130_fd_sc_hs__nand2_1_33/a_117_74#
+ prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_11/a_293_74# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_27/a_1178_124#
+ prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_11/a_132_392# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_13/a_437_503#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_51/a_437_503# prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_5/a_52_123#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_35/a_544_485# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_73/a_651_503#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_45/a_696_458# prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_15/a_52_123#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_47/a_1141_508# prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_47/a_112_119#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_4/a_1178_124# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_17/a_1034_424#
+ prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_23/B prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_37/a_376_368#
+ prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_15/B prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_7/Y
+ prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_29/a_138_385# prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_33/a_230_79#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_25/a_1178_124# prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_47/a_293_74#
+ prbs_generator_syn_23/sky130_fd_sc_hs__nand2_1_37/a_117_74# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_33/a_206_368#
+ prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_15/a_293_74# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_71/a_206_368#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_25/a_544_485# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_67/a_1034_424#
+ prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_13/a_222_392# prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_9/a_52_123#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_15/a_1034_424# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_57/a_1226_296#
+ prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_19/a_52_123# prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_23/X
+ prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_63/a_52_123# prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_19/a_138_385#
+ prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_9/a_376_368# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_21/a_206_368#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_33/a_437_503# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_71/a_437_503#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_53/a_651_503# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_15/a_544_485#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_63/a_696_458# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_65/a_1034_424#
+ prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_19/a_293_74# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_45/a_1141_508#
+ prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_27/a_112_119# prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_67/a_112_119#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_1/a_1178_124# prbs_generator_syn_23/sky130_fd_sc_hs__conb_1_1/a_21_290#
+ prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_63/a_293_74# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_8/a_206_368#
+ prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_17/a_376_368# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_63/a_27_74#
+ prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_21/A prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_55/a_376_368#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_1/a_696_458# prbs_generator_syn_23/sky130_fd_sc_hs__nor2b_1_1/a_278_368#
+ prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_47/a_138_385# prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_33/a_52_123#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_9/a_1034_424# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_21/a_437_503#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_1/a_27_74# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_43/a_651_503#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_1/Q prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_45/a_544_485#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_69/a_735_102# prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_57/a_112_119#
+ prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_31/a_222_392# prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_13/A
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_55/a_1226_296# prbs_generator_syn_23/sky130_fd_sc_hs__nand2_2_5/a_27_74#
+ prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_53/a_230_79# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_8/a_437_503#
+ prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_67/a_293_74# prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_33/a_293_74#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_7/a_735_102# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_23/a_1178_124#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_41/a_206_368# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_8/a_1034_424#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_63/a_1034_424# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_59/a_735_102#
+ prbs_generator_syn_23/sky130_fd_sc_hs__nand2_1_5/B prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_43/a_1141_508#
+ prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_46/a_112_119# prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_61/a_222_392#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_13/a_1034_424# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_73/a_1178_124#
+ prbs_generator_syn_23/sky130_fd_sc_hs__nand2_1_27/B prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_13/B
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_57/a_27_74# prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_57/a_230_79#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_21/a_1178_124# prbs_generator_syn_23/sky130_fd_sc_hs__nor2b_1_1/a_27_112#
+ prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_27/a_138_385# prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_23/a_230_79#
+ prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_67/a_138_385# prbs_generator_syn_23/sky130_fd_sc_hs__nand2_1_41/B
+ prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_9/a_222_392# prbs_generator_syn_23/sky130_fd_sc_hs__nand2_1_27/a_117_74#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_32/a_206_368# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_23/a_651_503#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_41/a_437_503# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_73/a_27_74#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_61/a_651_503# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_63/a_544_485#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_49/a_735_102# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_73/a_696_458#
+ prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_37/a_112_119# prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_51/a_222_392#
+ prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_43/X prbs_generator_syn_23/sky130_fd_sc_hs__nand2_2_1/B
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_9/a_651_503# prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_53/a_52_123#
+ prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_49/X prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_25/a_376_368#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_1/a_544_485# prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_65/a_376_368#
+ prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_57/a_138_385# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_27/a_27_74#
+ prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_39/a_132_392# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_7/a_1034_424#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_13/a_651_503# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_32/a_437_503#
+ prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_27/a_230_79# prbs_generator_syn_23/m3_13600_12265#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_51/a_651_503# prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_59/B
+ prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_47/A prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_61/a_1034_424#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_41/a_1141_508# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_59/a_1141_508#
+ prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_41/a_222_392# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_53/a_1226_296#
+ prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_3/A prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_71/a_1178_124#
+ prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_9/a_112_119# prbs_generator_syn_23/sky130_fd_sc_hs__nand2_1_3/a_117_74#
+ prbs_generator_syn_23/m3_13600_8483# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_39/a_1178_124#
+ prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_57/a_52_123# prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_46/a_138_385#
+ prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_23/a_52_123# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_67/a_27_74#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_53/a_696_458# prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_17/a_112_119#
+ prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_11/A prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_55/a_112_119#
+ prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_1/A prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_51/a_1226_296#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_29/a_1034_424# prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_59/A
+ prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_23/A prbs_generator_syn_23/sky130_fd_sc_hs__nand2_1_39/B
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_5/a_27_74# prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_57/a_293_74#
+ prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_37/a_138_385# prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_59/a_132_392#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_33/a_651_503# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_71/a_651_503#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_43/a_696_458# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_73/a_544_485#
+ prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_27/a_52_123# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_57/a_1141_508#
+ prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_21/a_222_392# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_35/a_27_74#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_69/a_1226_296# prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_37/B
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_19/a_1226_296# prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_35/a_376_368#
+ prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_47/a_230_79# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_37/a_1178_124#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_5/a_1034_424# prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_49/a_132_392#
+ prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_7/a_222_392# prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_27/a_293_74#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_21/a_651_503# prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_9/a_138_385#
+ prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_11/a_222_392# prbs_generator_syn_23/m3_13600_14095#
+ prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_50/A prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_27/a_1034_424#
+ prbs_generator_syn_23/sky130_fd_sc_hs__nand2_1_13/B prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_8/a_651_503#
+ prbs_generator_syn_23/m3_13600_9703# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_35/a_1178_124#
+ prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_17/a_138_385# prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_55/a_138_385#
+ prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_7/a_230_79# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_4/a_1034_424#
+ prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_7/a_376_368# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_69/a_206_368#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_23/a_696_458# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_53/a_544_485#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_39/a_735_102# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_61/a_696_458#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_55/a_1141_508# prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_25/a_112_119#
+ prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_65/a_112_119# prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_43/a_293_74#
+ prbs_generator_syn_23/sky130_fd_sc_hs__nand2_1_57/B prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_25/a_1034_424#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_7/a_206_368# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_17/a_1226_296#
+ prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_15/a_376_368# prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_53/a_376_368#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_9/a_696_458# prbs_generator_syn_23/m3_13600_431#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_45/a_27_74# prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_47/a_52_123#
+ prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_29/a_132_392# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_59/a_206_368#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_69/a_437_503# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_41/a_651_503#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_43/a_544_485# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_13/a_696_458#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_29/a_735_102# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_51/a_696_458#
+ prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_61/Y prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_67/a_1226_296#
+ prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_5/a_132_392# prbs_generator_syn_23/sky130_fd_sc_hs__and2b_2_1/a_198_48#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_7/a_437_503# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_15/a_1226_296#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_69/a_27_74# prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_46/a_293_74#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_1/a_1034_424# prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_19/a_132_392#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_49/a_206_368# prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_7/a_52_123#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_59/a_437_503# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_32/a_651_503#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_7/a_27_74# prbs_generator_syn_23/sky130_fd_sc_hs__nand2_2_1/a_27_74#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_19/a_735_102# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_57/a_735_102#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_65/a_1226_296# prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_37/A
+ prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_33/a_376_368# prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_37/a_230_79#
+ prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_25/a_138_385# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_39/a_27_74#
+ prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_65/a_138_385# prbs_generator_syn_23/sky130_fd_sc_hs__nor2b_1_9/a_278_368#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_49/a_437_503# prbs_generator_syn_23/sky130_fd_sc_hs__and2b_2_1/a_505_74#
+ prbs_generator_syn_23/sky130_fd_sc_hs__nand2_1_51/a_117_74# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_23/a_544_485#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_33/a_696_458# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_61/a_544_485#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_9/a_1226_296# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_53/a_1141_508#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_71/a_696_458# prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_35/a_112_119#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_23/a_1034_424# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_9/a_544_485#
+ prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_63/a_376_368# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_33/a_1178_124#
+ prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_5/a_376_368# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_13/a_544_485#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_73/a_1034_424# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_21/a_696_458#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_51/a_544_485# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_8/a_1226_296#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_51/a_1141_508# prbs_generator_syn_23/sky130_fd_sc_hs__nand2_1_55/a_117_74#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_21/a_1034_424# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_63/a_1226_296#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_23/a_27_74# prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_7/a_112_119#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_13/a_1226_296# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_8/a_696_458#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_32/a_1178_124# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_49/a_1178_124#
+ prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_37/a_52_123# prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_27/a_132_392#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_71/Q prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_67/a_735_102#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_69/a_1141_508# prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_15/a_112_119#
+ prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_53/a_112_119# prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_39/a_222_392#
+ prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_55/a_230_79# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_19/a_1141_508#
+ prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_37/a_293_74# prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_43/a_376_368#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_5/a_735_102# prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_35/a_138_385#
+ prbs_generator_syn_23/sky130_fd_sc_hs__sdlclkp_2_1/a_114_424# prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_57/a_132_392#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_71/a_1034_424# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_7/a_1226_296#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_33/a_544_485# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_41/a_696_458#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_71/a_544_485# prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_21/B
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_61/a_1226_296# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_39/a_1034_424#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_17/a_27_74# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_9/a_27_74#
+ prbs_generator_syn_23/sky130_fd_sc_hs__nor2b_1_5/a_27_112# prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_47/a_132_392#
+ prbs_generator_syn_23/sky130_fd_sc_hs__nor2b_1_8/a_278_368# prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_9/B
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_39/a_206_368# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_33/a_27_74#
+ prbs_generator_syn_23/sky130_fd_sc_hs__nand2_1_41/a_117_74# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_69/a_651_503#
+ prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_51/a_293_74# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_21/a_544_485#
+ prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_7/a_138_385# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_32/a_696_458#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_47/a_735_102# prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_33/a_112_119#
+ prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_59/a_222_392# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_17/a_1141_508#
+ prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_55/a_52_123# prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_3/a_293_74#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_7/a_651_503# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_29/a_1226_296#
+ prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_23/a_376_368# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_8/a_544_485#
+ prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_47/B prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_47/a_1178_124#
+ prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_15/a_138_385# prbs_generator_syn_23/sky130_fd_sc_hs__sdlclkp_2_1/a_1195_374#
+ prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_53/a_138_385# prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_37/a_132_392#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_29/a_206_368# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_39/a_437_503#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_59/a_651_503# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_37/a_735_102#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_67/a_1141_508# prbs_generator_syn_23/sky130_fd_sc_hs__and2b_2_1/a_27_74#
+ prbs_generator_syn_23/sky130_fd_sc_hs__conb_1_1/a_165_290# prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_55/a_293_74#
+ prbs_generator_syn_23/sky130_fd_sc_hs__nand2_1_45/a_117_74# prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_63/a_112_119#
+ prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_49/a_222_392# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_37/a_1034_424#
+ prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_23/a_293_74# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_15/a_1141_508#
+ prbs_generator_syn_23/sky130_fd_sc_hs__nand2_1_5/a_117_74# prbs_generator_syn_23/m3_13600_13485#
+ prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_5/a_112_119# prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_13/a_376_368#
+ prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_51/a_376_368# prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_7/a_293_74#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_19/a_206_368# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_57/a_206_368#
+ prbs_generator_syn_23/sky130_fd_sc_hs__sdlclkp_2_1/a_318_74# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_29/a_437_503#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_49/a_651_503# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_25/a_27_74#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_5/a_1226_296# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_41/a_544_485#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_27/a_735_102# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_65/a_1141_508#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_65/a_735_102# prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_3/a_230_79#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_35/a_1034_424# prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_13/a_230_79#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_41/a_27_74# prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_3/a_132_392#
+ prbs_generator_syn_23/sky130_fd_sc_hs__nand2_1_49/a_117_74# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_27/a_1226_296#
+ prbs_generator_syn_23/sky130_fd_sc_hs__nand2_1_15/a_117_74# prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_41/a_376_368#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_45/a_1178_124# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_4/a_735_102#
+ prbs_generator_syn_23/sky130_fd_sc_hs__nand2_1_9/a_117_74# prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_33/a_138_385#
+ prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_17/a_132_392# prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_55/a_132_392#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_9/a_1141_508# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_19/a_437_503#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_57/a_437_503# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_4/a_1226_296#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_32/a_544_485# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_17/a_735_102#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_55/a_735_102# prbs_generator_syn_23/m3_13600_2261#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_65/a_27_74# prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_29/a_222_392#
+ prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_43/a_112_119# prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_19/X
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_25/a_1226_296# prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_31/a_376_368#
+ prbs_generator_syn_23/sky130_fd_sc_hs__or2_1_1/a_63_368# prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_17/a_230_79#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_4/a_27_74# prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_61/a_230_79#
+ prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_63/a_138_385# prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_5/a_222_392#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_8/a_1141_508# prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_41/a_293_74#
+ prbs_generator_syn_23/sky130_fd_sc_hs__nand2_1_31/a_117_74# prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_5/a_138_385#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_63/a_1141_508# prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_19/a_222_392#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_13/a_1141_508# prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_3/a_52_123#
+ prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_13/a_52_123# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_43/a_1178_124#
+ prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_61/a_376_368# prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_35/a_132_392#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_67/a_206_368# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_1/a_1226_296#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_69/a_696_458# prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_31/a_230_79#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_35/a_735_102# prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_23/a_112_119#
+ prbs_generator_syn_23/sky130_fd_sc_hs__nand2_1_35/a_117_74# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_59/a_27_74#
+ prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_13/a_293_74# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_5/a_206_368#
+ prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_50/a_376_368# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_7/a_696_458#
+ prbs_generator_syn_23/sky130_fd_sc_hs__nor2b_1_7/a_278_368# prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_17/a_52_123#
+ prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_43/a_138_385# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_7/a_1141_508#
+ prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_61/a_52_123# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_67/a_437_503#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_61/a_1141_508# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_25/a_735_102#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_59/a_696_458# prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_13/a_112_119#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_33/a_1034_424# prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_51/a_112_119#
+ prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_35/a_230_79# prbs_generator_syn_23/m3_13600_4091#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_23/a_1226_296# prbs_generator_syn_23/sky130_fd_sc_hs__nand2_1_39/a_117_74#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_29/a_27_74# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_5/a_437_503#
+ prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_17/a_293_74# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_41/a_1178_124#
+ prbs_generator_syn_23/sky130_fd_sc_hs__or2_1_1/a_152_368# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_59/a_1178_124#
+ prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_61/a_293_74# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_47/a_206_368#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_39/a_651_503# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_49/a_696_458#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_15/a_735_102# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_32/a_1034_424#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_73/a_1226_296# prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_27/a_222_392#
+ prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_41/a_112_119# prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_31/a_52_123#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_49/a_1034_424# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_29/a_1141_508#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_21/a_1226_296# prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_39/a_230_79#
+ prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_23/a_138_385# prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_51/a_230_79#
+ prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_45/a_132_392# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_37/a_206_368#
+ prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_65/a_293_74# prbs_generator_syn_23/sky130_fd_sc_hs__nand2_1_53/a_117_74#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_47/a_437_503# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_29/a_651_503#
+ prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_31/a_293_74# prbs_generator_syn_23/sky130_fd_sc_hs__nand2_1_21/a_117_74#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_69/a_544_485# prbs_generator_syn_23/sky130_fd_sc_hs__clkbuf_16_1/a_114_74#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_45/a_735_102# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_13/a_27_74#
+ prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_31/a_112_119# prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_57/a_222_392#
+ prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_35/a_52_123# prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_21/a_376_368#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_7/a_544_485# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_57/a_1178_124#
+ prbs_generator_syn_23/m3_13600_6043# prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_13/a_138_385#
+ prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_51/a_138_385# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_5/a_1141_508#
+ prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_3/a_376_368# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_27/a_206_368#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_65/a_206_368# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_37/a_437_503#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_19/a_651_503# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_57/a_651_503#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_59/a_544_485# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_71/a_1226_296#
+ prbs_generator_syn_23/sky130_fd_sc_hs__nand2_1_25/a_117_74# prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_61/a_112_119#
+ prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_47/a_222_392# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_27/a_1141_508#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_53/a_27_74# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_4/a_206_368#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_39/a_1226_296# prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_11/a_376_368#
+ prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_39/a_52_123# prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_41/a_138_385#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_4/a_1141_508# prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_25/a_132_392#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_17/a_206_368# prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_41/A
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_55/a_206_368# prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_51/a_52_123#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_27/a_437_503# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_65/a_437_503#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_49/a_544_485# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_63/a_735_102#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_47/a_1034_424# prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_50/a_112_119#
+ prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_37/a_222_392# prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_59/a_230_79#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_25/a_1141_508# prbs_generator_syn_23/sky130_fd_sc_hs__nor2b_1_4/a_27_112#
+ prbs_generator_syn_23/sky130_fd_sc_hs__sdlclkp_2_1/a_685_81# prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_1/a_132_392#
+ prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_39/a_293_74# prbs_generator_syn_23/sky130_fd_sc_hs__nand2_1_29/a_117_74#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_4/a_437_503# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_55/a_1178_124#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_21/a_27_74# prbs_generator_syn_23/m3_13600_12875#
+ prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_50/a_293_74# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_1/a_735_102#
+ prbs_generator_syn_23/sky130_fd_sc_hs__xnor2_1_31/a_138_385# prbs_generator_syn_23/sky130_fd_sc_hs__a22o_1_15/a_132_392#
+ prbs_generator_syn_23/sky130_fd_sc_hs__nand2_1_1/a_117_74# prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_17/a_437_503#
+ prbs_generator_syn_23/sky130_fd_sc_hs__dfxtp_4_55/a_437_503# prbs_generator_syn
Xsky130_fd_sc_hs__conb_1_3 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__conb_1_3/LO sky130_fd_sc_hs__conb_1_3/HI
+ sky130_fd_sc_hs__conb_1_3/a_165_290# sky130_fd_sc_hs__conb_1_3/a_21_290# sky130_fd_sc_hs__conb_1
Xsky130_fd_sc_hs__buf_2_110 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__buf_2_111/A sky130_fd_sc_hs__buf_2_111/X
+ sky130_fd_sc_hs__buf_2_111/a_21_260# sky130_fd_sc_hs__buf_2
Xsky130_fd_sc_hs__buf_2_121 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__buf_2_121/A sky130_fd_sc_hs__buf_2_121/X
+ sky130_fd_sc_hs__buf_2_121/a_21_260# sky130_fd_sc_hs__buf_2
Xsky130_fd_sc_hs__buf_2_132 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__buf_2_133/A sky130_fd_sc_hs__buf_2_133/X
+ sky130_fd_sc_hs__buf_2_133/a_21_260# sky130_fd_sc_hs__buf_2
Xsky130_fd_sc_hs__buf_2_143 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__buf_2_143/A sky130_fd_sc_hs__buf_2_143/X
+ sky130_fd_sc_hs__buf_2_143/a_21_260# sky130_fd_sc_hs__buf_2
Xsky130_fd_sc_hs__buf_2_154 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__buf_2_155/A sky130_fd_sc_hs__buf_2_155/X
+ sky130_fd_sc_hs__buf_2_155/a_21_260# sky130_fd_sc_hs__buf_2
Xsky130_fd_sc_hs__einvp_2_11 DVSS: DVDD: DVDD: DVSS: dout_n sky130_fd_sc_hs__einvp_2_9/A
+ sky130_fd_sc_hs__dlrtp_1_8/Q sky130_fd_sc_hs__einvp_2_11/a_263_323# sky130_fd_sc_hs__einvp_2_11/a_36_74#
+ sky130_fd_sc_hs__einvp_2_11/a_27_368# sky130_fd_sc_hs__einvp_2
Xsky130_fd_sc_hs__einvp_2_22 DVSS: DVDD: DVDD: DVSS: dout_n sky130_fd_sc_hs__einvp_2_9/A
+ sky130_fd_sc_hs__dlrtp_1_17/Q sky130_fd_sc_hs__einvp_2_23/a_263_323# sky130_fd_sc_hs__einvp_2_23/a_36_74#
+ sky130_fd_sc_hs__einvp_2_23/a_27_368# sky130_fd_sc_hs__einvp_2
Xsky130_fd_sc_hs__einvp_2_33 DVSS: DVDD: DVDD: DVSS: dout_n sky130_fd_sc_hs__buf_8_1/A
+ sky130_fd_sc_hs__buf_2_125/X sky130_fd_sc_hs__einvp_2_33/a_263_323# sky130_fd_sc_hs__einvp_2_33/a_36_74#
+ sky130_fd_sc_hs__einvp_2_33/a_27_368# sky130_fd_sc_hs__einvp_2
Xsky130_fd_sc_hs__einvp_2_44 DVSS: DVDD: DVDD: DVSS: dout_n sky130_fd_sc_hs__buf_8_1/A
+ sky130_fd_sc_hs__dlrtp_1_29/Q sky130_fd_sc_hs__einvp_2_45/a_263_323# sky130_fd_sc_hs__einvp_2_45/a_36_74#
+ sky130_fd_sc_hs__einvp_2_45/a_27_368# sky130_fd_sc_hs__einvp_2
Xsky130_fd_sc_hs__einvp_2_55 DVSS: DVDD: DVDD: DVSS: dout_p sky130_fd_sc_hs__inv_4_9/Y
+ sky130_fd_sc_hs__dlrtp_1_39/Q sky130_fd_sc_hs__einvp_2_55/a_263_323# sky130_fd_sc_hs__einvp_2_55/a_36_74#
+ sky130_fd_sc_hs__einvp_2_55/a_27_368# sky130_fd_sc_hs__einvp_2
Xsky130_fd_sc_hs__einvp_2_66 DVSS: DVDD: DVDD: DVSS: dout_p sky130_fd_sc_hs__einvp_2_99/A
+ sky130_fd_sc_hs__dlrtp_1_47/Q sky130_fd_sc_hs__einvp_2_67/a_263_323# sky130_fd_sc_hs__einvp_2_67/a_36_74#
+ sky130_fd_sc_hs__einvp_2_67/a_27_368# sky130_fd_sc_hs__einvp_2
Xsky130_fd_sc_hs__einvp_2_77 DVSS: DVDD: DVDD: DVSS: dout_p sky130_fd_sc_hs__einvp_2_97/A
+ sky130_fd_sc_hs__dlrtp_1_65/Q sky130_fd_sc_hs__einvp_2_77/a_263_323# sky130_fd_sc_hs__einvp_2_77/a_36_74#
+ sky130_fd_sc_hs__einvp_2_77/a_27_368# sky130_fd_sc_hs__einvp_2
Xsky130_fd_sc_hs__einvp_2_88 DVSS: DVDD: DVDD: DVSS: dout_p sky130_fd_sc_hs__einvp_2_97/A
+ sky130_fd_sc_hs__einvp_2_89/TE sky130_fd_sc_hs__einvp_2_89/a_263_323# sky130_fd_sc_hs__einvp_2_89/a_36_74#
+ sky130_fd_sc_hs__einvp_2_89/a_27_368# sky130_fd_sc_hs__einvp_2
Xsky130_fd_sc_hs__einvp_2_99 DVSS: DVDD: DVDD: DVSS: dout_p sky130_fd_sc_hs__einvp_2_99/A
+ sky130_fd_sc_hs__dlrtp_1_81/Q sky130_fd_sc_hs__einvp_2_99/a_263_323# sky130_fd_sc_hs__einvp_2_99/a_36_74#
+ sky130_fd_sc_hs__einvp_2_99/a_27_368# sky130_fd_sc_hs__einvp_2
Xsky130_fd_sc_hs__or2b_2_3 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__or2b_2_3/X sky130_fd_sc_hs__or2b_2_1/A
+ sky130_fd_sc_hs__or2b_2_3/A sky130_fd_sc_hs__or2b_2_3/a_470_368# sky130_fd_sc_hs__or2b_2_3/a_27_368#
+ sky130_fd_sc_hs__or2b_2_3/a_187_48# sky130_fd_sc_hs__or2b_2
Xsky130_fd_sc_hs__conb_1_10 DVSS: DVDD: DVDD: DVSS: prbs_generator_syn_3/eqn[4] prbs_generator_syn_3/eqn[1]
+ sky130_fd_sc_hs__conb_1_11/a_165_290# sky130_fd_sc_hs__conb_1_11/a_21_290# sky130_fd_sc_hs__conb_1
Xsky130_fd_sc_hs__conb_1_21 DVSS: DVDD: DVDD: DVSS: prbs_generator_syn_9/eqn[2] prbs_generator_syn_9/eqn[1]
+ sky130_fd_sc_hs__conb_1_21/a_165_290# sky130_fd_sc_hs__conb_1_21/a_21_290# sky130_fd_sc_hs__conb_1
Xsky130_fd_sc_hs__conb_1_32 DVSS: DVDD: DVDD: DVSS: prbs_generator_syn_5/eqn[31] prbs_generator_syn_5/cke
+ sky130_fd_sc_hs__conb_1_33/a_165_290# sky130_fd_sc_hs__conb_1_33/a_21_290# sky130_fd_sc_hs__conb_1
Xsky130_fd_sc_hs__conb_1_43 DVSS: DVDD: DVDD: DVSS: prbs_generator_syn_5/eqn[5] prbs_generator_syn_5/eqn[1]
+ sky130_fd_sc_hs__conb_1_43/a_165_290# sky130_fd_sc_hs__conb_1_43/a_21_290# sky130_fd_sc_hs__conb_1
Xsky130_fd_sc_hs__conb_1_54 DVSS: DVDD: DVDD: DVSS: prbs_generator_syn_9/eqn[30] sky130_fd_sc_hs__conb_1_55/HI
+ sky130_fd_sc_hs__conb_1_55/a_165_290# sky130_fd_sc_hs__conb_1_55/a_21_290# sky130_fd_sc_hs__conb_1
Xsky130_fd_sc_hs__conb_1_65 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__conb_1_65/LO
+ sky130_fd_sc_hs__conb_1_65/HI sky130_fd_sc_hs__conb_1_65/a_165_290# sky130_fd_sc_hs__conb_1_65/a_21_290#
+ sky130_fd_sc_hs__conb_1
Xsky130_fd_sc_hs__conb_1_76 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__conb_1_77/LO
+ sky130_fd_sc_hs__conb_1_77/HI sky130_fd_sc_hs__conb_1_77/a_165_290# sky130_fd_sc_hs__conb_1_77/a_21_290#
+ sky130_fd_sc_hs__conb_1
Xsky130_fd_sc_hs__conb_1_87 DVSS: DVDD: DVDD: DVSS: prbs_generator_syn_11/eqn[2] prbs_generator_syn_11/eqn[1]
+ sky130_fd_sc_hs__conb_1_87/a_165_290# sky130_fd_sc_hs__conb_1_87/a_21_290# sky130_fd_sc_hs__conb_1
Xsky130_fd_sc_hs__conb_1_98 DVSS: DVDD: DVDD: DVSS: prbs_generator_syn_13/eqn[9] sky130_fd_sc_hs__conb_1_99/HI
+ sky130_fd_sc_hs__conb_1_99/a_165_290# sky130_fd_sc_hs__conb_1_99/a_21_290# sky130_fd_sc_hs__conb_1
Xsky130_fd_sc_hs__inv_4_50 DVSS: DVDD: DVDD: DVSS: osc_core_1/pi3_r[2] osc_core_1/pi3_l[2]
+ sky130_fd_sc_hs__inv_4
Xsky130_fd_sc_hs__inv_4_61 DVSS: DVDD: DVDD: DVSS: hr_16t4_mux_top_3/din[14] prbs_generator_syn_17/out
+ sky130_fd_sc_hs__inv_4
Xsky130_fd_sc_hs__inv_4_72 DVSS: DVDD: DVDD: DVSS: osc_core_1/pi5_r[2] osc_core_1/pi5_l[2]
+ sky130_fd_sc_hs__inv_4
Xsky130_fd_sc_hs__inv_4_83 DVSS: DVDD: DVDD: DVSS: hr_16t4_mux_top_3/din[6] hr_16t4_mux_top_1/din[6]
+ sky130_fd_sc_hs__inv_4
Xsky130_fd_sc_hs__dlrtp_1_12 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__dlrtp_1_13/Q
+ sky130_fd_sc_hs__dlrtp_1_9/GATE sky130_fd_sc_hs__conb_1_117/HI sky130_fd_sc_hs__buf_2_109/X
+ sky130_fd_sc_hs__dlrtp_1_13/a_216_424# sky130_fd_sc_hs__dlrtp_1_13/a_759_508# sky130_fd_sc_hs__dlrtp_1_13/a_565_74#
+ sky130_fd_sc_hs__dlrtp_1_13/a_27_424# sky130_fd_sc_hs__dlrtp_1_13/a_1045_74# sky130_fd_sc_hs__dlrtp_1_13/a_643_74#
+ sky130_fd_sc_hs__dlrtp_1_13/a_817_48# sky130_fd_sc_hs__dlrtp_1_13/a_568_392# sky130_fd_sc_hs__dlrtp_1_13/a_363_74#
+ sky130_fd_sc_hs__dlrtp_1_13/a_769_74# sky130_fd_sc_hs__dlrtp_1
Xsky130_fd_sc_hs__dlrtp_1_23 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__dlrtp_1_25/Q
+ sky130_fd_sc_hs__clkbuf_2_3/X sky130_fd_sc_hs__conb_1_119/HI sky130_fd_sc_hs__dlrtp_1_25/D
+ sky130_fd_sc_hs__dlrtp_1_25/a_216_424# sky130_fd_sc_hs__dlrtp_1_25/a_759_508# sky130_fd_sc_hs__dlrtp_1_25/a_565_74#
+ sky130_fd_sc_hs__dlrtp_1_25/a_27_424# sky130_fd_sc_hs__dlrtp_1_25/a_1045_74# sky130_fd_sc_hs__dlrtp_1_25/a_643_74#
+ sky130_fd_sc_hs__dlrtp_1_25/a_817_48# sky130_fd_sc_hs__dlrtp_1_25/a_568_392# sky130_fd_sc_hs__dlrtp_1_25/a_363_74#
+ sky130_fd_sc_hs__dlrtp_1_25/a_769_74# sky130_fd_sc_hs__dlrtp_1
Xsky130_fd_sc_hs__dlrtp_1_34 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__dlrtp_1_35/Q
+ sky130_fd_sc_hs__clkbuf_2_3/A sky130_fd_sc_hs__conb_1_121/HI sky130_fd_sc_hs__dlrtp_1_35/D
+ sky130_fd_sc_hs__dlrtp_1_35/a_216_424# sky130_fd_sc_hs__dlrtp_1_35/a_759_508# sky130_fd_sc_hs__dlrtp_1_35/a_565_74#
+ sky130_fd_sc_hs__dlrtp_1_35/a_27_424# sky130_fd_sc_hs__dlrtp_1_35/a_1045_74# sky130_fd_sc_hs__dlrtp_1_35/a_643_74#
+ sky130_fd_sc_hs__dlrtp_1_35/a_817_48# sky130_fd_sc_hs__dlrtp_1_35/a_568_392# sky130_fd_sc_hs__dlrtp_1_35/a_363_74#
+ sky130_fd_sc_hs__dlrtp_1_35/a_769_74# sky130_fd_sc_hs__dlrtp_1
Xsky130_fd_sc_hs__dlrtp_1_45 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__dlrtp_1_45/Q
+ sky130_fd_sc_hs__clkbuf_16_53/A sky130_fd_sc_hs__conb_1_123/HI sky130_fd_sc_hs__buf_2_49/X
+ sky130_fd_sc_hs__dlrtp_1_45/a_216_424# sky130_fd_sc_hs__dlrtp_1_45/a_759_508# sky130_fd_sc_hs__dlrtp_1_45/a_565_74#
+ sky130_fd_sc_hs__dlrtp_1_45/a_27_424# sky130_fd_sc_hs__dlrtp_1_45/a_1045_74# sky130_fd_sc_hs__dlrtp_1_45/a_643_74#
+ sky130_fd_sc_hs__dlrtp_1_45/a_817_48# sky130_fd_sc_hs__dlrtp_1_45/a_568_392# sky130_fd_sc_hs__dlrtp_1_45/a_363_74#
+ sky130_fd_sc_hs__dlrtp_1_45/a_769_74# sky130_fd_sc_hs__dlrtp_1
Xsky130_fd_sc_hs__dlrtp_1_56 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__dlrtp_1_58/Q
+ sky130_fd_sc_hs__clkbuf_16_53/A sky130_fd_sc_hs__conb_1_125/HI sky130_fd_sc_hs__dlrtp_1_58/D
+ sky130_fd_sc_hs__dlrtp_1_58/a_216_424# sky130_fd_sc_hs__dlrtp_1_58/a_759_508# sky130_fd_sc_hs__dlrtp_1_58/a_565_74#
+ sky130_fd_sc_hs__dlrtp_1_58/a_27_424# sky130_fd_sc_hs__dlrtp_1_58/a_1045_74# sky130_fd_sc_hs__dlrtp_1_58/a_643_74#
+ sky130_fd_sc_hs__dlrtp_1_58/a_817_48# sky130_fd_sc_hs__dlrtp_1_58/a_568_392# sky130_fd_sc_hs__dlrtp_1_58/a_363_74#
+ sky130_fd_sc_hs__dlrtp_1_58/a_769_74# sky130_fd_sc_hs__dlrtp_1
Xsky130_fd_sc_hs__dlrtp_1_67 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__dlrtp_1_67/Q
+ sky130_fd_sc_hs__clkbuf_16_53/A sky130_fd_sc_hs__conb_1_129/HI sky130_fd_sc_hs__buf_2_57/X
+ sky130_fd_sc_hs__dlrtp_1_67/a_216_424# sky130_fd_sc_hs__dlrtp_1_67/a_759_508# sky130_fd_sc_hs__dlrtp_1_67/a_565_74#
+ sky130_fd_sc_hs__dlrtp_1_67/a_27_424# sky130_fd_sc_hs__dlrtp_1_67/a_1045_74# sky130_fd_sc_hs__dlrtp_1_67/a_643_74#
+ sky130_fd_sc_hs__dlrtp_1_67/a_817_48# sky130_fd_sc_hs__dlrtp_1_67/a_568_392# sky130_fd_sc_hs__dlrtp_1_67/a_363_74#
+ sky130_fd_sc_hs__dlrtp_1_67/a_769_74# sky130_fd_sc_hs__dlrtp_1
Xsky130_fd_sc_hs__dlrtp_1_78 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__dlrtp_1_79/Q
+ sky130_fd_sc_hs__clkbuf_16_53/X sky130_fd_sc_hs__conb_1_129/HI sky130_fd_sc_hs__dlrtp_1_79/D
+ sky130_fd_sc_hs__dlrtp_1_79/a_216_424# sky130_fd_sc_hs__dlrtp_1_79/a_759_508# sky130_fd_sc_hs__dlrtp_1_79/a_565_74#
+ sky130_fd_sc_hs__dlrtp_1_79/a_27_424# sky130_fd_sc_hs__dlrtp_1_79/a_1045_74# sky130_fd_sc_hs__dlrtp_1_79/a_643_74#
+ sky130_fd_sc_hs__dlrtp_1_79/a_817_48# sky130_fd_sc_hs__dlrtp_1_79/a_568_392# sky130_fd_sc_hs__dlrtp_1_79/a_363_74#
+ sky130_fd_sc_hs__dlrtp_1_79/a_769_74# sky130_fd_sc_hs__dlrtp_1
Xsky130_fd_sc_hs__dlrtp_1_89 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__buf_2_71/A sky130_fd_sc_hs__clkbuf_16_53/A
+ sky130_fd_sc_hs__conb_1_137/HI sky130_fd_sc_hs__dlrtp_1_89/D sky130_fd_sc_hs__dlrtp_1_89/a_216_424#
+ sky130_fd_sc_hs__dlrtp_1_89/a_759_508# sky130_fd_sc_hs__dlrtp_1_89/a_565_74# sky130_fd_sc_hs__dlrtp_1_89/a_27_424#
+ sky130_fd_sc_hs__dlrtp_1_89/a_1045_74# sky130_fd_sc_hs__dlrtp_1_89/a_643_74# sky130_fd_sc_hs__dlrtp_1_89/a_817_48#
+ sky130_fd_sc_hs__dlrtp_1_89/a_568_392# sky130_fd_sc_hs__dlrtp_1_89/a_363_74# sky130_fd_sc_hs__dlrtp_1_89/a_769_74#
+ sky130_fd_sc_hs__dlrtp_1
Xsky130_fd_sc_hs__einvp_2_5 DVSS: DVDD: DVDD: DVSS: dout_n sky130_fd_sc_hs__buf_8_1/A
+ sky130_fd_sc_hs__dlrtp_1_7/Q sky130_fd_sc_hs__einvp_2_5/a_263_323# sky130_fd_sc_hs__einvp_2_5/a_36_74#
+ sky130_fd_sc_hs__einvp_2_5/a_27_368# sky130_fd_sc_hs__einvp_2
Xsky130_fd_sc_hs__clkbuf_2_8 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__dlrtp_1_58/D
+ sky130_fd_sc_hs__o21bai_2_3/Y sky130_fd_sc_hs__clkbuf_2_9/a_43_192# sky130_fd_sc_hs__clkbuf_2
Xsky130_fd_sc_hs__clkbuf_2_19 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__dlrtp_1_65/D
+ sky130_fd_sc_hs__o21ai_2_15/Y sky130_fd_sc_hs__clkbuf_2_19/a_43_192# sky130_fd_sc_hs__clkbuf_2
Xsky130_fd_sc_hs__einvp_8_10 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__inv_4_39/A sky130_fd_sc_hs__einvp_8_11/TE
+ osc_core_1/inj_out sky130_fd_sc_hs__einvp_8_11/a_802_323# sky130_fd_sc_hs__einvp_8_11/a_27_74#
+ sky130_fd_sc_hs__einvp_8_11/a_27_368# sky130_fd_sc_hs__einvp_8
Xsky130_fd_sc_hs__buf_2_15 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__buf_2_15/A sky130_fd_sc_hs__buf_2_15/X
+ sky130_fd_sc_hs__buf_2_15/a_21_260# sky130_fd_sc_hs__buf_2
Xsky130_fd_sc_hs__buf_2_26 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__buf_2_39/X sky130_fd_sc_hs__buf_2_29/X
+ sky130_fd_sc_hs__buf_2_29/a_21_260# sky130_fd_sc_hs__buf_2
Xsky130_fd_sc_hs__buf_2_37 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__buf_2_37/A sky130_fd_sc_hs__buf_2_37/X
+ sky130_fd_sc_hs__buf_2_37/a_21_260# sky130_fd_sc_hs__buf_2
Xsky130_fd_sc_hs__buf_2_48 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__buf_2_51/X sky130_fd_sc_hs__buf_2_49/X
+ sky130_fd_sc_hs__buf_2_49/a_21_260# sky130_fd_sc_hs__buf_2
Xsky130_fd_sc_hs__buf_2_59 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__buf_2_59/A sky130_fd_sc_hs__buf_2_59/X
+ sky130_fd_sc_hs__buf_2_59/a_21_260# sky130_fd_sc_hs__buf_2
Xsky130_fd_sc_hs__o21bai_2_17 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__o21bai_2_5/A1
+ sky130_fd_sc_hs__nand2_2_11/B sky130_fd_sc_hs__dlrtp_1_157/D sky130_fd_sc_hs__buf_2_69/A
+ sky130_fd_sc_hs__o21bai_2_17/a_27_74# sky130_fd_sc_hs__o21bai_2_17/a_225_74# sky130_fd_sc_hs__o21bai_2_17/a_507_368#
+ sky130_fd_sc_hs__o21bai_2
Xsky130_fd_sc_hs__o21bai_2_28 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__clkinv_4_5/Y
+ sky130_fd_sc_hs__buf_8_3/X sky130_fd_sc_hs__buf_2_103/X sky130_fd_sc_hs__buf_2_109/A
+ sky130_fd_sc_hs__o21bai_2_29/a_27_74# sky130_fd_sc_hs__o21bai_2_29/a_225_74# sky130_fd_sc_hs__o21bai_2_29/a_507_368#
+ sky130_fd_sc_hs__o21bai_2
Xsky130_fd_sc_hs__o21bai_2_39 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__o21ai_4_1/A1
+ sky130_fd_sc_hs__clkinv_4_5/Y sky130_fd_sc_hs__dlrtp_1_19/D sky130_fd_sc_hs__buf_2_113/A
+ sky130_fd_sc_hs__o21bai_2_39/a_27_74# sky130_fd_sc_hs__o21bai_2_39/a_225_74# sky130_fd_sc_hs__o21bai_2_39/a_507_368#
+ sky130_fd_sc_hs__o21bai_2
Xsky130_fd_sc_hs__o21bai_4_6 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__buf_2_151/A
+ sky130_fd_sc_hs__o21bai_4_7/A1 sky130_fd_sc_hs__nand2_2_3/B sky130_fd_sc_hs__dlrtp_1_55/D
+ sky130_fd_sc_hs__o21bai_4_7/a_28_368# sky130_fd_sc_hs__o21bai_4_7/a_27_74# sky130_fd_sc_hs__o21bai_4_7/a_828_48#
+ sky130_fd_sc_hs__o21bai_4
Xsky130_fd_sc_hs__conb_1_204 DVSS: DVDD: DVDD: DVSS: prbs_generator_syn_29/eqn[2]
+ prbs_generator_syn_29/eqn[1] sky130_fd_sc_hs__conb_1_205/a_165_290# sky130_fd_sc_hs__conb_1_205/a_21_290#
+ sky130_fd_sc_hs__conb_1
Xsky130_fd_sc_hs__conb_1_215 DVSS: DVDD: DVDD: DVSS: prbs_generator_syn_25/eqn[9]
+ sky130_fd_sc_hs__conb_1_215/HI sky130_fd_sc_hs__conb_1_215/a_165_290# sky130_fd_sc_hs__conb_1_215/a_21_290#
+ sky130_fd_sc_hs__conb_1
Xsky130_fd_sc_hs__conb_1_226 DVSS: DVDD: DVDD: DVSS: prbs_generator_syn_23/eqn[30]
+ sky130_fd_sc_hs__conb_1_227/HI sky130_fd_sc_hs__conb_1_227/a_165_290# sky130_fd_sc_hs__conb_1_227/a_21_290#
+ sky130_fd_sc_hs__conb_1
Xsky130_fd_sc_hs__conb_1_237 DVSS: DVDD: DVDD: DVSS: prbs_generator_syn_27/eqn[22]
+ prbs_generator_syn_27/eqn[20] sky130_fd_sc_hs__conb_1_237/a_165_290# sky130_fd_sc_hs__conb_1_237/a_21_290#
+ sky130_fd_sc_hs__conb_1
Xsky130_fd_sc_hs__conb_1_248 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__conb_1_249/LO
+ sky130_fd_sc_hs__conb_1_249/HI sky130_fd_sc_hs__conb_1_249/a_165_290# sky130_fd_sc_hs__conb_1_249/a_21_290#
+ sky130_fd_sc_hs__conb_1
Xsky130_fd_sc_hs__conb_1_259 DVSS: DVDD: DVDD: DVSS: prbs_generator_syn_31/eqn[30]
+ sky130_fd_sc_hs__conb_1_259/HI sky130_fd_sc_hs__conb_1_259/a_165_290# sky130_fd_sc_hs__conb_1_259/a_21_290#
+ sky130_fd_sc_hs__conb_1
Xsky130_fd_sc_hs__clkbuf_8_18 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__clkbuf_8_19/X
+ sky130_fd_sc_hs__clkbuf_8_19/A sky130_fd_sc_hs__clkbuf_8_19/a_125_368# sky130_fd_sc_hs__clkbuf_8
Xsky130_fd_sc_hs__clkbuf_8_29 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__clkbuf_8_29/X
+ sky130_fd_sc_hs__clkbuf_8_29/A sky130_fd_sc_hs__clkbuf_8_29/a_125_368# sky130_fd_sc_hs__clkbuf_8
Xsky130_fd_sc_hs__diode_2_0 hr_16t4_mux_top_1/din[1] DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__diode_2
Xsky130_fd_sc_hs__o21bai_2_3 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__nand2_2_5/B
+ sky130_fd_sc_hs__o21bai_2_3/A2 sky130_fd_sc_hs__buf_2_55/X sky130_fd_sc_hs__o21bai_2_3/Y
+ sky130_fd_sc_hs__o21bai_2_3/a_27_74# sky130_fd_sc_hs__o21bai_2_3/a_225_74# sky130_fd_sc_hs__o21bai_2_3/a_507_368#
+ sky130_fd_sc_hs__o21bai_2
Xsky130_fd_sc_hs__o21ai_2_30 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__inv_4_19/Y sky130_fd_sc_hs__o21ai_2_31/A2
+ sky130_fd_sc_hs__o21ai_4_1/A1 sky130_fd_sc_hs__buf_2_83/A sky130_fd_sc_hs__o21ai_2_31/a_116_368#
+ sky130_fd_sc_hs__o21ai_2_31/a_27_74# sky130_fd_sc_hs__o21ai_2
Xsky130_fd_sc_hs__o21ai_2_41 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__inv_4_23/Y sky130_fd_sc_hs__nand2_2_15/B
+ sky130_fd_sc_hs__clkinv_4_7/Y sky130_fd_sc_hs__o21ai_2_41/Y sky130_fd_sc_hs__o21ai_2_41/a_116_368#
+ sky130_fd_sc_hs__o21ai_2_41/a_27_74# sky130_fd_sc_hs__o21ai_2
Xsky130_fd_sc_hs__o21ai_2_52 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__nand2_2_27/B
+ sky130_fd_sc_hs__or2b_4_1/X sky130_fd_sc_hs__nand2_2_21/B sky130_fd_sc_hs__buf_2_137/A
+ sky130_fd_sc_hs__o21ai_2_53/a_116_368# sky130_fd_sc_hs__o21ai_2_53/a_27_74# sky130_fd_sc_hs__o21ai_2
Xsky130_fd_sc_hs__clkinv_4_11 DVSS: DVDD: DVDD: DVSS: osc_core_1/pi2_r[3] osc_core_1/pi2_l[3]
+ sky130_fd_sc_hs__clkinv_4
Xsky130_fd_sc_hs__einvn_1_0 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__inv_4_49/Y sky130_fd_sc_hs__buf_1_1/A
+ sky130_fd_sc_hs__clkinv_8_15/Y sky130_fd_sc_hs__einvn_1_1/a_281_100# sky130_fd_sc_hs__einvn_1_1/a_278_368#
+ sky130_fd_sc_hs__einvn_1_1/a_22_46# sky130_fd_sc_hs__einvn_1
Xprbs_generator_syn_13 prbs_generator_syn_19/clk prbs_generator_syn_13/rst prbs_generator_syn_13/cke
+ sky130_fd_sc_hs__conb_1_109/LO sky130_fd_sc_hs__conb_1_109/LO sky130_fd_sc_hs__conb_1_109/LO
+ sky130_fd_sc_hs__conb_1_109/LO sky130_fd_sc_hs__conb_1_109/LO sky130_fd_sc_hs__conb_1_109/LO
+ sky130_fd_sc_hs__conb_1_109/HI sky130_fd_sc_hs__conb_1_109/HI sky130_fd_sc_hs__conb_1_109/HI
+ sky130_fd_sc_hs__conb_1_109/HI sky130_fd_sc_hs__conb_1_109/HI prbs_generator_syn_13/cke
+ sky130_fd_sc_hs__conb_1_111/HI sky130_fd_sc_hs__conb_1_111/HI sky130_fd_sc_hs__conb_1_111/HI
+ sky130_fd_sc_hs__conb_1_111/HI prbs_generator_syn_15/eqn[13] sky130_fd_sc_hs__conb_1_111/HI
+ prbs_generator_syn_13/eqn[2] prbs_generator_syn_13/eqn[1] prbs_generator_syn_13/eqn[2]
+ prbs_generator_syn_13/eqn[1] prbs_generator_syn_13/eqn[2] prbs_generator_syn_13/eqn[1]
+ sky130_fd_sc_hs__conb_1_115/LO sky130_fd_sc_hs__conb_1_115/HI sky130_fd_sc_hs__conb_1_115/LO
+ sky130_fd_sc_hs__conb_1_115/LO sky130_fd_sc_hs__conb_1_115/HI sky130_fd_sc_hs__conb_1_115/HI
+ sky130_fd_sc_hs__conb_1_115/LO sky130_fd_sc_hs__conb_1_115/LO prbs_generator_syn_13/eqn[31]
+ prbs_generator_syn_13/eqn[30] prbs_generator_syn_13/eqn[30] prbs_generator_syn_13/eqn[30]
+ prbs_generator_syn_13/eqn[30] prbs_generator_syn_13/eqn[30] prbs_generator_syn_13/eqn[30]
+ prbs_generator_syn_13/eqn[30] prbs_generator_syn_13/eqn[30] prbs_generator_syn_13/eqn[22]
+ prbs_generator_syn_13/eqn[22] prbs_generator_syn_13/eqn[20] prbs_generator_syn_13/eqn[22]
+ prbs_generator_syn_13/eqn[22] prbs_generator_syn_13/eqn[22] prbs_generator_syn_13/eqn[22]
+ prbs_generator_syn_13/eqn[22] prbs_generator_syn_13/eqn[22] sky130_fd_sc_hs__conb_1_97/LO
+ sky130_fd_sc_hs__conb_1_97/LO sky130_fd_sc_hs__conb_1_97/LO prbs_generator_syn_13/eqn[9]
+ prbs_generator_syn_13/eqn[9] prbs_generator_syn_13/eqn[9] prbs_generator_syn_13/eqn[9]
+ prbs_generator_syn_13/eqn[9] prbs_generator_syn_13/eqn[9] prbs_generator_syn_13/eqn[9]
+ prbs_generator_syn_13/eqn[9] prbs_generator_syn_13/eqn[2] prbs_generator_syn_13/eqn[1]
+ prbs_generator_syn_13/eqn[2] prbs_generator_syn_19/inj_err prbs_generator_syn_13/eqn[31]
+ prbs_generator_syn_13/eqn[31] hr_16t4_mux_top_1/din[5] DVSS: DVDD: prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_1/a_293_74#
+ prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_15/X prbs_generator_syn_13/sky130_fd_sc_hs__nand2_1_35/B
+ prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_51/Y prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_9/A
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_9/CLK prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_47/a_27_74#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_37/a_1226_296# prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_3/B
+ prbs_generator_syn_13/sky130_fd_sc_hs__nor2b_1_7/a_27_112# prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_29/B
+ prbs_generator_syn_13/sky130_fd_sc_hs__sdlclkp_2_1/a_580_74# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_1/a_1141_508#
+ prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_5/Y prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_41/a_230_79#
+ prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_61/a_138_385# prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_43/a_132_392#
+ prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_3/a_222_392# prbs_generator_syn_13/sky130_fd_sc_hs__nor2b_1_9/a_27_112#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_61/a_27_74# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_35/a_206_368#
+ prbs_generator_syn_13/sky130_fd_sc_hs__nand2_2_3/Y prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_25/B
+ prbs_generator_syn_13/sky130_fd_sc_hs__nand2_1_11/a_117_74# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_67/a_651_503#
+ prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_45/X prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_39/a_696_458#
+ prbs_generator_syn_13/sky130_fd_sc_hs__sdlclkp_2_1/a_1198_74# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_45/a_1034_424#
+ prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_17/a_222_392# prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_55/a_222_392#
+ prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_53/Y prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_35/A
+ prbs_generator_syn_13/m3_13600_1651# prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_59/a_52_123#
+ prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_5/a_293_74# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_35/a_1226_296#
+ prbs_generator_syn_13/sky130_fd_sc_hs__nand2_1_51/B prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_5/a_651_503#
+ prbs_generator_syn_13/sky130_fd_sc_hs__nand2_1_21/B prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_8/a_27_74#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_15/a_27_74# prbs_generator_syn_13/sky130_fd_sc_hs__and2b_2_1/X
+ prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_13/X prbs_generator_syn_13/sky130_fd_sc_hs__nand2_2_3/a_27_74#
+ prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_50/a_138_385# prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_33/a_132_392#
+ prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_1/a_376_368# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_25/a_206_368#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_35/a_437_503# prbs_generator_syn_13/sky130_fd_sc_hs__sdlclkp_2_1/a_708_451#
+ prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_45/a_230_79# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_29/a_696_458#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_32/a_27_74# prbs_generator_syn_13/sky130_fd_sc_hs__nor2b_1_4/Y
+ prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_59/a_293_74# prbs_generator_syn_13/sky130_fd_sc_hs__nand2_1_47/a_117_74#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_73/a_735_102# prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_21/a_112_119#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_23/a_1141_508# prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_25/a_293_74#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_7/Q prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_3/a_112_119#
+ prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_35/B prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_51/X
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_53/a_1178_124# prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_23/a_132_392#
+ prbs_generator_syn_13/sky130_fd_sc_hs__nand2_1_3/B prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_15/a_206_368#
+ prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_63/a_132_392# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_55/a_27_74#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_25/a_437_503# prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_41/a_52_123#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_47/a_651_503# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_73/a_1141_508#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_19/a_696_458# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_57/a_696_458#
+ prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_7/X prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_43/a_1034_424#
+ prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_55/A prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_11/a_112_119#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_21/a_1141_508# prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_35/a_222_392#
+ prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_49/a_230_79# prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_67/Y
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_71/a_27_74# prbs_generator_syn_13/sky130_fd_sc_hs__nand2_1_33/B
+ prbs_generator_syn_13/sky130_fd_sc_hs__conb_1_1/LO prbs_generator_syn_13/sky130_fd_sc_hs__nand2_1_19/a_117_74#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_51/a_1178_124# prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_33/X
+ prbs_generator_syn_13/sky130_fd_sc_hs__nand2_1_29/B prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_41/Y
+ prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_53/a_132_392# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_45/a_206_368#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_15/a_437_503# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_37/a_651_503#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_39/a_544_485# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_53/a_735_102#
+ prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_45/a_52_123# prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_1/B
+ prbs_generator_syn_13/sky130_fd_sc_hs__nand2_2_3/B prbs_generator_syn_13/sky130_fd_sc_hs__clkbuf_16_1/A
+ prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_21/X prbs_generator_syn_13/sky130_fd_sc_hs__nand2_1_25/B
+ prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_39/a_376_368# prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_63/X
+ prbs_generator_syn_13/m3_13600_3481# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_69/a_1178_124#
+ prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_21/a_138_385# prbs_generator_syn_13/sky130_fd_sc_hs__nor2b_1_8/Y
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_19/a_1178_124# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_49/a_27_74#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_45/a_437_503# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_27/a_651_503#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_71/a_1141_508# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_65/a_651_503#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_29/a_544_485# prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_3/a_138_385#
+ prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_55/X prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_43/a_735_102#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_41/a_1034_424# prbs_generator_syn_13/sky130_fd_sc_hs__nand2_1_9/B
+ prbs_generator_syn_13/sky130_fd_sc_hs__nor2b_1_9/Y prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_59/a_1034_424#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_39/a_1141_508# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_33/a_1226_296#
+ prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_49/a_52_123# prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_47/Y
+ prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_43/Y prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_4/a_651_503#
+ prbs_generator_syn_13/sky130_fd_sc_hs__nand2_1_49/B prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_19/A
+ prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_11/a_138_385# prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_5/X
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_63/a_206_368# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_17/a_651_503#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_19/a_544_485# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_55/a_651_503#
+ prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_9/Y prbs_generator_syn_13/sky130_fd_sc_hs__nand2_1_17/B
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_57/a_544_485# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_67/a_696_458#
+ prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_35/X prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_19/a_27_74#
+ prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_45/a_222_392# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_32/a_1226_296#
+ prbs_generator_syn_13/sky130_fd_sc_hs__nand2_1_43/B prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_25/A
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_1/a_206_368# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_49/a_1226_296#
+ prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_1/a_112_119# prbs_generator_syn_13/sky130_fd_sc_hs__or2_1_1/X
+ prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_59/a_376_368# prbs_generator_syn_13/sky130_fd_sc_hs__nand2_1_19/B
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_5/a_696_458# prbs_generator_syn_13/sky130_fd_sc_hs__nor2b_1_1/Y
+ prbs_generator_syn_13/sky130_fd_sc_hs__nor2b_1_5/a_278_368# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_17/a_1178_124#
+ prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_39/X prbs_generator_syn_13/m3_13600_5433#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_63/a_437_503# prbs_generator_syn_13/sky130_fd_sc_hs__nand2_2_5/B
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_23/a_735_102# prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_53/A
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_61/a_735_102# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_57/a_1034_424#
+ prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_63/B prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_37/a_1141_508#
+ prbs_generator_syn_13/sky130_fd_sc_hs__nand2_1_47/B prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_29/X
+ prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_65/Y prbs_generator_syn_13/m3_13600_4701#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_1/a_437_503# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_67/a_1178_124#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_9/a_735_102# prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_13/a_132_392#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_15/a_1178_124# prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_15/A
+ prbs_generator_syn_13/sky130_fd_sc_hs__nand2_1_1/B prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_43/B
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_35/a_651_503# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_8/D
+ prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_29/A prbs_generator_syn_13/sky130_fd_sc_hs__nand2_1_7/B
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_13/a_735_102# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_47/a_696_458#
+ prbs_generator_syn_13/sky130_fd_sc_hs__nand2_1_31/B prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_51/a_735_102#
+ prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_59/X prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_35/a_1141_508#
+ prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_25/a_222_392# prbs_generator_syn_13/sky130_fd_sc_hs__sdlclkp_2_1/a_288_48#
+ prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_55/B prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_17/B
+ prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_43/A prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_7/A
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_65/a_1178_124# prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_59/Y
+ prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_41/X prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_21/a_230_79#
+ prbs_generator_syn_13/sky130_fd_sc_hs__nand2_1_57/a_117_74# prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_1/a_222_392#
+ prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_19/B prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_35/a_293_74#
+ prbs_generator_syn_13/sky130_fd_sc_hs__nand2_1_23/a_117_74# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_73/a_206_368#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_25/a_651_503# prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_1/a_138_385#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_37/a_696_458# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_67/a_544_485#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_43/a_27_74# prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_9/X
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_55/a_1034_424# prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_39/a_112_119#
+ prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_15/a_222_392# prbs_generator_syn_13/sky130_fd_sc_hs__conb_1_1/HI
+ prbs_generator_syn_13/sky130_fd_sc_hs__nand2_1_23/B prbs_generator_syn_13/sky130_fd_sc_hs__nand2_1_53/B
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_9/a_1178_124# prbs_generator_syn_13/sky130_fd_sc_hs__nor2b_1_4/A
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_47/a_1226_296# prbs_generator_syn_13/m3_13600_11045#
+ prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_17/X prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_29/a_376_368#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_5/a_544_485# prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_3/X
+ prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_31/a_132_392# prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_61/A
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_15/a_651_503# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_73/a_437_503#
+ prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_25/a_230_79# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_27/a_696_458#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_65/a_696_458# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_33/a_735_102#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_71/a_735_102# prbs_generator_syn_13/m3_13600_7263#
+ prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_43/a_222_392# prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_50/Y
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_8/a_1178_124# prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_53/B
+ prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_19/a_376_368# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_63/a_1178_124#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_4/a_696_458# prbs_generator_syn_13/sky130_fd_sc_hs__nor2b_1_4/a_278_368#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_13/a_1178_124# prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_61/a_132_392#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_53/a_206_368# prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_21/a_52_123#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_45/a_651_503# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_17/a_696_458#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_47/a_544_485# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_55/a_696_458#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_21/a_735_102# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_37/a_27_74#
+ prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_61/B prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_61/X
+ prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_59/a_112_119# prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_31/A
+ prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_33/a_222_392# prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_29/a_230_79#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_45/a_1226_296# prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_9/a_132_392#
+ prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_5/A prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_57/Y
+ prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_31/X prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_51/a_27_74#
+ prbs_generator_syn_13/sky130_fd_sc_hs__nor2b_1_8/a_27_112# prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_47/a_376_368#
+ prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_53/a_293_74# prbs_generator_syn_13/sky130_fd_sc_hs__nand2_1_43/a_117_74#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_8/a_735_102# prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_21/a_293_74#
+ prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_39/a_138_385# prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_63/Y
+ prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_51/a_132_392# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_43/a_206_368#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_53/a_437_503# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_37/a_544_485#
+ prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_57/X prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_53/a_1034_424#
+ prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_25/a_52_123# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_33/a_1141_508#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_63/Q prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_23/a_222_392#
+ prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_63/a_222_392# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_7/a_1178_124#
+ prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_53/X prbs_generator_syn_13/sky130_fd_sc_hs__nand2_2_5/Y
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_61/a_1178_124# prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_1/a_230_79#
+ prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_43/a_230_79# prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_11/a_230_79#
+ prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_41/a_132_392# prbs_generator_syn_13/sky130_fd_sc_hs__nand2_1_13/a_117_74#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_43/a_437_503# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_27/a_544_485#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_63/a_651_503# prbs_generator_syn_13/sky130_fd_sc_hs__nand2_1_7/a_117_74#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_35/a_696_458# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_65/a_544_485#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_51/a_1034_424# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_41/a_735_102#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_32/a_1141_508# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_49/a_1141_508#
+ prbs_generator_syn_13/sky130_fd_sc_hs__nand2_1_55/B prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_53/a_222_392#
+ prbs_generator_syn_13/sky130_fd_sc_hs__sdlclkp_2_1/a_114_112# prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_9/a_293_74#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_43/a_1226_296# prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_29/a_52_123#
+ prbs_generator_syn_13/sky130_fd_sc_hs__nand2_1_37/B prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_1/a_651_503#
+ prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_27/a_376_368# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_4/a_544_485#
+ prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_67/a_376_368# prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_27/X
+ prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_1/X prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_59/a_138_385#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_29/a_1178_124# prbs_generator_syn_13/m3_13600_2871#
+ prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_5/a_230_79# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_23/a_206_368#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_61/a_206_368# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_17/a_544_485#
+ prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_15/a_230_79# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_25/a_696_458#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_55/a_544_485# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_32/a_735_102#
+ prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_29/a_293_74# prbs_generator_syn_13/sky130_fd_sc_hs__nand2_1_17/a_117_74#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_69/a_1034_424# prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_29/a_112_119#
+ prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_37/X prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_31/B
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_19/a_1034_424# prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_33/A
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_9/a_206_368# prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_57/a_376_368#
+ prbs_generator_syn_13/sky130_fd_sc_hs__sdlclkp_2_1/a_706_317# prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_11/B
+ prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_1/a_52_123# prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_39/B
+ prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_21/a_132_392# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_13/a_206_368#
+ prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_43/a_52_123# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_51/a_206_368#
+ prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_47/X prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_23/a_437_503#
+ prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_11/a_52_123# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_61/a_437_503#
+ prbs_generator_syn_13/sky130_fd_sc_hs__nor2b_1_7/Y prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_51/A
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_15/a_696_458# prbs_generator_syn_13/sky130_fd_sc_hs__nor2b_1_5/Y
+ prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_9/a_230_79# prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_25/X
+ prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_19/a_112_119# prbs_generator_syn_13/sky130_fd_sc_hs__nand2_1_45/B
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_5/a_1178_124# prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_19/a_230_79#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_41/a_1226_296# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_59/a_1226_296#
+ prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_63/a_230_79# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_51/Q
+ prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_7/a_132_392# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_9/a_437_503#
+ prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_46/a_376_368# prbs_generator_syn_13/sky130_fd_sc_hs__nand2_1_33/a_117_74#
+ prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_11/a_293_74# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_27/a_1178_124#
+ prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_11/a_132_392# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_13/a_437_503#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_51/a_437_503# prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_5/a_52_123#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_35/a_544_485# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_73/a_651_503#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_45/a_696_458# prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_15/a_52_123#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_47/a_1141_508# prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_47/a_112_119#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_4/a_1178_124# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_17/a_1034_424#
+ prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_23/B prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_37/a_376_368#
+ prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_15/B prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_7/Y
+ prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_29/a_138_385# prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_33/a_230_79#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_25/a_1178_124# prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_47/a_293_74#
+ prbs_generator_syn_13/sky130_fd_sc_hs__nand2_1_37/a_117_74# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_33/a_206_368#
+ prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_15/a_293_74# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_71/a_206_368#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_25/a_544_485# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_67/a_1034_424#
+ prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_13/a_222_392# prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_9/a_52_123#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_15/a_1034_424# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_57/a_1226_296#
+ prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_19/a_52_123# prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_23/X
+ prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_63/a_52_123# prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_19/a_138_385#
+ prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_9/a_376_368# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_21/a_206_368#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_33/a_437_503# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_71/a_437_503#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_53/a_651_503# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_15/a_544_485#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_63/a_696_458# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_65/a_1034_424#
+ prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_19/a_293_74# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_45/a_1141_508#
+ prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_27/a_112_119# prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_67/a_112_119#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_1/a_1178_124# prbs_generator_syn_13/sky130_fd_sc_hs__conb_1_1/a_21_290#
+ prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_63/a_293_74# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_8/a_206_368#
+ prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_17/a_376_368# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_63/a_27_74#
+ prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_21/A prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_55/a_376_368#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_1/a_696_458# prbs_generator_syn_13/sky130_fd_sc_hs__nor2b_1_1/a_278_368#
+ prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_47/a_138_385# prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_33/a_52_123#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_9/a_1034_424# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_21/a_437_503#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_1/a_27_74# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_43/a_651_503#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_1/Q prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_45/a_544_485#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_69/a_735_102# prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_57/a_112_119#
+ prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_31/a_222_392# prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_13/A
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_55/a_1226_296# prbs_generator_syn_13/sky130_fd_sc_hs__nand2_2_5/a_27_74#
+ prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_53/a_230_79# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_8/a_437_503#
+ prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_67/a_293_74# prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_33/a_293_74#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_7/a_735_102# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_23/a_1178_124#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_41/a_206_368# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_8/a_1034_424#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_63/a_1034_424# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_59/a_735_102#
+ prbs_generator_syn_13/sky130_fd_sc_hs__nand2_1_5/B prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_43/a_1141_508#
+ prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_46/a_112_119# prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_61/a_222_392#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_13/a_1034_424# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_73/a_1178_124#
+ prbs_generator_syn_13/sky130_fd_sc_hs__nand2_1_27/B prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_13/B
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_57/a_27_74# prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_57/a_230_79#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_21/a_1178_124# prbs_generator_syn_13/sky130_fd_sc_hs__nor2b_1_1/a_27_112#
+ prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_27/a_138_385# prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_23/a_230_79#
+ prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_67/a_138_385# prbs_generator_syn_13/sky130_fd_sc_hs__nand2_1_41/B
+ prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_9/a_222_392# prbs_generator_syn_13/sky130_fd_sc_hs__nand2_1_27/a_117_74#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_32/a_206_368# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_23/a_651_503#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_41/a_437_503# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_73/a_27_74#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_61/a_651_503# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_63/a_544_485#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_49/a_735_102# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_73/a_696_458#
+ prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_37/a_112_119# prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_51/a_222_392#
+ prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_43/X prbs_generator_syn_13/sky130_fd_sc_hs__nand2_2_1/B
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_9/a_651_503# prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_53/a_52_123#
+ prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_49/X prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_25/a_376_368#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_1/a_544_485# prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_65/a_376_368#
+ prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_57/a_138_385# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_27/a_27_74#
+ prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_39/a_132_392# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_7/a_1034_424#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_13/a_651_503# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_32/a_437_503#
+ prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_27/a_230_79# prbs_generator_syn_13/m3_13600_12265#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_51/a_651_503# prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_59/B
+ prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_47/A prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_61/a_1034_424#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_41/a_1141_508# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_59/a_1141_508#
+ prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_41/a_222_392# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_53/a_1226_296#
+ prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_3/A prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_71/a_1178_124#
+ prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_9/a_112_119# prbs_generator_syn_13/sky130_fd_sc_hs__nand2_1_3/a_117_74#
+ prbs_generator_syn_13/m3_13600_8483# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_39/a_1178_124#
+ prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_57/a_52_123# prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_46/a_138_385#
+ prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_23/a_52_123# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_67/a_27_74#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_53/a_696_458# prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_17/a_112_119#
+ prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_11/A prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_55/a_112_119#
+ prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_1/A prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_51/a_1226_296#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_29/a_1034_424# prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_59/A
+ prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_23/A prbs_generator_syn_13/sky130_fd_sc_hs__nand2_1_39/B
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_5/a_27_74# prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_57/a_293_74#
+ prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_37/a_138_385# prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_59/a_132_392#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_33/a_651_503# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_71/a_651_503#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_43/a_696_458# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_73/a_544_485#
+ prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_27/a_52_123# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_57/a_1141_508#
+ prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_21/a_222_392# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_35/a_27_74#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_69/a_1226_296# prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_37/B
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_19/a_1226_296# prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_35/a_376_368#
+ prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_47/a_230_79# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_37/a_1178_124#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_5/a_1034_424# prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_49/a_132_392#
+ prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_7/a_222_392# prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_27/a_293_74#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_21/a_651_503# prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_9/a_138_385#
+ prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_11/a_222_392# prbs_generator_syn_13/m3_13600_14095#
+ prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_50/A prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_27/a_1034_424#
+ prbs_generator_syn_13/sky130_fd_sc_hs__nand2_1_13/B prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_8/a_651_503#
+ prbs_generator_syn_13/m3_13600_9703# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_35/a_1178_124#
+ prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_17/a_138_385# prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_55/a_138_385#
+ prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_7/a_230_79# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_4/a_1034_424#
+ prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_7/a_376_368# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_69/a_206_368#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_23/a_696_458# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_53/a_544_485#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_39/a_735_102# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_61/a_696_458#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_55/a_1141_508# prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_25/a_112_119#
+ prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_65/a_112_119# prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_43/a_293_74#
+ prbs_generator_syn_13/sky130_fd_sc_hs__nand2_1_57/B prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_25/a_1034_424#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_7/a_206_368# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_17/a_1226_296#
+ prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_15/a_376_368# prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_53/a_376_368#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_9/a_696_458# prbs_generator_syn_13/m3_13600_431#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_45/a_27_74# prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_47/a_52_123#
+ prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_29/a_132_392# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_59/a_206_368#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_69/a_437_503# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_41/a_651_503#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_43/a_544_485# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_13/a_696_458#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_29/a_735_102# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_51/a_696_458#
+ prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_61/Y prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_67/a_1226_296#
+ prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_5/a_132_392# prbs_generator_syn_13/sky130_fd_sc_hs__and2b_2_1/a_198_48#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_7/a_437_503# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_15/a_1226_296#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_69/a_27_74# prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_46/a_293_74#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_1/a_1034_424# prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_19/a_132_392#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_49/a_206_368# prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_7/a_52_123#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_59/a_437_503# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_32/a_651_503#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_7/a_27_74# prbs_generator_syn_13/sky130_fd_sc_hs__nand2_2_1/a_27_74#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_19/a_735_102# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_57/a_735_102#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_65/a_1226_296# prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_37/A
+ prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_33/a_376_368# prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_37/a_230_79#
+ prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_25/a_138_385# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_39/a_27_74#
+ prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_65/a_138_385# prbs_generator_syn_13/sky130_fd_sc_hs__nor2b_1_9/a_278_368#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_49/a_437_503# prbs_generator_syn_13/sky130_fd_sc_hs__and2b_2_1/a_505_74#
+ prbs_generator_syn_13/sky130_fd_sc_hs__nand2_1_51/a_117_74# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_23/a_544_485#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_33/a_696_458# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_61/a_544_485#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_9/a_1226_296# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_53/a_1141_508#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_71/a_696_458# prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_35/a_112_119#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_23/a_1034_424# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_9/a_544_485#
+ prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_63/a_376_368# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_33/a_1178_124#
+ prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_5/a_376_368# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_13/a_544_485#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_73/a_1034_424# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_21/a_696_458#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_51/a_544_485# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_8/a_1226_296#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_51/a_1141_508# prbs_generator_syn_13/sky130_fd_sc_hs__nand2_1_55/a_117_74#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_21/a_1034_424# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_63/a_1226_296#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_23/a_27_74# prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_7/a_112_119#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_13/a_1226_296# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_8/a_696_458#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_32/a_1178_124# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_49/a_1178_124#
+ prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_37/a_52_123# prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_27/a_132_392#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_71/Q prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_67/a_735_102#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_69/a_1141_508# prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_15/a_112_119#
+ prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_53/a_112_119# prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_39/a_222_392#
+ prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_55/a_230_79# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_19/a_1141_508#
+ prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_37/a_293_74# prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_43/a_376_368#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_5/a_735_102# prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_35/a_138_385#
+ prbs_generator_syn_13/sky130_fd_sc_hs__sdlclkp_2_1/a_114_424# prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_57/a_132_392#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_71/a_1034_424# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_7/a_1226_296#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_33/a_544_485# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_41/a_696_458#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_71/a_544_485# prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_21/B
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_61/a_1226_296# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_39/a_1034_424#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_17/a_27_74# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_9/a_27_74#
+ prbs_generator_syn_13/sky130_fd_sc_hs__nor2b_1_5/a_27_112# prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_47/a_132_392#
+ prbs_generator_syn_13/sky130_fd_sc_hs__nor2b_1_8/a_278_368# prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_9/B
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_39/a_206_368# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_33/a_27_74#
+ prbs_generator_syn_13/sky130_fd_sc_hs__nand2_1_41/a_117_74# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_69/a_651_503#
+ prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_51/a_293_74# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_21/a_544_485#
+ prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_7/a_138_385# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_32/a_696_458#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_47/a_735_102# prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_33/a_112_119#
+ prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_59/a_222_392# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_17/a_1141_508#
+ prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_55/a_52_123# prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_3/a_293_74#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_7/a_651_503# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_29/a_1226_296#
+ prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_23/a_376_368# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_8/a_544_485#
+ prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_47/B prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_47/a_1178_124#
+ prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_15/a_138_385# prbs_generator_syn_13/sky130_fd_sc_hs__sdlclkp_2_1/a_1195_374#
+ prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_53/a_138_385# prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_37/a_132_392#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_29/a_206_368# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_39/a_437_503#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_59/a_651_503# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_37/a_735_102#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_67/a_1141_508# prbs_generator_syn_13/sky130_fd_sc_hs__and2b_2_1/a_27_74#
+ prbs_generator_syn_13/sky130_fd_sc_hs__conb_1_1/a_165_290# prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_55/a_293_74#
+ prbs_generator_syn_13/sky130_fd_sc_hs__nand2_1_45/a_117_74# prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_63/a_112_119#
+ prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_49/a_222_392# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_37/a_1034_424#
+ prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_23/a_293_74# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_15/a_1141_508#
+ prbs_generator_syn_13/sky130_fd_sc_hs__nand2_1_5/a_117_74# prbs_generator_syn_13/m3_13600_13485#
+ prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_5/a_112_119# prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_13/a_376_368#
+ prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_51/a_376_368# prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_7/a_293_74#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_19/a_206_368# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_57/a_206_368#
+ prbs_generator_syn_13/sky130_fd_sc_hs__sdlclkp_2_1/a_318_74# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_29/a_437_503#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_49/a_651_503# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_25/a_27_74#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_5/a_1226_296# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_41/a_544_485#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_27/a_735_102# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_65/a_1141_508#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_65/a_735_102# prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_3/a_230_79#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_35/a_1034_424# prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_13/a_230_79#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_41/a_27_74# prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_3/a_132_392#
+ prbs_generator_syn_13/sky130_fd_sc_hs__nand2_1_49/a_117_74# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_27/a_1226_296#
+ prbs_generator_syn_13/sky130_fd_sc_hs__nand2_1_15/a_117_74# prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_41/a_376_368#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_45/a_1178_124# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_4/a_735_102#
+ prbs_generator_syn_13/sky130_fd_sc_hs__nand2_1_9/a_117_74# prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_33/a_138_385#
+ prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_17/a_132_392# prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_55/a_132_392#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_9/a_1141_508# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_19/a_437_503#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_57/a_437_503# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_4/a_1226_296#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_32/a_544_485# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_17/a_735_102#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_55/a_735_102# prbs_generator_syn_13/m3_13600_2261#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_65/a_27_74# prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_29/a_222_392#
+ prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_43/a_112_119# prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_19/X
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_25/a_1226_296# prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_31/a_376_368#
+ prbs_generator_syn_13/sky130_fd_sc_hs__or2_1_1/a_63_368# prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_17/a_230_79#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_4/a_27_74# prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_61/a_230_79#
+ prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_63/a_138_385# prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_5/a_222_392#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_8/a_1141_508# prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_41/a_293_74#
+ prbs_generator_syn_13/sky130_fd_sc_hs__nand2_1_31/a_117_74# prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_5/a_138_385#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_63/a_1141_508# prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_19/a_222_392#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_13/a_1141_508# prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_3/a_52_123#
+ prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_13/a_52_123# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_43/a_1178_124#
+ prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_61/a_376_368# prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_35/a_132_392#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_67/a_206_368# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_1/a_1226_296#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_69/a_696_458# prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_31/a_230_79#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_35/a_735_102# prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_23/a_112_119#
+ prbs_generator_syn_13/sky130_fd_sc_hs__nand2_1_35/a_117_74# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_59/a_27_74#
+ prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_13/a_293_74# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_5/a_206_368#
+ prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_50/a_376_368# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_7/a_696_458#
+ prbs_generator_syn_13/sky130_fd_sc_hs__nor2b_1_7/a_278_368# prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_17/a_52_123#
+ prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_43/a_138_385# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_7/a_1141_508#
+ prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_61/a_52_123# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_67/a_437_503#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_61/a_1141_508# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_25/a_735_102#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_59/a_696_458# prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_13/a_112_119#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_33/a_1034_424# prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_51/a_112_119#
+ prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_35/a_230_79# prbs_generator_syn_13/m3_13600_4091#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_23/a_1226_296# prbs_generator_syn_13/sky130_fd_sc_hs__nand2_1_39/a_117_74#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_29/a_27_74# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_5/a_437_503#
+ prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_17/a_293_74# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_41/a_1178_124#
+ prbs_generator_syn_13/sky130_fd_sc_hs__or2_1_1/a_152_368# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_59/a_1178_124#
+ prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_61/a_293_74# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_47/a_206_368#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_39/a_651_503# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_49/a_696_458#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_15/a_735_102# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_32/a_1034_424#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_73/a_1226_296# prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_27/a_222_392#
+ prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_41/a_112_119# prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_31/a_52_123#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_49/a_1034_424# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_29/a_1141_508#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_21/a_1226_296# prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_39/a_230_79#
+ prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_23/a_138_385# prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_51/a_230_79#
+ prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_45/a_132_392# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_37/a_206_368#
+ prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_65/a_293_74# prbs_generator_syn_13/sky130_fd_sc_hs__nand2_1_53/a_117_74#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_47/a_437_503# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_29/a_651_503#
+ prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_31/a_293_74# prbs_generator_syn_13/sky130_fd_sc_hs__nand2_1_21/a_117_74#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_69/a_544_485# prbs_generator_syn_13/sky130_fd_sc_hs__clkbuf_16_1/a_114_74#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_45/a_735_102# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_13/a_27_74#
+ prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_31/a_112_119# prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_57/a_222_392#
+ prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_35/a_52_123# prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_21/a_376_368#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_7/a_544_485# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_57/a_1178_124#
+ prbs_generator_syn_13/m3_13600_6043# prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_13/a_138_385#
+ prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_51/a_138_385# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_5/a_1141_508#
+ prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_3/a_376_368# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_27/a_206_368#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_65/a_206_368# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_37/a_437_503#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_19/a_651_503# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_57/a_651_503#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_59/a_544_485# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_71/a_1226_296#
+ prbs_generator_syn_13/sky130_fd_sc_hs__nand2_1_25/a_117_74# prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_61/a_112_119#
+ prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_47/a_222_392# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_27/a_1141_508#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_53/a_27_74# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_4/a_206_368#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_39/a_1226_296# prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_11/a_376_368#
+ prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_39/a_52_123# prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_41/a_138_385#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_4/a_1141_508# prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_25/a_132_392#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_17/a_206_368# prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_41/A
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_55/a_206_368# prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_51/a_52_123#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_27/a_437_503# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_65/a_437_503#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_49/a_544_485# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_63/a_735_102#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_47/a_1034_424# prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_50/a_112_119#
+ prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_37/a_222_392# prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_59/a_230_79#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_25/a_1141_508# prbs_generator_syn_13/sky130_fd_sc_hs__nor2b_1_4/a_27_112#
+ prbs_generator_syn_13/sky130_fd_sc_hs__sdlclkp_2_1/a_685_81# prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_1/a_132_392#
+ prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_39/a_293_74# prbs_generator_syn_13/sky130_fd_sc_hs__nand2_1_29/a_117_74#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_4/a_437_503# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_55/a_1178_124#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_21/a_27_74# prbs_generator_syn_13/m3_13600_12875#
+ prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_50/a_293_74# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_1/a_735_102#
+ prbs_generator_syn_13/sky130_fd_sc_hs__xnor2_1_31/a_138_385# prbs_generator_syn_13/sky130_fd_sc_hs__a22o_1_15/a_132_392#
+ prbs_generator_syn_13/sky130_fd_sc_hs__nand2_1_1/a_117_74# prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_17/a_437_503#
+ prbs_generator_syn_13/sky130_fd_sc_hs__dfxtp_4_55/a_437_503# prbs_generator_syn
Xprbs_generator_syn_24 prbs_generator_syn_31/clk prbs_generator_syn_27/rst prbs_generator_syn_25/cke
+ sky130_fd_sc_hs__conb_1_249/LO sky130_fd_sc_hs__conb_1_249/HI sky130_fd_sc_hs__conb_1_249/HI
+ sky130_fd_sc_hs__conb_1_249/HI sky130_fd_sc_hs__conb_1_249/HI sky130_fd_sc_hs__conb_1_249/HI
+ sky130_fd_sc_hs__conb_1_249/HI sky130_fd_sc_hs__conb_1_249/HI sky130_fd_sc_hs__conb_1_249/HI
+ sky130_fd_sc_hs__conb_1_249/LO sky130_fd_sc_hs__conb_1_249/LO prbs_generator_syn_25/eqn[31]
+ prbs_generator_syn_25/cke prbs_generator_syn_25/eqn[31] prbs_generator_syn_25/cke
+ prbs_generator_syn_25/eqn[31] prbs_generator_syn_25/cke prbs_generator_syn_25/cke
+ sky130_fd_sc_hs__conb_1_233/HI prbs_generator_syn_27/eqn[20] prbs_generator_syn_27/eqn[20]
+ prbs_generator_syn_27/eqn[20] prbs_generator_syn_27/eqn[22] prbs_generator_syn_27/eqn[28]
+ sky130_fd_sc_hs__conb_1_251/HI sky130_fd_sc_hs__conb_1_251/HI prbs_generator_syn_27/eqn[28]
+ prbs_generator_syn_27/eqn[30] sky130_fd_sc_hs__conb_1_253/HI sky130_fd_sc_hs__conb_1_253/HI
+ sky130_fd_sc_hs__conb_1_253/HI sky130_fd_sc_hs__conb_1_253/HI prbs_generator_syn_25/eqn[31]
+ prbs_generator_syn_25/eqn[30] prbs_generator_syn_25/eqn[30] prbs_generator_syn_25/eqn[30]
+ prbs_generator_syn_25/eqn[30] prbs_generator_syn_25/eqn[30] prbs_generator_syn_25/eqn[30]
+ prbs_generator_syn_25/eqn[30] prbs_generator_syn_25/eqn[30] prbs_generator_syn_25/eqn[22]
+ prbs_generator_syn_25/eqn[22] prbs_generator_syn_25/eqn[20] prbs_generator_syn_25/eqn[22]
+ prbs_generator_syn_25/eqn[22] prbs_generator_syn_25/eqn[22] prbs_generator_syn_25/eqn[22]
+ prbs_generator_syn_25/eqn[22] prbs_generator_syn_25/eqn[22] prbs_generator_syn_25/eqn[9]
+ prbs_generator_syn_25/eqn[9] prbs_generator_syn_25/eqn[9] prbs_generator_syn_25/eqn[9]
+ prbs_generator_syn_25/eqn[9] prbs_generator_syn_25/eqn[8] prbs_generator_syn_25/eqn[8]
+ prbs_generator_syn_25/eqn[8] prbs_generator_syn_25/eqn[8] prbs_generator_syn_25/eqn[8]
+ prbs_generator_syn_25/eqn[8] prbs_generator_syn_25/eqn[8] prbs_generator_syn_25/eqn[1]
+ prbs_generator_syn_27/eqn[9] prbs_generator_syn_27/inj_err prbs_generator_syn_25/eqn[31]
+ prbs_generator_syn_25/eqn[31] hr_16t4_mux_top_1/din[0] DVSS: DVDD: prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_1/a_293_74#
+ prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_15/X prbs_generator_syn_25/sky130_fd_sc_hs__nand2_1_35/B
+ prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_51/Y prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_9/A
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_9/CLK prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_47/a_27_74#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_37/a_1226_296# prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_3/B
+ prbs_generator_syn_25/sky130_fd_sc_hs__nor2b_1_7/a_27_112# prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_29/B
+ prbs_generator_syn_25/sky130_fd_sc_hs__sdlclkp_2_1/a_580_74# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_1/a_1141_508#
+ prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_5/Y prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_41/a_230_79#
+ prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_61/a_138_385# prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_43/a_132_392#
+ prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_3/a_222_392# prbs_generator_syn_25/sky130_fd_sc_hs__nor2b_1_9/a_27_112#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_61/a_27_74# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_35/a_206_368#
+ prbs_generator_syn_25/sky130_fd_sc_hs__nand2_2_3/Y prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_25/B
+ prbs_generator_syn_25/sky130_fd_sc_hs__nand2_1_11/a_117_74# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_67/a_651_503#
+ prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_45/X prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_39/a_696_458#
+ prbs_generator_syn_25/sky130_fd_sc_hs__sdlclkp_2_1/a_1198_74# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_45/a_1034_424#
+ prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_17/a_222_392# prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_55/a_222_392#
+ prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_53/Y prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_35/A
+ prbs_generator_syn_25/m3_13600_1651# prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_59/a_52_123#
+ prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_5/a_293_74# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_35/a_1226_296#
+ prbs_generator_syn_25/sky130_fd_sc_hs__nand2_1_51/B prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_5/a_651_503#
+ prbs_generator_syn_25/sky130_fd_sc_hs__nand2_1_21/B prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_8/a_27_74#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_15/a_27_74# prbs_generator_syn_25/sky130_fd_sc_hs__and2b_2_1/X
+ prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_13/X prbs_generator_syn_25/sky130_fd_sc_hs__nand2_2_3/a_27_74#
+ prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_50/a_138_385# prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_33/a_132_392#
+ prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_1/a_376_368# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_25/a_206_368#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_35/a_437_503# prbs_generator_syn_25/sky130_fd_sc_hs__sdlclkp_2_1/a_708_451#
+ prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_45/a_230_79# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_29/a_696_458#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_32/a_27_74# prbs_generator_syn_25/sky130_fd_sc_hs__nor2b_1_4/Y
+ prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_59/a_293_74# prbs_generator_syn_25/sky130_fd_sc_hs__nand2_1_47/a_117_74#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_73/a_735_102# prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_21/a_112_119#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_23/a_1141_508# prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_25/a_293_74#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_7/Q prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_3/a_112_119#
+ prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_35/B prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_51/X
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_53/a_1178_124# prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_23/a_132_392#
+ prbs_generator_syn_25/sky130_fd_sc_hs__nand2_1_3/B prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_15/a_206_368#
+ prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_63/a_132_392# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_55/a_27_74#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_25/a_437_503# prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_41/a_52_123#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_47/a_651_503# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_73/a_1141_508#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_19/a_696_458# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_57/a_696_458#
+ prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_7/X prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_43/a_1034_424#
+ prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_55/A prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_11/a_112_119#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_21/a_1141_508# prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_35/a_222_392#
+ prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_49/a_230_79# prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_67/Y
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_71/a_27_74# prbs_generator_syn_25/sky130_fd_sc_hs__nand2_1_33/B
+ prbs_generator_syn_25/sky130_fd_sc_hs__conb_1_1/LO prbs_generator_syn_25/sky130_fd_sc_hs__nand2_1_19/a_117_74#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_51/a_1178_124# prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_33/X
+ prbs_generator_syn_25/sky130_fd_sc_hs__nand2_1_29/B prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_41/Y
+ prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_53/a_132_392# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_45/a_206_368#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_15/a_437_503# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_37/a_651_503#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_39/a_544_485# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_53/a_735_102#
+ prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_45/a_52_123# prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_1/B
+ prbs_generator_syn_25/sky130_fd_sc_hs__nand2_2_3/B prbs_generator_syn_25/sky130_fd_sc_hs__clkbuf_16_1/A
+ prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_21/X prbs_generator_syn_25/sky130_fd_sc_hs__nand2_1_25/B
+ prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_39/a_376_368# prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_63/X
+ prbs_generator_syn_25/m3_13600_3481# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_69/a_1178_124#
+ prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_21/a_138_385# prbs_generator_syn_25/sky130_fd_sc_hs__nor2b_1_8/Y
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_19/a_1178_124# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_49/a_27_74#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_45/a_437_503# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_27/a_651_503#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_71/a_1141_508# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_65/a_651_503#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_29/a_544_485# prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_3/a_138_385#
+ prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_55/X prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_43/a_735_102#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_41/a_1034_424# prbs_generator_syn_25/sky130_fd_sc_hs__nand2_1_9/B
+ prbs_generator_syn_25/sky130_fd_sc_hs__nor2b_1_9/Y prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_59/a_1034_424#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_39/a_1141_508# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_33/a_1226_296#
+ prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_49/a_52_123# prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_47/Y
+ prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_43/Y prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_4/a_651_503#
+ prbs_generator_syn_25/sky130_fd_sc_hs__nand2_1_49/B prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_19/A
+ prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_11/a_138_385# prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_5/X
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_63/a_206_368# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_17/a_651_503#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_19/a_544_485# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_55/a_651_503#
+ prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_9/Y prbs_generator_syn_25/sky130_fd_sc_hs__nand2_1_17/B
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_57/a_544_485# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_67/a_696_458#
+ prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_35/X prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_19/a_27_74#
+ prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_45/a_222_392# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_32/a_1226_296#
+ prbs_generator_syn_25/sky130_fd_sc_hs__nand2_1_43/B prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_25/A
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_1/a_206_368# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_49/a_1226_296#
+ prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_1/a_112_119# prbs_generator_syn_25/sky130_fd_sc_hs__or2_1_1/X
+ prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_59/a_376_368# prbs_generator_syn_25/sky130_fd_sc_hs__nand2_1_19/B
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_5/a_696_458# prbs_generator_syn_25/sky130_fd_sc_hs__nor2b_1_1/Y
+ prbs_generator_syn_25/sky130_fd_sc_hs__nor2b_1_5/a_278_368# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_17/a_1178_124#
+ prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_39/X prbs_generator_syn_25/m3_13600_5433#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_63/a_437_503# prbs_generator_syn_25/sky130_fd_sc_hs__nand2_2_5/B
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_23/a_735_102# prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_53/A
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_61/a_735_102# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_57/a_1034_424#
+ prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_63/B prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_37/a_1141_508#
+ prbs_generator_syn_25/sky130_fd_sc_hs__nand2_1_47/B prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_29/X
+ prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_65/Y prbs_generator_syn_25/m3_13600_4701#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_1/a_437_503# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_67/a_1178_124#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_9/a_735_102# prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_13/a_132_392#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_15/a_1178_124# prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_15/A
+ prbs_generator_syn_25/sky130_fd_sc_hs__nand2_1_1/B prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_43/B
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_35/a_651_503# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_8/D
+ prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_29/A prbs_generator_syn_25/sky130_fd_sc_hs__nand2_1_7/B
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_13/a_735_102# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_47/a_696_458#
+ prbs_generator_syn_25/sky130_fd_sc_hs__nand2_1_31/B prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_51/a_735_102#
+ prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_59/X prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_35/a_1141_508#
+ prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_25/a_222_392# prbs_generator_syn_25/sky130_fd_sc_hs__sdlclkp_2_1/a_288_48#
+ prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_55/B prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_17/B
+ prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_43/A prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_7/A
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_65/a_1178_124# prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_59/Y
+ prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_41/X prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_21/a_230_79#
+ prbs_generator_syn_25/sky130_fd_sc_hs__nand2_1_57/a_117_74# prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_1/a_222_392#
+ prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_19/B prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_35/a_293_74#
+ prbs_generator_syn_25/sky130_fd_sc_hs__nand2_1_23/a_117_74# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_73/a_206_368#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_25/a_651_503# prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_1/a_138_385#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_37/a_696_458# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_67/a_544_485#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_43/a_27_74# prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_9/X
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_55/a_1034_424# prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_39/a_112_119#
+ prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_15/a_222_392# prbs_generator_syn_25/sky130_fd_sc_hs__conb_1_1/HI
+ prbs_generator_syn_25/sky130_fd_sc_hs__nand2_1_23/B prbs_generator_syn_25/sky130_fd_sc_hs__nand2_1_53/B
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_9/a_1178_124# prbs_generator_syn_25/sky130_fd_sc_hs__nor2b_1_4/A
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_47/a_1226_296# prbs_generator_syn_25/m3_13600_11045#
+ prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_17/X prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_29/a_376_368#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_5/a_544_485# prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_3/X
+ prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_31/a_132_392# prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_61/A
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_15/a_651_503# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_73/a_437_503#
+ prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_25/a_230_79# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_27/a_696_458#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_65/a_696_458# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_33/a_735_102#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_71/a_735_102# prbs_generator_syn_25/m3_13600_7263#
+ prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_43/a_222_392# prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_50/Y
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_8/a_1178_124# prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_53/B
+ prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_19/a_376_368# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_63/a_1178_124#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_4/a_696_458# prbs_generator_syn_25/sky130_fd_sc_hs__nor2b_1_4/a_278_368#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_13/a_1178_124# prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_61/a_132_392#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_53/a_206_368# prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_21/a_52_123#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_45/a_651_503# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_17/a_696_458#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_47/a_544_485# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_55/a_696_458#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_21/a_735_102# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_37/a_27_74#
+ prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_61/B prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_61/X
+ prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_59/a_112_119# prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_31/A
+ prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_33/a_222_392# prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_29/a_230_79#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_45/a_1226_296# prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_9/a_132_392#
+ prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_5/A prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_57/Y
+ prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_31/X prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_51/a_27_74#
+ prbs_generator_syn_25/sky130_fd_sc_hs__nor2b_1_8/a_27_112# prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_47/a_376_368#
+ prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_53/a_293_74# prbs_generator_syn_25/sky130_fd_sc_hs__nand2_1_43/a_117_74#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_8/a_735_102# prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_21/a_293_74#
+ prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_39/a_138_385# prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_63/Y
+ prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_51/a_132_392# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_43/a_206_368#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_53/a_437_503# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_37/a_544_485#
+ prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_57/X prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_53/a_1034_424#
+ prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_25/a_52_123# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_33/a_1141_508#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_63/Q prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_23/a_222_392#
+ prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_63/a_222_392# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_7/a_1178_124#
+ prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_53/X prbs_generator_syn_25/sky130_fd_sc_hs__nand2_2_5/Y
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_61/a_1178_124# prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_1/a_230_79#
+ prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_43/a_230_79# prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_11/a_230_79#
+ prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_41/a_132_392# prbs_generator_syn_25/sky130_fd_sc_hs__nand2_1_13/a_117_74#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_43/a_437_503# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_27/a_544_485#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_63/a_651_503# prbs_generator_syn_25/sky130_fd_sc_hs__nand2_1_7/a_117_74#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_35/a_696_458# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_65/a_544_485#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_51/a_1034_424# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_41/a_735_102#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_32/a_1141_508# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_49/a_1141_508#
+ prbs_generator_syn_25/sky130_fd_sc_hs__nand2_1_55/B prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_53/a_222_392#
+ prbs_generator_syn_25/sky130_fd_sc_hs__sdlclkp_2_1/a_114_112# prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_9/a_293_74#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_43/a_1226_296# prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_29/a_52_123#
+ prbs_generator_syn_25/sky130_fd_sc_hs__nand2_1_37/B prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_1/a_651_503#
+ prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_27/a_376_368# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_4/a_544_485#
+ prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_67/a_376_368# prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_27/X
+ prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_1/X prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_59/a_138_385#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_29/a_1178_124# prbs_generator_syn_25/m3_13600_2871#
+ prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_5/a_230_79# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_23/a_206_368#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_61/a_206_368# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_17/a_544_485#
+ prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_15/a_230_79# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_25/a_696_458#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_55/a_544_485# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_32/a_735_102#
+ prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_29/a_293_74# prbs_generator_syn_25/sky130_fd_sc_hs__nand2_1_17/a_117_74#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_69/a_1034_424# prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_29/a_112_119#
+ prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_37/X prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_31/B
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_19/a_1034_424# prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_33/A
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_9/a_206_368# prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_57/a_376_368#
+ prbs_generator_syn_25/sky130_fd_sc_hs__sdlclkp_2_1/a_706_317# prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_11/B
+ prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_1/a_52_123# prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_39/B
+ prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_21/a_132_392# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_13/a_206_368#
+ prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_43/a_52_123# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_51/a_206_368#
+ prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_47/X prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_23/a_437_503#
+ prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_11/a_52_123# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_61/a_437_503#
+ prbs_generator_syn_25/sky130_fd_sc_hs__nor2b_1_7/Y prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_51/A
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_15/a_696_458# prbs_generator_syn_25/sky130_fd_sc_hs__nor2b_1_5/Y
+ prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_9/a_230_79# prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_25/X
+ prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_19/a_112_119# prbs_generator_syn_25/sky130_fd_sc_hs__nand2_1_45/B
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_5/a_1178_124# prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_19/a_230_79#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_41/a_1226_296# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_59/a_1226_296#
+ prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_63/a_230_79# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_51/Q
+ prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_7/a_132_392# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_9/a_437_503#
+ prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_46/a_376_368# prbs_generator_syn_25/sky130_fd_sc_hs__nand2_1_33/a_117_74#
+ prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_11/a_293_74# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_27/a_1178_124#
+ prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_11/a_132_392# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_13/a_437_503#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_51/a_437_503# prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_5/a_52_123#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_35/a_544_485# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_73/a_651_503#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_45/a_696_458# prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_15/a_52_123#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_47/a_1141_508# prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_47/a_112_119#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_4/a_1178_124# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_17/a_1034_424#
+ prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_23/B prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_37/a_376_368#
+ prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_15/B prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_7/Y
+ prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_29/a_138_385# prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_33/a_230_79#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_25/a_1178_124# prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_47/a_293_74#
+ prbs_generator_syn_25/sky130_fd_sc_hs__nand2_1_37/a_117_74# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_33/a_206_368#
+ prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_15/a_293_74# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_71/a_206_368#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_25/a_544_485# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_67/a_1034_424#
+ prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_13/a_222_392# prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_9/a_52_123#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_15/a_1034_424# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_57/a_1226_296#
+ prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_19/a_52_123# prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_23/X
+ prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_63/a_52_123# prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_19/a_138_385#
+ prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_9/a_376_368# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_21/a_206_368#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_33/a_437_503# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_71/a_437_503#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_53/a_651_503# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_15/a_544_485#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_63/a_696_458# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_65/a_1034_424#
+ prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_19/a_293_74# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_45/a_1141_508#
+ prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_27/a_112_119# prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_67/a_112_119#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_1/a_1178_124# prbs_generator_syn_25/sky130_fd_sc_hs__conb_1_1/a_21_290#
+ prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_63/a_293_74# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_8/a_206_368#
+ prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_17/a_376_368# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_63/a_27_74#
+ prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_21/A prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_55/a_376_368#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_1/a_696_458# prbs_generator_syn_25/sky130_fd_sc_hs__nor2b_1_1/a_278_368#
+ prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_47/a_138_385# prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_33/a_52_123#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_9/a_1034_424# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_21/a_437_503#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_1/a_27_74# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_43/a_651_503#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_1/Q prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_45/a_544_485#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_69/a_735_102# prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_57/a_112_119#
+ prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_31/a_222_392# prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_13/A
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_55/a_1226_296# prbs_generator_syn_25/sky130_fd_sc_hs__nand2_2_5/a_27_74#
+ prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_53/a_230_79# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_8/a_437_503#
+ prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_67/a_293_74# prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_33/a_293_74#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_7/a_735_102# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_23/a_1178_124#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_41/a_206_368# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_8/a_1034_424#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_63/a_1034_424# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_59/a_735_102#
+ prbs_generator_syn_25/sky130_fd_sc_hs__nand2_1_5/B prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_43/a_1141_508#
+ prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_46/a_112_119# prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_61/a_222_392#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_13/a_1034_424# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_73/a_1178_124#
+ prbs_generator_syn_25/sky130_fd_sc_hs__nand2_1_27/B prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_13/B
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_57/a_27_74# prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_57/a_230_79#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_21/a_1178_124# prbs_generator_syn_25/sky130_fd_sc_hs__nor2b_1_1/a_27_112#
+ prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_27/a_138_385# prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_23/a_230_79#
+ prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_67/a_138_385# prbs_generator_syn_25/sky130_fd_sc_hs__nand2_1_41/B
+ prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_9/a_222_392# prbs_generator_syn_25/sky130_fd_sc_hs__nand2_1_27/a_117_74#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_32/a_206_368# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_23/a_651_503#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_41/a_437_503# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_73/a_27_74#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_61/a_651_503# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_63/a_544_485#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_49/a_735_102# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_73/a_696_458#
+ prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_37/a_112_119# prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_51/a_222_392#
+ prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_43/X prbs_generator_syn_25/sky130_fd_sc_hs__nand2_2_1/B
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_9/a_651_503# prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_53/a_52_123#
+ prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_49/X prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_25/a_376_368#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_1/a_544_485# prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_65/a_376_368#
+ prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_57/a_138_385# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_27/a_27_74#
+ prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_39/a_132_392# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_7/a_1034_424#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_13/a_651_503# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_32/a_437_503#
+ prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_27/a_230_79# prbs_generator_syn_25/m3_13600_12265#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_51/a_651_503# prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_59/B
+ prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_47/A prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_61/a_1034_424#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_41/a_1141_508# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_59/a_1141_508#
+ prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_41/a_222_392# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_53/a_1226_296#
+ prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_3/A prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_71/a_1178_124#
+ prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_9/a_112_119# prbs_generator_syn_25/sky130_fd_sc_hs__nand2_1_3/a_117_74#
+ prbs_generator_syn_25/m3_13600_8483# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_39/a_1178_124#
+ prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_57/a_52_123# prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_46/a_138_385#
+ prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_23/a_52_123# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_67/a_27_74#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_53/a_696_458# prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_17/a_112_119#
+ prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_11/A prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_55/a_112_119#
+ prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_1/A prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_51/a_1226_296#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_29/a_1034_424# prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_59/A
+ prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_23/A prbs_generator_syn_25/sky130_fd_sc_hs__nand2_1_39/B
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_5/a_27_74# prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_57/a_293_74#
+ prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_37/a_138_385# prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_59/a_132_392#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_33/a_651_503# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_71/a_651_503#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_43/a_696_458# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_73/a_544_485#
+ prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_27/a_52_123# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_57/a_1141_508#
+ prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_21/a_222_392# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_35/a_27_74#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_69/a_1226_296# prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_37/B
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_19/a_1226_296# prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_35/a_376_368#
+ prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_47/a_230_79# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_37/a_1178_124#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_5/a_1034_424# prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_49/a_132_392#
+ prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_7/a_222_392# prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_27/a_293_74#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_21/a_651_503# prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_9/a_138_385#
+ prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_11/a_222_392# prbs_generator_syn_25/m3_13600_14095#
+ prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_50/A prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_27/a_1034_424#
+ prbs_generator_syn_25/sky130_fd_sc_hs__nand2_1_13/B prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_8/a_651_503#
+ prbs_generator_syn_25/m3_13600_9703# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_35/a_1178_124#
+ prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_17/a_138_385# prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_55/a_138_385#
+ prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_7/a_230_79# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_4/a_1034_424#
+ prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_7/a_376_368# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_69/a_206_368#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_23/a_696_458# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_53/a_544_485#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_39/a_735_102# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_61/a_696_458#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_55/a_1141_508# prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_25/a_112_119#
+ prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_65/a_112_119# prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_43/a_293_74#
+ prbs_generator_syn_25/sky130_fd_sc_hs__nand2_1_57/B prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_25/a_1034_424#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_7/a_206_368# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_17/a_1226_296#
+ prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_15/a_376_368# prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_53/a_376_368#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_9/a_696_458# prbs_generator_syn_25/m3_13600_431#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_45/a_27_74# prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_47/a_52_123#
+ prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_29/a_132_392# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_59/a_206_368#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_69/a_437_503# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_41/a_651_503#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_43/a_544_485# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_13/a_696_458#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_29/a_735_102# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_51/a_696_458#
+ prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_61/Y prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_67/a_1226_296#
+ prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_5/a_132_392# prbs_generator_syn_25/sky130_fd_sc_hs__and2b_2_1/a_198_48#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_7/a_437_503# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_15/a_1226_296#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_69/a_27_74# prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_46/a_293_74#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_1/a_1034_424# prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_19/a_132_392#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_49/a_206_368# prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_7/a_52_123#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_59/a_437_503# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_32/a_651_503#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_7/a_27_74# prbs_generator_syn_25/sky130_fd_sc_hs__nand2_2_1/a_27_74#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_19/a_735_102# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_57/a_735_102#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_65/a_1226_296# prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_37/A
+ prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_33/a_376_368# prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_37/a_230_79#
+ prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_25/a_138_385# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_39/a_27_74#
+ prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_65/a_138_385# prbs_generator_syn_25/sky130_fd_sc_hs__nor2b_1_9/a_278_368#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_49/a_437_503# prbs_generator_syn_25/sky130_fd_sc_hs__and2b_2_1/a_505_74#
+ prbs_generator_syn_25/sky130_fd_sc_hs__nand2_1_51/a_117_74# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_23/a_544_485#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_33/a_696_458# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_61/a_544_485#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_9/a_1226_296# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_53/a_1141_508#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_71/a_696_458# prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_35/a_112_119#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_23/a_1034_424# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_9/a_544_485#
+ prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_63/a_376_368# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_33/a_1178_124#
+ prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_5/a_376_368# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_13/a_544_485#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_73/a_1034_424# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_21/a_696_458#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_51/a_544_485# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_8/a_1226_296#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_51/a_1141_508# prbs_generator_syn_25/sky130_fd_sc_hs__nand2_1_55/a_117_74#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_21/a_1034_424# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_63/a_1226_296#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_23/a_27_74# prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_7/a_112_119#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_13/a_1226_296# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_8/a_696_458#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_32/a_1178_124# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_49/a_1178_124#
+ prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_37/a_52_123# prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_27/a_132_392#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_71/Q prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_67/a_735_102#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_69/a_1141_508# prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_15/a_112_119#
+ prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_53/a_112_119# prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_39/a_222_392#
+ prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_55/a_230_79# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_19/a_1141_508#
+ prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_37/a_293_74# prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_43/a_376_368#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_5/a_735_102# prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_35/a_138_385#
+ prbs_generator_syn_25/sky130_fd_sc_hs__sdlclkp_2_1/a_114_424# prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_57/a_132_392#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_71/a_1034_424# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_7/a_1226_296#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_33/a_544_485# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_41/a_696_458#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_71/a_544_485# prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_21/B
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_61/a_1226_296# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_39/a_1034_424#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_17/a_27_74# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_9/a_27_74#
+ prbs_generator_syn_25/sky130_fd_sc_hs__nor2b_1_5/a_27_112# prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_47/a_132_392#
+ prbs_generator_syn_25/sky130_fd_sc_hs__nor2b_1_8/a_278_368# prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_9/B
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_39/a_206_368# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_33/a_27_74#
+ prbs_generator_syn_25/sky130_fd_sc_hs__nand2_1_41/a_117_74# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_69/a_651_503#
+ prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_51/a_293_74# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_21/a_544_485#
+ prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_7/a_138_385# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_32/a_696_458#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_47/a_735_102# prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_33/a_112_119#
+ prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_59/a_222_392# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_17/a_1141_508#
+ prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_55/a_52_123# prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_3/a_293_74#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_7/a_651_503# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_29/a_1226_296#
+ prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_23/a_376_368# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_8/a_544_485#
+ prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_47/B prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_47/a_1178_124#
+ prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_15/a_138_385# prbs_generator_syn_25/sky130_fd_sc_hs__sdlclkp_2_1/a_1195_374#
+ prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_53/a_138_385# prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_37/a_132_392#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_29/a_206_368# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_39/a_437_503#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_59/a_651_503# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_37/a_735_102#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_67/a_1141_508# prbs_generator_syn_25/sky130_fd_sc_hs__and2b_2_1/a_27_74#
+ prbs_generator_syn_25/sky130_fd_sc_hs__conb_1_1/a_165_290# prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_55/a_293_74#
+ prbs_generator_syn_25/sky130_fd_sc_hs__nand2_1_45/a_117_74# prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_63/a_112_119#
+ prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_49/a_222_392# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_37/a_1034_424#
+ prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_23/a_293_74# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_15/a_1141_508#
+ prbs_generator_syn_25/sky130_fd_sc_hs__nand2_1_5/a_117_74# prbs_generator_syn_25/m3_13600_13485#
+ prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_5/a_112_119# prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_13/a_376_368#
+ prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_51/a_376_368# prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_7/a_293_74#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_19/a_206_368# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_57/a_206_368#
+ prbs_generator_syn_25/sky130_fd_sc_hs__sdlclkp_2_1/a_318_74# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_29/a_437_503#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_49/a_651_503# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_25/a_27_74#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_5/a_1226_296# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_41/a_544_485#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_27/a_735_102# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_65/a_1141_508#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_65/a_735_102# prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_3/a_230_79#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_35/a_1034_424# prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_13/a_230_79#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_41/a_27_74# prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_3/a_132_392#
+ prbs_generator_syn_25/sky130_fd_sc_hs__nand2_1_49/a_117_74# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_27/a_1226_296#
+ prbs_generator_syn_25/sky130_fd_sc_hs__nand2_1_15/a_117_74# prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_41/a_376_368#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_45/a_1178_124# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_4/a_735_102#
+ prbs_generator_syn_25/sky130_fd_sc_hs__nand2_1_9/a_117_74# prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_33/a_138_385#
+ prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_17/a_132_392# prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_55/a_132_392#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_9/a_1141_508# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_19/a_437_503#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_57/a_437_503# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_4/a_1226_296#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_32/a_544_485# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_17/a_735_102#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_55/a_735_102# prbs_generator_syn_25/m3_13600_2261#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_65/a_27_74# prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_29/a_222_392#
+ prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_43/a_112_119# prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_19/X
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_25/a_1226_296# prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_31/a_376_368#
+ prbs_generator_syn_25/sky130_fd_sc_hs__or2_1_1/a_63_368# prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_17/a_230_79#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_4/a_27_74# prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_61/a_230_79#
+ prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_63/a_138_385# prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_5/a_222_392#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_8/a_1141_508# prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_41/a_293_74#
+ prbs_generator_syn_25/sky130_fd_sc_hs__nand2_1_31/a_117_74# prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_5/a_138_385#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_63/a_1141_508# prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_19/a_222_392#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_13/a_1141_508# prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_3/a_52_123#
+ prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_13/a_52_123# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_43/a_1178_124#
+ prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_61/a_376_368# prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_35/a_132_392#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_67/a_206_368# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_1/a_1226_296#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_69/a_696_458# prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_31/a_230_79#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_35/a_735_102# prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_23/a_112_119#
+ prbs_generator_syn_25/sky130_fd_sc_hs__nand2_1_35/a_117_74# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_59/a_27_74#
+ prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_13/a_293_74# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_5/a_206_368#
+ prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_50/a_376_368# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_7/a_696_458#
+ prbs_generator_syn_25/sky130_fd_sc_hs__nor2b_1_7/a_278_368# prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_17/a_52_123#
+ prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_43/a_138_385# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_7/a_1141_508#
+ prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_61/a_52_123# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_67/a_437_503#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_61/a_1141_508# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_25/a_735_102#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_59/a_696_458# prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_13/a_112_119#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_33/a_1034_424# prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_51/a_112_119#
+ prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_35/a_230_79# prbs_generator_syn_25/m3_13600_4091#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_23/a_1226_296# prbs_generator_syn_25/sky130_fd_sc_hs__nand2_1_39/a_117_74#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_29/a_27_74# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_5/a_437_503#
+ prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_17/a_293_74# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_41/a_1178_124#
+ prbs_generator_syn_25/sky130_fd_sc_hs__or2_1_1/a_152_368# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_59/a_1178_124#
+ prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_61/a_293_74# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_47/a_206_368#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_39/a_651_503# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_49/a_696_458#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_15/a_735_102# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_32/a_1034_424#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_73/a_1226_296# prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_27/a_222_392#
+ prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_41/a_112_119# prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_31/a_52_123#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_49/a_1034_424# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_29/a_1141_508#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_21/a_1226_296# prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_39/a_230_79#
+ prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_23/a_138_385# prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_51/a_230_79#
+ prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_45/a_132_392# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_37/a_206_368#
+ prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_65/a_293_74# prbs_generator_syn_25/sky130_fd_sc_hs__nand2_1_53/a_117_74#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_47/a_437_503# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_29/a_651_503#
+ prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_31/a_293_74# prbs_generator_syn_25/sky130_fd_sc_hs__nand2_1_21/a_117_74#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_69/a_544_485# prbs_generator_syn_25/sky130_fd_sc_hs__clkbuf_16_1/a_114_74#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_45/a_735_102# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_13/a_27_74#
+ prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_31/a_112_119# prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_57/a_222_392#
+ prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_35/a_52_123# prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_21/a_376_368#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_7/a_544_485# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_57/a_1178_124#
+ prbs_generator_syn_25/m3_13600_6043# prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_13/a_138_385#
+ prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_51/a_138_385# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_5/a_1141_508#
+ prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_3/a_376_368# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_27/a_206_368#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_65/a_206_368# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_37/a_437_503#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_19/a_651_503# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_57/a_651_503#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_59/a_544_485# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_71/a_1226_296#
+ prbs_generator_syn_25/sky130_fd_sc_hs__nand2_1_25/a_117_74# prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_61/a_112_119#
+ prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_47/a_222_392# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_27/a_1141_508#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_53/a_27_74# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_4/a_206_368#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_39/a_1226_296# prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_11/a_376_368#
+ prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_39/a_52_123# prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_41/a_138_385#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_4/a_1141_508# prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_25/a_132_392#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_17/a_206_368# prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_41/A
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_55/a_206_368# prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_51/a_52_123#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_27/a_437_503# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_65/a_437_503#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_49/a_544_485# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_63/a_735_102#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_47/a_1034_424# prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_50/a_112_119#
+ prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_37/a_222_392# prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_59/a_230_79#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_25/a_1141_508# prbs_generator_syn_25/sky130_fd_sc_hs__nor2b_1_4/a_27_112#
+ prbs_generator_syn_25/sky130_fd_sc_hs__sdlclkp_2_1/a_685_81# prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_1/a_132_392#
+ prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_39/a_293_74# prbs_generator_syn_25/sky130_fd_sc_hs__nand2_1_29/a_117_74#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_4/a_437_503# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_55/a_1178_124#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_21/a_27_74# prbs_generator_syn_25/m3_13600_12875#
+ prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_50/a_293_74# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_1/a_735_102#
+ prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_31/a_138_385# prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_15/a_132_392#
+ prbs_generator_syn_25/sky130_fd_sc_hs__nand2_1_1/a_117_74# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_17/a_437_503#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_55/a_437_503# prbs_generator_syn
Xsky130_fd_sc_hs__conb_1_4 DVSS: DVDD: DVDD: DVSS: prbs_generator_syn_1/eqn[8] prbs_generator_syn_1/eqn[1]
+ sky130_fd_sc_hs__conb_1_5/a_165_290# sky130_fd_sc_hs__conb_1_5/a_21_290# sky130_fd_sc_hs__conb_1
Xsky130_fd_sc_hs__buf_2_100 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__buf_2_91/X sky130_fd_sc_hs__buf_2_101/X
+ sky130_fd_sc_hs__buf_2_101/a_21_260# sky130_fd_sc_hs__buf_2
Xsky130_fd_sc_hs__buf_2_111 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__buf_2_111/A sky130_fd_sc_hs__buf_2_111/X
+ sky130_fd_sc_hs__buf_2_111/a_21_260# sky130_fd_sc_hs__buf_2
Xsky130_fd_sc_hs__buf_2_122 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__buf_2_123/A sky130_fd_sc_hs__buf_2_123/X
+ sky130_fd_sc_hs__buf_2_123/a_21_260# sky130_fd_sc_hs__buf_2
Xsky130_fd_sc_hs__buf_2_133 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__buf_2_133/A sky130_fd_sc_hs__buf_2_133/X
+ sky130_fd_sc_hs__buf_2_133/a_21_260# sky130_fd_sc_hs__buf_2
Xsky130_fd_sc_hs__buf_2_144 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__buf_2_151/X sky130_fd_sc_hs__buf_2_145/X
+ sky130_fd_sc_hs__buf_2_145/a_21_260# sky130_fd_sc_hs__buf_2
Xsky130_fd_sc_hs__buf_2_155 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__buf_2_155/A sky130_fd_sc_hs__buf_2_155/X
+ sky130_fd_sc_hs__buf_2_155/a_21_260# sky130_fd_sc_hs__buf_2
Xsky130_fd_sc_hs__einvp_2_12 DVSS: DVDD: DVDD: DVSS: dout_n sky130_fd_sc_hs__buf_8_1/A
+ sky130_fd_sc_hs__dlrtp_1_15/Q sky130_fd_sc_hs__einvp_2_13/a_263_323# sky130_fd_sc_hs__einvp_2_13/a_36_74#
+ sky130_fd_sc_hs__einvp_2_13/a_27_368# sky130_fd_sc_hs__einvp_2
Xsky130_fd_sc_hs__einvp_2_23 DVSS: DVDD: DVDD: DVSS: dout_n sky130_fd_sc_hs__einvp_2_9/A
+ sky130_fd_sc_hs__dlrtp_1_17/Q sky130_fd_sc_hs__einvp_2_23/a_263_323# sky130_fd_sc_hs__einvp_2_23/a_36_74#
+ sky130_fd_sc_hs__einvp_2_23/a_27_368# sky130_fd_sc_hs__einvp_2
Xsky130_fd_sc_hs__einvp_2_34 DVSS: DVDD: DVDD: DVSS: dout_n sky130_fd_sc_hs__buf_8_1/X
+ sky130_fd_sc_hs__buf_2_123/X sky130_fd_sc_hs__einvp_2_35/a_263_323# sky130_fd_sc_hs__einvp_2_35/a_36_74#
+ sky130_fd_sc_hs__einvp_2_35/a_27_368# sky130_fd_sc_hs__einvp_2
Xsky130_fd_sc_hs__einvp_2_45 DVSS: DVDD: DVDD: DVSS: dout_n sky130_fd_sc_hs__buf_8_1/A
+ sky130_fd_sc_hs__dlrtp_1_29/Q sky130_fd_sc_hs__einvp_2_45/a_263_323# sky130_fd_sc_hs__einvp_2_45/a_36_74#
+ sky130_fd_sc_hs__einvp_2_45/a_27_368# sky130_fd_sc_hs__einvp_2
Xsky130_fd_sc_hs__einvp_2_56 DVSS: DVDD: DVDD: DVSS: dout_p sky130_fd_sc_hs__einvp_2_65/A
+ sky130_fd_sc_hs__dlrtp_1_41/Q sky130_fd_sc_hs__einvp_2_57/a_263_323# sky130_fd_sc_hs__einvp_2_57/a_36_74#
+ sky130_fd_sc_hs__einvp_2_57/a_27_368# sky130_fd_sc_hs__einvp_2
Xsky130_fd_sc_hs__einvp_2_67 DVSS: DVDD: DVDD: DVSS: dout_p sky130_fd_sc_hs__einvp_2_99/A
+ sky130_fd_sc_hs__dlrtp_1_47/Q sky130_fd_sc_hs__einvp_2_67/a_263_323# sky130_fd_sc_hs__einvp_2_67/a_36_74#
+ sky130_fd_sc_hs__einvp_2_67/a_27_368# sky130_fd_sc_hs__einvp_2
Xsky130_fd_sc_hs__einvp_2_78 DVSS: DVDD: DVDD: DVSS: dout_p sky130_fd_sc_hs__einvp_2_97/A
+ sky130_fd_sc_hs__dlrtp_1_67/Q sky130_fd_sc_hs__einvp_2_79/a_263_323# sky130_fd_sc_hs__einvp_2_79/a_36_74#
+ sky130_fd_sc_hs__einvp_2_79/a_27_368# sky130_fd_sc_hs__einvp_2
Xsky130_fd_sc_hs__einvp_2_89 DVSS: DVDD: DVDD: DVSS: dout_p sky130_fd_sc_hs__einvp_2_97/A
+ sky130_fd_sc_hs__einvp_2_89/TE sky130_fd_sc_hs__einvp_2_89/a_263_323# sky130_fd_sc_hs__einvp_2_89/a_36_74#
+ sky130_fd_sc_hs__einvp_2_89/a_27_368# sky130_fd_sc_hs__einvp_2
Xsky130_fd_sc_hs__or2b_2_4 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__or2b_2_5/X sky130_fd_sc_hs__or2b_4_3/A
+ sky130_fd_sc_hs__or2b_2_5/A sky130_fd_sc_hs__or2b_2_5/a_470_368# sky130_fd_sc_hs__or2b_2_5/a_27_368#
+ sky130_fd_sc_hs__or2b_2_5/a_187_48# sky130_fd_sc_hs__or2b_2
Xsky130_fd_sc_hs__conb_1_11 DVSS: DVDD: DVDD: DVSS: prbs_generator_syn_3/eqn[4] prbs_generator_syn_3/eqn[1]
+ sky130_fd_sc_hs__conb_1_11/a_165_290# sky130_fd_sc_hs__conb_1_11/a_21_290# sky130_fd_sc_hs__conb_1
Xsky130_fd_sc_hs__conb_1_22 DVSS: DVDD: DVDD: DVSS: prbs_generator_syn_1/eqn[30] sky130_fd_sc_hs__conb_1_23/HI
+ sky130_fd_sc_hs__conb_1_23/a_165_290# sky130_fd_sc_hs__conb_1_23/a_21_290# sky130_fd_sc_hs__conb_1
Xsky130_fd_sc_hs__conb_1_33 DVSS: DVDD: DVDD: DVSS: prbs_generator_syn_5/eqn[31] prbs_generator_syn_5/cke
+ sky130_fd_sc_hs__conb_1_33/a_165_290# sky130_fd_sc_hs__conb_1_33/a_21_290# sky130_fd_sc_hs__conb_1
Xsky130_fd_sc_hs__conb_1_44 DVSS: DVDD: DVDD: DVSS: prbs_generator_syn_3/eqn[30] sky130_fd_sc_hs__conb_1_45/HI
+ sky130_fd_sc_hs__conb_1_45/a_165_290# sky130_fd_sc_hs__conb_1_45/a_21_290# sky130_fd_sc_hs__conb_1
Xsky130_fd_sc_hs__conb_1_55 DVSS: DVDD: DVDD: DVSS: prbs_generator_syn_9/eqn[30] sky130_fd_sc_hs__conb_1_55/HI
+ sky130_fd_sc_hs__conb_1_55/a_165_290# sky130_fd_sc_hs__conb_1_55/a_21_290# sky130_fd_sc_hs__conb_1
Xsky130_fd_sc_hs__conb_1_66 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__conb_1_67/LO
+ sky130_fd_sc_hs__conb_1_67/HI sky130_fd_sc_hs__conb_1_67/a_165_290# sky130_fd_sc_hs__conb_1_67/a_21_290#
+ sky130_fd_sc_hs__conb_1
Xsky130_fd_sc_hs__conb_1_77 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__conb_1_77/LO
+ sky130_fd_sc_hs__conb_1_77/HI sky130_fd_sc_hs__conb_1_77/a_165_290# sky130_fd_sc_hs__conb_1_77/a_21_290#
+ sky130_fd_sc_hs__conb_1
Xsky130_fd_sc_hs__inv_4_40 DVSS: DVDD: DVDD: DVSS: osc_core_1/pi2_r[2] osc_core_1/pi2_l[2]
+ sky130_fd_sc_hs__inv_4
Xsky130_fd_sc_hs__conb_1_88 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__conb_1_89/LO
+ sky130_fd_sc_hs__conb_1_89/HI sky130_fd_sc_hs__conb_1_89/a_165_290# sky130_fd_sc_hs__conb_1_89/a_21_290#
+ sky130_fd_sc_hs__conb_1
Xsky130_fd_sc_hs__conb_1_99 DVSS: DVDD: DVDD: DVSS: prbs_generator_syn_13/eqn[9] sky130_fd_sc_hs__conb_1_99/HI
+ sky130_fd_sc_hs__conb_1_99/a_165_290# sky130_fd_sc_hs__conb_1_99/a_21_290# sky130_fd_sc_hs__conb_1
Xsky130_fd_sc_hs__inv_4_51 DVSS: DVDD: DVDD: DVSS: osc_core_1/pi3_r[2] osc_core_1/pi3_l[2]
+ sky130_fd_sc_hs__inv_4
Xsky130_fd_sc_hs__inv_4_62 DVSS: DVDD: DVDD: DVSS: osc_core_1/pi4_r[1] osc_core_1/pi4_l[1]
+ sky130_fd_sc_hs__inv_4
Xsky130_fd_sc_hs__inv_4_73 DVSS: DVDD: DVDD: DVSS: osc_core_1/pi5_r[2] osc_core_1/pi5_l[2]
+ sky130_fd_sc_hs__inv_4
Xsky130_fd_sc_hs__inv_4_84 DVSS: DVDD: DVDD: DVSS: hr_16t4_mux_top_3/din[4] hr_16t4_mux_top_1/din[4]
+ sky130_fd_sc_hs__inv_4
Xsky130_fd_sc_hs__dlrtp_1_13 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__dlrtp_1_13/Q
+ sky130_fd_sc_hs__dlrtp_1_9/GATE sky130_fd_sc_hs__conb_1_117/HI sky130_fd_sc_hs__buf_2_109/X
+ sky130_fd_sc_hs__dlrtp_1_13/a_216_424# sky130_fd_sc_hs__dlrtp_1_13/a_759_508# sky130_fd_sc_hs__dlrtp_1_13/a_565_74#
+ sky130_fd_sc_hs__dlrtp_1_13/a_27_424# sky130_fd_sc_hs__dlrtp_1_13/a_1045_74# sky130_fd_sc_hs__dlrtp_1_13/a_643_74#
+ sky130_fd_sc_hs__dlrtp_1_13/a_817_48# sky130_fd_sc_hs__dlrtp_1_13/a_568_392# sky130_fd_sc_hs__dlrtp_1_13/a_363_74#
+ sky130_fd_sc_hs__dlrtp_1_13/a_769_74# sky130_fd_sc_hs__dlrtp_1
Xsky130_fd_sc_hs__dlrtp_1_24 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__dlrtp_1_24/Q
+ sky130_fd_sc_hs__clkbuf_2_3/X sky130_fd_sc_hs__conb_1_119/HI sky130_fd_sc_hs__dlrtp_1_24/D
+ sky130_fd_sc_hs__dlrtp_1_24/a_216_424# sky130_fd_sc_hs__dlrtp_1_24/a_759_508# sky130_fd_sc_hs__dlrtp_1_24/a_565_74#
+ sky130_fd_sc_hs__dlrtp_1_24/a_27_424# sky130_fd_sc_hs__dlrtp_1_24/a_1045_74# sky130_fd_sc_hs__dlrtp_1_24/a_643_74#
+ sky130_fd_sc_hs__dlrtp_1_24/a_817_48# sky130_fd_sc_hs__dlrtp_1_24/a_568_392# sky130_fd_sc_hs__dlrtp_1_24/a_363_74#
+ sky130_fd_sc_hs__dlrtp_1_24/a_769_74# sky130_fd_sc_hs__dlrtp_1
Xsky130_fd_sc_hs__dlrtp_1_35 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__dlrtp_1_35/Q
+ sky130_fd_sc_hs__clkbuf_2_3/A sky130_fd_sc_hs__conb_1_121/HI sky130_fd_sc_hs__dlrtp_1_35/D
+ sky130_fd_sc_hs__dlrtp_1_35/a_216_424# sky130_fd_sc_hs__dlrtp_1_35/a_759_508# sky130_fd_sc_hs__dlrtp_1_35/a_565_74#
+ sky130_fd_sc_hs__dlrtp_1_35/a_27_424# sky130_fd_sc_hs__dlrtp_1_35/a_1045_74# sky130_fd_sc_hs__dlrtp_1_35/a_643_74#
+ sky130_fd_sc_hs__dlrtp_1_35/a_817_48# sky130_fd_sc_hs__dlrtp_1_35/a_568_392# sky130_fd_sc_hs__dlrtp_1_35/a_363_74#
+ sky130_fd_sc_hs__dlrtp_1_35/a_769_74# sky130_fd_sc_hs__dlrtp_1
Xsky130_fd_sc_hs__dlrtp_1_46 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__dlrtp_1_47/Q
+ sky130_fd_sc_hs__clkbuf_16_53/A sky130_fd_sc_hs__conb_1_121/HI sky130_fd_sc_hs__buf_2_21/X
+ sky130_fd_sc_hs__dlrtp_1_47/a_216_424# sky130_fd_sc_hs__dlrtp_1_47/a_759_508# sky130_fd_sc_hs__dlrtp_1_47/a_565_74#
+ sky130_fd_sc_hs__dlrtp_1_47/a_27_424# sky130_fd_sc_hs__dlrtp_1_47/a_1045_74# sky130_fd_sc_hs__dlrtp_1_47/a_643_74#
+ sky130_fd_sc_hs__dlrtp_1_47/a_817_48# sky130_fd_sc_hs__dlrtp_1_47/a_568_392# sky130_fd_sc_hs__dlrtp_1_47/a_363_74#
+ sky130_fd_sc_hs__dlrtp_1_47/a_769_74# sky130_fd_sc_hs__dlrtp_1
Xsky130_fd_sc_hs__dlrtp_1_57 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__dlrtp_1_59/Q
+ sky130_fd_sc_hs__clkbuf_16_53/A sky130_fd_sc_hs__conb_1_125/HI sky130_fd_sc_hs__buf_2_55/X
+ sky130_fd_sc_hs__dlrtp_1_59/a_216_424# sky130_fd_sc_hs__dlrtp_1_59/a_759_508# sky130_fd_sc_hs__dlrtp_1_59/a_565_74#
+ sky130_fd_sc_hs__dlrtp_1_59/a_27_424# sky130_fd_sc_hs__dlrtp_1_59/a_1045_74# sky130_fd_sc_hs__dlrtp_1_59/a_643_74#
+ sky130_fd_sc_hs__dlrtp_1_59/a_817_48# sky130_fd_sc_hs__dlrtp_1_59/a_568_392# sky130_fd_sc_hs__dlrtp_1_59/a_363_74#
+ sky130_fd_sc_hs__dlrtp_1_59/a_769_74# sky130_fd_sc_hs__dlrtp_1
Xsky130_fd_sc_hs__dlrtp_1_68 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__dlrtp_1_69/Q
+ sky130_fd_sc_hs__clkbuf_16_53/A sky130_fd_sc_hs__conb_1_129/HI sky130_fd_sc_hs__dlrtp_1_69/D
+ sky130_fd_sc_hs__dlrtp_1_69/a_216_424# sky130_fd_sc_hs__dlrtp_1_69/a_759_508# sky130_fd_sc_hs__dlrtp_1_69/a_565_74#
+ sky130_fd_sc_hs__dlrtp_1_69/a_27_424# sky130_fd_sc_hs__dlrtp_1_69/a_1045_74# sky130_fd_sc_hs__dlrtp_1_69/a_643_74#
+ sky130_fd_sc_hs__dlrtp_1_69/a_817_48# sky130_fd_sc_hs__dlrtp_1_69/a_568_392# sky130_fd_sc_hs__dlrtp_1_69/a_363_74#
+ sky130_fd_sc_hs__dlrtp_1_69/a_769_74# sky130_fd_sc_hs__dlrtp_1
Xsky130_fd_sc_hs__dlrtp_1_79 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__dlrtp_1_79/Q
+ sky130_fd_sc_hs__clkbuf_16_53/X sky130_fd_sc_hs__conb_1_129/HI sky130_fd_sc_hs__dlrtp_1_79/D
+ sky130_fd_sc_hs__dlrtp_1_79/a_216_424# sky130_fd_sc_hs__dlrtp_1_79/a_759_508# sky130_fd_sc_hs__dlrtp_1_79/a_565_74#
+ sky130_fd_sc_hs__dlrtp_1_79/a_27_424# sky130_fd_sc_hs__dlrtp_1_79/a_1045_74# sky130_fd_sc_hs__dlrtp_1_79/a_643_74#
+ sky130_fd_sc_hs__dlrtp_1_79/a_817_48# sky130_fd_sc_hs__dlrtp_1_79/a_568_392# sky130_fd_sc_hs__dlrtp_1_79/a_363_74#
+ sky130_fd_sc_hs__dlrtp_1_79/a_769_74# sky130_fd_sc_hs__dlrtp_1
Xsky130_fd_sc_hs__einvp_2_6 DVSS: DVDD: DVDD: DVSS: dout_n sky130_fd_sc_hs__buf_8_1/A
+ sky130_fd_sc_hs__dlrtp_1_3/Q sky130_fd_sc_hs__einvp_2_7/a_263_323# sky130_fd_sc_hs__einvp_2_7/a_36_74#
+ sky130_fd_sc_hs__einvp_2_7/a_27_368# sky130_fd_sc_hs__einvp_2
Xsky130_fd_sc_hs__clkbuf_2_9 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__dlrtp_1_58/D
+ sky130_fd_sc_hs__o21bai_2_3/Y sky130_fd_sc_hs__clkbuf_2_9/a_43_192# sky130_fd_sc_hs__clkbuf_2
Xfine_freq_track_0 osc_core_1/p3 sky130_fd_sc_hs__clkbuf_4_89/X sky130_fd_sc_hs__clkbuf_4_91/X
+ sky130_fd_sc_hs__clkbuf_4_93/X sky130_fd_sc_hs__clkbuf_4_95/X sky130_fd_sc_hs__clkbuf_4_97/X
+ sky130_fd_sc_hs__clkbuf_4_99/X osc_core_1/ref_clk qr_4t1_mux_top_1/rst fine_freq_track_1/aux_osc_en
+ fine_freq_track_1/fftl_en sky130_fd_sc_hs__clkbuf_4_65/X sky130_fd_sc_hs__clkbuf_4_61/X
+ sky130_fd_sc_hs__clkbuf_4_63/X sky130_fd_sc_hs__clkinv_2_3/Y sky130_fd_sc_hs__clkbuf_4_67/X
+ sky130_fd_sc_hs__clkbuf_4_53/X sky130_fd_sc_hs__clkbuf_4_57/X sky130_fd_sc_hs__clkbuf_4_59/X
+ sky130_fd_sc_hs__clkbuf_4_55/X sky130_fd_sc_hs__clkbuf_8_15/X sky130_fd_sc_hs__clkbuf_8_17/X
+ sky130_fd_sc_hs__clkbuf_8_19/X sky130_fd_sc_hs__clkbuf_8_13/X sky130_fd_sc_hs__clkbuf_8_21/X
+ sky130_fd_sc_hs__clkbuf_16_19/X sky130_fd_sc_hs__clkbuf_16_17/X sky130_fd_sc_hs__clkbuf_8_23/X
+ sky130_fd_sc_hs__clkbuf_8_25/X sky130_fd_sc_hs__clkbuf_8_27/X sky130_fd_sc_hs__clkbuf_8_29/X
+ sky130_fd_sc_hs__clkbuf_8_31/X sky130_fd_sc_hs__clkbuf_4_41/X sky130_fd_sc_hs__einvp_8_5/A
+ fine_freq_track_1/out_star osc_core_1/delay_con_msb[7] osc_core_1/delay_con_msb[6]
+ osc_core_1/delay_con_msb[5] osc_core_1/delay_con_msb[4] osc_core_1/delay_con_msb[3]
+ osc_core_1/delay_con_msb[2] osc_core_1/delay_con_msb[1] osc_core_1/delay_con_msb[0]
+ osc_core_1/delay_con_lsb[4] osc_core_1/delay_con_lsb[3] osc_core_1/delay_con_lsb[2]
+ osc_core_1/delay_con_lsb[1] osc_core_1/delay_con_lsb[0] DVSS: DVDD: fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_9/a_1827_81#
+ fine_freq_track_1/sky130_fd_sc_hs__nor2b_1_23/Y fine_freq_track_1/sky130_fd_sc_hs__o21a_1_51/B1
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_19/a_498_360# fine_freq_track_1/sky130_fd_sc_hs__inv_4_65/Y
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_79/a_1350_392# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_63/a_789_463#
+ fine_freq_track_1/sky130_fd_sc_hs__dfstp_2_4/a_2022_94# fine_freq_track_1/sky130_fd_sc_hs__nor2_1_35/B
+ fine_freq_track_1/sky130_fd_sc_hs__dfstp_2_7/a_1278_74# fine_freq_track_1/sky130_fd_sc_hs__nor2_1_3/a_116_368#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_15/a_706_463# fine_freq_track_1/sky130_fd_sc_hs__inv_2_7/Y
+ fine_freq_track_1/sky130_fd_sc_hs__a22o_1_27/a_222_392# fine_freq_track_1/sky130_fd_sc_hs__a32oi_1_3/Y
+ fine_freq_track_1/sky130_fd_sc_hs__a22o_1_21/a_52_123# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_3/a_37_78#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_75/a_1678_395# fine_freq_track_1/sky130_fd_sc_hs__inv_4_45/A
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_45/a_834_355# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_37/a_1627_493#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_45/a_319_360# fine_freq_track_1/sky130_fd_sc_hs__fa_2_11/a_1205_79#
+ fine_freq_track_1/sky130_fd_sc_hs__fa_2_1/CIN fine_freq_track_1/sky130_fd_sc_hs__nor2_1_31/Y
+ fine_freq_track_1/sky130_fd_sc_hs__a32oi_1_3/B1 fine_freq_track_1/sky130_fd_sc_hs__nand2_4_13/Y
+ fine_freq_track_1/sky130_fd_sc_hs__nand3_1_1/a_155_74# fine_freq_track_1/sky130_fd_sc_hs__nor2_1_37/B
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_59/a_313_74# fine_freq_track_1/sky130_fd_sc_hs__sdlclkp_1_1/a_114_112#
+ fine_freq_track_1/sky130_fd_sc_hs__nor2b_1_25/Y fine_freq_track_1/sky130_fd_sc_hs__o21a_1_7/A1
+ fine_freq_track_1/sky130_fd_sc_hs__sdlclkp_4_1/a_634_74# fine_freq_track_1/sky130_fd_sc_hs__nor4_1_1/D
+ fine_freq_track_1/sky130_fd_sc_hs__inv_4_63/Y fine_freq_track_1/sky130_fd_sc_hs__inv_4_125/A
+ fine_freq_track_1/sky130_fd_sc_hs__inv_4_59/A fine_freq_track_1/sky130_fd_sc_hs__dfxtp_2_3/a_1217_314#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_25/a_313_74# fine_freq_track_1/sky130_fd_sc_hs__clkbuf_8_1/X
+ fine_freq_track_1/sky130_fd_sc_hs__inv_4_47/A fine_freq_track_1/sky130_fd_sc_hs__o21a_1_5/X
+ fine_freq_track_1/sky130_fd_sc_hs__o21a_1_37/a_376_387# fine_freq_track_1/sky130_fd_sc_hs__inv_4_55/Y
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_39/a_890_138# fine_freq_track_1/sky130_fd_sc_hs__clkbuf_2_1/X
+ fine_freq_track_1/sky130_fd_sc_hs__dfxtp_2_9/a_206_368# fine_freq_track_1/sky130_fd_sc_hs__xnor2_1_3/B
+ fine_freq_track_1/sky130_fd_sc_hs__nor2_1_61/B fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_25/a_125_78#
+ fine_freq_track_1/sky130_fd_sc_hs__o21a_1_77/a_376_387# fine_freq_track_1/sky130_fd_sc_hs__dfsbp_2_1/a_225_74#
+ fine_freq_track_1/sky130_fd_sc_hs__nor2b_1_7/a_27_112# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_7/a_714_127#
+ fine_freq_track_1/sky130_fd_sc_hs__o21a_1_77/a_83_244# fine_freq_track_1/sky130_fd_sc_hs__nand2_1_9/A
+ fine_freq_track_1/sky130_fd_sc_hs__nand2_1_113/a_117_74# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_15/a_38_78#
+ fine_freq_track_1/sky130_fd_sc_hs__inv_4_135/Y fine_freq_track_1/sky130_fd_sc_hs__nand4_2_1/B
+ fine_freq_track_1/sky130_fd_sc_hs__inv_4_73/A fine_freq_track_1/sky130_fd_sc_hs__nand2_1_47/B
+ fine_freq_track_1/sky130_fd_sc_hs__nor2_1_43/a_116_368# fine_freq_track_1/sky130_fd_sc_hs__a22oi_1_19/a_339_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_5/a_1224_74# fine_freq_track_1/sky130_fd_sc_hs__xnor2_1_15/Y
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_43/D fine_freq_track_1/sky130_fd_sc_hs__inv_4_137/A
+ fine_freq_track_1/sky130_fd_sc_hs__dfstp_2_1/CLK fine_freq_track_1/sky130_fd_sc_hs__nor2_1_41/Y
+ fine_freq_track_1/sky130_fd_sc_hs__dfxtp_4_2/a_1141_508# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_5/a_124_78#
+ fine_freq_track_1/sky130_fd_sc_hs__inv_4_103/A fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_23/D
+ fine_freq_track_1/sky130_fd_sc_hs__nor2_1_45/B fine_freq_track_1/sky130_fd_sc_hs__nor2b_1_45/a_27_112#
+ fine_freq_track_1/sky130_fd_sc_hs__dfstp_2_7/Q fine_freq_track_1/sky130_fd_sc_hs__a31oi_2_1/Y
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_81/a_699_463# fine_freq_track_1/sky130_fd_sc_hs__o22ai_1_9/B1
+ fine_freq_track_1/sky130_fd_sc_hs__xnor2_1_1/B fine_freq_track_1/sky130_fd_sc_hs__nor2b_1_19/a_278_368#
+ fine_freq_track_1/sky130_fd_sc_hs__nor3_1_5/Y fine_freq_track_1/sky130_fd_sc_hs__inv_4_87/Y
+ fine_freq_track_1/sky130_fd_sc_hs__nand2_1_77/a_117_74# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_43/a_841_401#
+ fine_freq_track_1/sky130_fd_sc_hs__o22ai_1_9/a_27_74# fine_freq_track_1/sky130_fd_sc_hs__inv_4_133/Y
+ fine_freq_track_1/sky130_fd_sc_hs__nor3_1_1/a_198_368# fine_freq_track_1/sky130_fd_sc_hs__o21a_1_71/A1
+ fine_freq_track_1/sky130_fd_sc_hs__a22o_1_3/a_222_392# fine_freq_track_1/sky130_fd_sc_hs__a21oi_1_97/Y
+ fine_freq_track_1/sky130_fd_sc_hs__nor3_1_13/A fine_freq_track_1/sky130_fd_sc_hs__inv_4_17/Y
+ fine_freq_track_1/sky130_fd_sc_hs__nand2_1_43/a_117_74# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_45/a_812_138#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_23/a_856_304# fine_freq_track_1/sky130_fd_sc_hs__o31ai_1_1/a_119_368#
+ fine_freq_track_1/sky130_fd_sc_hs__fa_2_21/a_27_79# fine_freq_track_1/sky130_fd_sc_hs__o211ai_1_7/a_311_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_23/a_850_127# fine_freq_track_1/sky130_fd_sc_hs__nor3_1_13/C
+ fine_freq_track_1/sky130_fd_sc_hs__nand2_1_11/a_117_74# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_17/a_33_74#
+ fine_freq_track_1/sky130_fd_sc_hs__nand4_1_5/C fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_29/a_1647_81#
+ fine_freq_track_1/sky130_fd_sc_hs__fa_2_21/a_484_347# fine_freq_track_1/sky130_fd_sc_hs__dfxtp_2_3/a_695_459#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_81/a_124_78# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_31/a_38_78#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_67/a_1647_81# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_29/a_1224_74#
+ fine_freq_track_1/sky130_fd_sc_hs__inv_4_75/A fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_5/a_38_78#
+ fine_freq_track_1/sky130_fd_sc_hs__nand2_1_5/a_117_74# fine_freq_track_1/sky130_fd_sc_hs__nor2_1_51/Y
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_41/a_507_368# fine_freq_track_1/sky130_fd_sc_hs__or3b_2_1/a_458_368#
+ fine_freq_track_1/sky130_fd_sc_hs__o21a_1_71/a_320_74# fine_freq_track_1/sky130_fd_sc_hs__a21oi_1_27/a_29_368#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_43/Q_N fine_freq_track_1/sky130_fd_sc_hs__nor2_1_37/Y
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_53/a_789_463# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_47/a_498_360#
+ fine_freq_track_1/sky130_fd_sc_hs__dfstp_2_1/a_767_384# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_49/a_1547_508#
+ fine_freq_track_1/sky130_fd_sc_hs__a22o_1_17/a_222_392# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_35/Q_N
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_73/a_1678_395# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_35/a_834_355#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_91/a_37_78# fine_freq_track_1/sky130_fd_sc_hs__fa_2_7/a_27_79#
+ fine_freq_track_1/sky130_fd_sc_hs__xnor2_1_7/Y fine_freq_track_1/sky130_fd_sc_hs__a21oi_1_9/a_29_368#
+ fine_freq_track_1/sky130_fd_sc_hs__a21oi_1_71/a_29_368# fine_freq_track_1/sky130_fd_sc_hs__xor2_1_5/a_455_87#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_25/Q_N fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_43/D
+ fine_freq_track_1/sky130_fd_sc_hs__inv_4_85/Y fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_73/a_834_355#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_39/a_922_127# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_27/a_1350_392#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_21/D fine_freq_track_1/sky130_fd_sc_hs__maj3_1_3/a_598_384#
+ fine_freq_track_1/sky130_fd_sc_hs__nor2_1_47/B fine_freq_track_1/sky130_fd_sc_hs__o21a_1_15/A1
+ fine_freq_track_1/sky130_fd_sc_hs__inv_4_65/A fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_33/a_33_74#
+ fine_freq_track_1/sky130_fd_sc_hs__a22oi_1_15/Y fine_freq_track_1/sky130_fd_sc_hs__o21a_1_9/a_83_244#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_23/a_1678_395# fine_freq_track_1/sky130_fd_sc_hs__o21a_1_27/a_376_387#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_41/a_2026_424# fine_freq_track_1/sky130_fd_sc_hs__inv_4_37/A
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_23/a_832_118# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_29/a_890_138#
+ fine_freq_track_1/sky130_fd_sc_hs__a22oi_1_21/Y fine_freq_track_1/sky130_fd_sc_hs__o21a_1_67/a_376_387#
+ fine_freq_track_1/sky130_fd_sc_hs__maj3_1_1/a_595_136# fine_freq_track_1/sky130_fd_sc_hs__or2_1_3/A
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_25/a_1465_471# fine_freq_track_1/sky130_fd_sc_hs__a21oi_1_17/Y
+ fine_freq_track_1/sky130_fd_sc_hs__inv_4_45/Y fine_freq_track_1/sky130_fd_sc_hs__nor3_1_5/A
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_67/a_890_138# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_13/D
+ fine_freq_track_1/sky130_fd_sc_hs__xor2_1_11/B fine_freq_track_1/sky130_fd_sc_hs__o21a_1_35/X
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_57/a_2010_409# fine_freq_track_1/sky130_fd_sc_hs__nor4_1_1/C
+ fine_freq_track_1/sky130_fd_sc_hs__a21oi_1_57/a_117_74# fine_freq_track_1/sky130_fd_sc_hs__or3b_2_1/B
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_37/a_817_508# fine_freq_track_1/sky130_fd_sc_hs__a211oi_1_1/Y
+ fine_freq_track_1/sky130_fd_sc_hs__nor2_1_97/A fine_freq_track_1/sky130_fd_sc_hs__inv_4_79/Y
+ fine_freq_track_1/sky130_fd_sc_hs__dfxtp_4_9/a_27_74# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_41/a_910_118#
+ fine_freq_track_1/sky130_fd_sc_hs__nor2_1_33/a_116_368# fine_freq_track_1/sky130_fd_sc_hs__inv_4_43/Y
+ fine_freq_track_1/sky130_fd_sc_hs__nor2_1_71/a_116_368# fine_freq_track_1/sky130_fd_sc_hs__nand2_2_3/A
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_7/a_699_463# fine_freq_track_1/sky130_fd_sc_hs__nand2_2_3/a_27_74#
+ fine_freq_track_1/sky130_fd_sc_hs__inv_4_41/Y fine_freq_track_1/sky130_fd_sc_hs__o21ai_2_1/B1
+ fine_freq_track_1/sky130_fd_sc_hs__a31oi_2_1/A1 fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_71/a_699_463#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_31/a_300_74# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_59/D
+ fine_freq_track_1/sky130_fd_sc_hs__a21oi_1_105/a_29_368# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_73/a_313_74#
+ fine_freq_track_1/sky130_fd_sc_hs__nor2_1_87/Y fine_freq_track_1/sky130_fd_sc_hs__nand2_1_117/a_117_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_37/a_1624_74# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_1/a_319_360#
+ fine_freq_track_1/sky130_fd_sc_hs__nor3_1_9/Y fine_freq_track_1/sky130_fd_sc_hs__inv_4_129/A
+ fine_freq_track_1/sky130_fd_sc_hs__dfstp_2_5/a_27_74# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_3/a_1736_119#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_35/a_812_138# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_41/a_313_74#
+ fine_freq_track_1/sky130_fd_sc_hs__inv_4_69/A fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_37/D
+ fine_freq_track_1/sky130_fd_sc_hs__inv_4_129/Y fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_3/a_1266_119#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_73/a_812_138# fine_freq_track_1/sky130_fd_sc_hs__nor2_1_35/Y
+ fine_freq_track_1/sky130_fd_sc_hs__fa_2_3/a_27_378# fine_freq_track_1/sky130_fd_sc_hs__o21a_1_15/a_83_244#
+ fine_freq_track_1/sky130_fd_sc_hs__or2_1_1/A fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_9/a_124_78#
+ fine_freq_track_1/sky130_fd_sc_hs__xor2_1_9/A fine_freq_track_1/sky130_fd_sc_hs__inv_4_77/Y
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_19/a_1647_81# fine_freq_track_1/sky130_fd_sc_hs__maj3_1_1/A
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_87/a_1627_493# fine_freq_track_1/sky130_fd_sc_hs__o21a_1_23/A1
+ fine_freq_track_1/sky130_fd_sc_hs__nor4_1_3/Y fine_freq_track_1/sky130_fd_sc_hs__nor2_2_1/Y
+ fine_freq_track_1/sky130_fd_sc_hs__inv_4_55/A fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_45/a_37_78#
+ fine_freq_track_1/sky130_fd_sc_hs__inv_4_113/Y fine_freq_track_1/sky130_fd_sc_hs__maj3_1_3/A
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_19/a_1224_74# fine_freq_track_1/sky130_fd_sc_hs__fa_2_3/CIN
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_31/a_507_368# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_77/a_1350_392#
+ fine_freq_track_1/sky130_fd_sc_hs__nor4_1_1/a_342_368# fine_freq_track_1/sky130_fd_sc_hs__o21a_1_65/B1
+ fine_freq_track_1/sky130_fd_sc_hs__xor2_1_11/a_455_87# fine_freq_track_1/sky130_fd_sc_hs__xor2_1_9/a_158_392#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_47/a_1547_508# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_83/a_789_463#
+ fine_freq_track_1/sky130_fd_sc_hs__a22oi_1_5/Y fine_freq_track_1/sky130_fd_sc_hs__inv_4_11/A
+ fine_freq_track_1/sky130_fd_sc_hs__nand2_1_15/a_117_74# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_35/a_706_463#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_25/a_319_360# fine_freq_track_1/sky130_fd_sc_hs__inv_4_49/Y
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_63/a_834_355# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_49/a_494_366#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_85/a_124_78# fine_freq_track_1/sky130_fd_sc_hs__and2_2_5/a_31_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_7/a_1934_94# fine_freq_track_1/sky130_fd_sc_hs__nand2_4_9/Y
+ fine_freq_track_1/sky130_fd_sc_hs__fa_2_3/a_701_79# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_29/a_922_127#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_9/a_1598_93# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_25/a_1350_392#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_89/a_494_366# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_7/D
+ fine_freq_track_1/sky130_fd_sc_hs__o211ai_1_9/a_116_368# fine_freq_track_1/sky130_fd_sc_hs__o21a_1_75/a_320_74#
+ fine_freq_track_1/sky130_fd_sc_hs__nor2_1_31/B fine_freq_track_1/sky130_fd_sc_hs__fa_2_11/SUM
+ fine_freq_track_1/sky130_fd_sc_hs__dfxtp_2_1/a_1217_314# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_43/a_1434_74#
+ fine_freq_track_1/sky130_fd_sc_hs__xnor2_1_3/A fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_3/a_1624_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfxtp_4_3/a_206_368# fine_freq_track_1/sky130_fd_sc_hs__nor2_1_27/B
+ fine_freq_track_1/sky130_fd_sc_hs__a22o_1_29/X fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_21/a_1678_395#
+ fine_freq_track_1/sky130_fd_sc_hs__xnor2_1_3/a_112_119# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_13/a_832_118#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_19/a_890_138# fine_freq_track_1/sky130_fd_sc_hs__a21oi_1_75/a_29_368#
+ fine_freq_track_1/sky130_fd_sc_hs__xor2_1_9/a_455_87# fine_freq_track_1/sky130_fd_sc_hs__o21a_1_57/a_376_387#
+ fine_freq_track_1/sky130_fd_sc_hs__a31oi_2_1/a_200_74# fine_freq_track_1/sky130_fd_sc_hs__inv_4_63/A
+ fine_freq_track_1/sky130_fd_sc_hs__xor2_1_9/X fine_freq_track_1/sky130_fd_sc_hs__o21a_1_65/X
+ fine_freq_track_1/sky130_fd_sc_hs__a32oi_1_7/B1 fine_freq_track_1/sky130_fd_sc_hs__fa_2_5/a_992_347#
+ fine_freq_track_1/sky130_fd_sc_hs__or2_1_3/X fine_freq_track_1/sky130_fd_sc_hs__dfxtp_4_5/a_696_458#
+ fine_freq_track_1/sky130_fd_sc_hs__nor2_1_7/Y fine_freq_track_1/sky130_fd_sc_hs__o21ai_1_3/B1
+ fine_freq_track_1/sky130_fd_sc_hs__inv_2_1/A fine_freq_track_1/sky130_fd_sc_hs__nor2_1_23/a_116_368#
+ fine_freq_track_1/sky130_fd_sc_hs__o21a_1_3/a_376_387# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_21/a_699_463#
+ fine_freq_track_1/sky130_fd_sc_hs__nor2b_1_5/a_278_368# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_7/D
+ fine_freq_track_1/sky130_fd_sc_hs__nand2_4_9/a_27_74# fine_freq_track_1/sky130_fd_sc_hs__o21a_1_73/A2
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_61/a_699_463# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_37/a_1550_119#
+ fine_freq_track_1/sky130_fd_sc_hs__nor2_1_107/a_116_368# fine_freq_track_1/sky130_fd_sc_hs__nor2_1_65/Y
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_23/a_841_401# fine_freq_track_1/sky130_fd_sc_hs__nand2_1_59/Y
+ fine_freq_track_1/sky130_fd_sc_hs__fa_2_15/a_336_347# fine_freq_track_1/sky130_fd_sc_hs__nor2_1_63/B
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_1/a_1736_119# fine_freq_track_1/sky130_fd_sc_hs__inv_4_3/A
+ fine_freq_track_1/sky130_fd_sc_hs__inv_4_105/A fine_freq_track_1/sky130_fd_sc_hs__dfxtp_2_9/a_708_101#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_1/a_1266_119# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_63/a_812_138#
+ fine_freq_track_1/sky130_fd_sc_hs__nor2_1_25/B fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_41/a_856_304#
+ fine_freq_track_1/sky130_fd_sc_hs__a32oi_1_9/Y fine_freq_track_1/sky130_fd_sc_hs__o21a_1_25/A1
+ fine_freq_track_1/sky130_fd_sc_hs__fa_2_15/a_27_79# fine_freq_track_1/sky130_fd_sc_hs__o21a_1_27/X
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_41/a_850_127# fine_freq_track_1/sky130_fd_sc_hs__o31ai_1_1/B1
+ fine_freq_track_1/sky130_fd_sc_hs__a21oi_1_109/a_29_368# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_7/a_125_78#
+ fine_freq_track_1/sky130_fd_sc_hs__inv_4_81/Y fine_freq_track_1/sky130_fd_sc_hs__o22ai_1_11/a_340_368#
+ fine_freq_track_1/sky130_fd_sc_hs__fa_2_7/a_683_347# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_47/a_1647_81#
+ fine_freq_track_1/sky130_fd_sc_hs__o22ai_1_1/a_340_368# fine_freq_track_1/sky130_fd_sc_hs__fa_2_19/CIN
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_43/a_1827_81# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_21/a_507_368#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_87/a_1647_81# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_47/a_1224_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfxtp_4_7/D fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_45/a_313_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_9/a_789_463# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_27/a_498_360#
+ fine_freq_track_1/sky130_fd_sc_hs__nor3_1_11/a_114_368# fine_freq_track_1/sky130_fd_sc_hs__nor2_1_27/Y
+ fine_freq_track_1/sky130_fd_sc_hs__xnor2_1_11/a_112_119# fine_freq_track_1/sky130_fd_sc_hs__a222oi_1_3/a_116_392#
+ fine_freq_track_1/sky130_fd_sc_hs__xnor2_1_1/A fine_freq_track_1/sky130_fd_sc_hs__fa_2_7/a_27_378#
+ fine_freq_track_1/sky130_fd_sc_hs__o21a_1_19/a_83_244# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_35/a_1627_493#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_15/a_319_360# fine_freq_track_1/sky130_fd_sc_hs__maj3_1_1/C
+ fine_freq_track_1/sky130_fd_sc_hs__clkbuf_8_1/A fine_freq_track_1/sky130_fd_sc_hs__nor2_1_17/Y
+ fine_freq_track_1/sky130_fd_sc_hs__a21oi_1_121/a_29_368# fine_freq_track_1/sky130_fd_sc_hs__fa_2_17/a_683_347#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_53/a_834_355# fine_freq_track_1/sky130_fd_sc_hs__maj3_1_3/B
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_85/a_37_78# fine_freq_track_1/sky130_fd_sc_hs__nor3_1_3/A
+ fine_freq_track_1/sky130_fd_sc_hs__nor4_1_1/a_144_368# fine_freq_track_1/sky130_fd_sc_hs__fa_2_21/a_1205_79#
+ fine_freq_track_1/sky130_fd_sc_hs__o21a_1_59/A1 fine_freq_track_1/sky130_fd_sc_hs__o21ai_1_7/a_162_368#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_19/a_922_127# fine_freq_track_1/sky130_fd_sc_hs__o21a_1_63/a_83_244#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_79/a_494_366# fine_freq_track_1/sky130_fd_sc_hs__maj3_1_1/a_223_120#
+ fine_freq_track_1/sky130_fd_sc_hs__inv_4_79/A fine_freq_track_1/sky130_fd_sc_hs__inv_4_21/Y
+ fine_freq_track_1/sky130_fd_sc_hs__nand4_1_3/a_373_74# fine_freq_track_1/sky130_fd_sc_hs__fa_2_21/a_487_79#
+ fine_freq_track_1/sky130_fd_sc_hs__nor2_1_9/Y fine_freq_track_1/sky130_fd_sc_hs__inv_4_13/A
+ fine_freq_track_1/sky130_fd_sc_hs__nand2_1_19/a_117_74# fine_freq_track_1/sky130_fd_sc_hs__dfstp_2_1/a_612_74#
+ fine_freq_track_1/sky130_fd_sc_hs__nor3_1_1/Y fine_freq_track_1/sky130_fd_sc_hs__o21a_1_47/a_376_387#
+ fine_freq_track_1/sky130_fd_sc_hs__o21ai_1_3/a_27_74# fine_freq_track_1/sky130_fd_sc_hs__inv_4_125/Y
+ fine_freq_track_1/sky130_fd_sc_hs__dfxtp_4_3/a_437_503# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_23/a_1465_471#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_47/a_890_138# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_89/a_124_78#
+ fine_freq_track_1/sky130_fd_sc_hs__nor2b_1_31/a_27_112# fine_freq_track_1/sky130_fd_sc_hs__nor2_4_1/B
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_55/a_2010_409# fine_freq_track_1/sky130_fd_sc_hs__fa_2_7/a_701_79#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_87/a_890_138# fine_freq_track_1/sky130_fd_sc_hs__nor3_1_9/B
+ fine_freq_track_1/sky130_fd_sc_hs__o21a_1_73/B1 fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_37/D
+ fine_freq_track_1/sky130_fd_sc_hs__nor2_1_13/a_116_368# fine_freq_track_1/sky130_fd_sc_hs__nor4_1_3/B
+ fine_freq_track_1/sky130_fd_sc_hs__or3b_2_1/X fine_freq_track_1/sky130_fd_sc_hs__nor3_1_11/B
+ fine_freq_track_1/sky130_fd_sc_hs__inv_4_39/A fine_freq_track_1/sky130_fd_sc_hs__nor2_1_83/B
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_23/a_124_78# fine_freq_track_1/sky130_fd_sc_hs__dfsbp_2_1/a_2221_74#
+ fine_freq_track_1/sky130_fd_sc_hs__fa_2_19/SUM fine_freq_track_1/sky130_fd_sc_hs__nor2b_1_7/Y
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_51/a_699_463# fine_freq_track_1/sky130_fd_sc_hs__nor2_1_91/a_116_368#
+ fine_freq_track_1/sky130_fd_sc_hs__inv_4_67/Y fine_freq_track_1/sky130_fd_sc_hs__nand2_4_7/Y
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_13/a_841_401# fine_freq_track_1/sky130_fd_sc_hs__a32oi_1_7/A1
+ fine_freq_track_1/sky130_fd_sc_hs__a22o_1_13/a_132_392# fine_freq_track_1/sky130_fd_sc_hs__o31ai_1_1/a_203_368#
+ fine_freq_track_1/sky130_fd_sc_hs__o21a_1_75/B1 fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_3/D
+ fine_freq_track_1/sky130_fd_sc_hs__nor2_1_45/Y fine_freq_track_1/sky130_fd_sc_hs__a21oi_1_13/a_29_368#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_41/a_33_74# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_53/a_812_138#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_31/a_856_304# fine_freq_track_1/sky130_fd_sc_hs__nor2_1_5/Y
+ fine_freq_track_1/sky130_fd_sc_hs__nor4_1_1/a_228_368# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_31/a_850_127#
+ fine_freq_track_1/sky130_fd_sc_hs__nor3_1_1/B fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_85/a_1627_493#
+ fine_freq_track_1/sky130_fd_sc_hs__or3b_2_1/a_542_368# fine_freq_track_1/sky130_fd_sc_hs__o21a_1_53/B1
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_37/a_1647_81# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_3/a_1647_81#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_33/a_1827_81# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_39/a_714_127#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_11/a_507_368# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_77/a_1647_81#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_39/a_37_78# fine_freq_track_1/sky130_fd_sc_hs__inv_2_5/Y
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_75/a_1350_392# fine_freq_track_1/sky130_fd_sc_hs__a32oi_1_1/Y
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_17/a_498_360# fine_freq_track_1/sky130_fd_sc_hs__fa_2_11/B
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_31/a_796_463# fine_freq_track_1/sky130_fd_sc_hs__o211ai_1_3/Y
+ fine_freq_track_1/sky130_fd_sc_hs__nor2_1_25/Y fine_freq_track_1/sky130_fd_sc_hs__dfstp_2_1/a_2022_94#
+ fine_freq_track_1/sky130_fd_sc_hs__o22ai_1_11/a_142_368# fine_freq_track_1/sky130_fd_sc_hs__o22ai_1_1/a_142_368#
+ fine_freq_track_1/sky130_fd_sc_hs__nor2_1_1/a_116_368# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_71/a_1678_395#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_39/a_300_74# fine_freq_track_1/sky130_fd_sc_hs__nor2_1_87/B
+ fine_freq_track_1/sky130_fd_sc_hs__fa_2_13/B fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_83/a_834_355#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_69/a_494_366# fine_freq_track_1/sky130_fd_sc_hs__a21oi_1_1/Y
+ fine_freq_track_1/sky130_fd_sc_hs__inv_4_53/Y fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_49/a_922_127#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_23/a_1434_74# fine_freq_track_1/sky130_fd_sc_hs__a21oi_1_43/a_117_74#
+ fine_freq_track_1/sky130_fd_sc_hs__o22ai_1_1/Y fine_freq_track_1/sky130_fd_sc_hs__a32oi_1_3/a_469_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_15/a_313_74# fine_freq_track_1/sky130_fd_sc_hs__dfxtp_4_9/CLK
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_39/a_1678_395# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_33/a_832_118#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_37/a_890_138# fine_freq_track_1/sky130_fd_sc_hs__dfxtp_2_7/a_206_368#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_53/a_37_78# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_15/a_125_78#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_3/a_890_138# fine_freq_track_1/sky130_fd_sc_hs__inv_4_87/A
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_53/a_2010_409# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_77/a_890_138#
+ fine_freq_track_1/sky130_fd_sc_hs__o21a_1_67/a_83_244# fine_freq_track_1/sky130_fd_sc_hs__nand4_2_1/C
+ fine_freq_track_1/sky130_fd_sc_hs__inv_4_59/Y fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_41/D
+ fine_freq_track_1/sky130_fd_sc_hs__nand2_2_1/Y fine_freq_track_1/sky130_fd_sc_hs__nand2_1_103/a_117_74#
+ fine_freq_track_1/sky130_fd_sc_hs__o21a_1_63/A1 fine_freq_track_1/sky130_fd_sc_hs__maj3_1_1/B
+ fine_freq_track_1/sky130_fd_sc_hs__fa_2_3/B fine_freq_track_1/sky130_fd_sc_hs__nor2_1_41/a_116_368#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_7/a_796_463# fine_freq_track_1/sky130_fd_sc_hs__dfsbp_2_1/a_1339_74#
+ fine_freq_track_1/sky130_fd_sc_hs__o21a_1_67/B1 fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_41/a_699_463#
+ fine_freq_track_1/sky130_fd_sc_hs__nand2_1_99/a_117_74# fine_freq_track_1/sky130_fd_sc_hs__nor2_1_81/a_116_368#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_35/a_1550_119# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_5/a_37_78#
+ fine_freq_track_1/sky130_fd_sc_hs__nor2_4_3/a_27_368# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_29/Q_N
+ fine_freq_track_1/sky130_fd_sc_hs__nand2_1_67/a_117_74# fine_freq_track_1/sky130_fd_sc_hs__o21a_1_59/X
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_45/a_1624_74# fine_freq_track_1/sky130_fd_sc_hs__nor2_1_29/Y
+ fine_freq_track_1/sky130_fd_sc_hs__or2_1_3/B fine_freq_track_1/sky130_fd_sc_hs__xnor2_1_5/B
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_27/a_124_78# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_21/a_856_304#
+ fine_freq_track_1/sky130_fd_sc_hs__fa_2_15/B fine_freq_track_1/sky130_fd_sc_hs__dfxtp_2_5/a_431_508#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_83/a_812_138# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_21/a_850_127#
+ fine_freq_track_1/sky130_fd_sc_hs__a22oi_1_3/a_159_74# fine_freq_track_1/sky130_fd_sc_hs__o21a_1_17/a_320_74#
+ fine_freq_track_1/sky130_fd_sc_hs__inv_4_33/Y fine_freq_track_1/sky130_fd_sc_hs__xnor2_1_3/a_138_385#
+ fine_freq_track_1/sky130_fd_sc_hs__nand3_1_1/A fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_23/a_1827_81#
+ fine_freq_track_1/sky130_fd_sc_hs__a21oi_1_49/a_29_368# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_29/a_714_127#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_3/D fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_71/a_124_78#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_9/a_832_118# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_27/a_1224_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_73/a_1350_392# fine_freq_track_1/sky130_fd_sc_hs__nor2_1_99/Y
+ fine_freq_track_1/sky130_fd_sc_hs__o21a_1_61/a_320_74# fine_freq_track_1/sky130_fd_sc_hs__a21oi_1_17/a_29_368#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_21/a_796_463# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_19/a_38_78#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_45/a_1547_508# fine_freq_track_1/sky130_fd_sc_hs__o21a_1_17/X
+ fine_freq_track_1/sky130_fd_sc_hs__inv_4_83/Y fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_33/a_1627_493#
+ fine_freq_track_1/sky130_fd_sc_hs__inv_4_61/A fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_31/D
+ fine_freq_track_1/sky130_fd_sc_hs__xnor2_1_13/A fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_43/a_706_463#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_35/a_319_360# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_9/a_834_355#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_89/a_1678_395# fine_freq_track_1/sky130_fd_sc_hs__fa_2_11/a_27_378#
+ fine_freq_track_1/sky130_fd_sc_hs__a21oi_1_61/a_29_368# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_23/a_1350_392#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_59/a_494_366# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_79/a_37_78#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_13/a_1434_74# fine_freq_track_1/sky130_fd_sc_hs__maj3_1_1/a_598_384#
+ fine_freq_track_1/sky130_fd_sc_hs__and2_2_5/X fine_freq_track_1/sky130_fd_sc_hs__o21a_1_17/A1
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_39/a_1482_48# fine_freq_track_1/sky130_fd_sc_hs__fa_2_3/A
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_37/a_1678_395# fine_freq_track_1/sky130_fd_sc_hs__o22ai_1_7/A1
+ fine_freq_track_1/sky130_fd_sc_hs__nor3_1_15/A fine_freq_track_1/sky130_fd_sc_hs__fa_2_21/CIN
+ fine_freq_track_1/sky130_fd_sc_hs__a21oi_1_79/a_117_74# fine_freq_track_1/sky130_fd_sc_hs__fa_2_19/B
+ fine_freq_track_1/sky130_fd_sc_hs__dfxtp_4_5/a_544_485# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_7/a_38_78#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_27/a_120_74# fine_freq_track_1/sky130_fd_sc_hs__nand2_2_1/B
+ fine_freq_track_1/sky130_fd_sc_hs__a21oi_1_47/a_117_74# fine_freq_track_1/sky130_fd_sc_hs__o21a_1_33/X
+ fine_freq_track_1/sky130_fd_sc_hs__inv_4_25/A fine_freq_track_1/sky130_fd_sc_hs__fa_2_11/a_701_79#
+ fine_freq_track_1/sky130_fd_sc_hs__a32oi_1_7/a_469_74# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_31/a_699_463#
+ fine_freq_track_1/sky130_fd_sc_hs__xnor2_1_11/a_138_385# fine_freq_track_1/sky130_fd_sc_hs__a21oi_1_91/a_117_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_23/a_37_78# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_21/a_300_74#
+ fine_freq_track_1/sky130_fd_sc_hs__nor2_1_117/a_116_368# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_7/Q
+ fine_freq_track_1/sky130_fd_sc_hs__a211oi_1_1/a_159_74# fine_freq_track_1/sky130_fd_sc_hs__dfxtp_4_3/a_27_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_63/a_313_74# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_33/a_841_401#
+ fine_freq_track_1/sky130_fd_sc_hs__o21a_1_63/X fine_freq_track_1/sky130_fd_sc_hs__o21a_1_63/A2
+ fine_freq_track_1/sky130_fd_sc_hs__nand2_1_107/a_117_74# fine_freq_track_1/sky130_fd_sc_hs__nor2_1_33/Y
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_39/a_1934_94# fine_freq_track_1/sky130_fd_sc_hs__xnor2_1_1/a_376_368#
+ fine_freq_track_1/sky130_fd_sc_hs__nor2b_1_47/a_278_368# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_1/a_120_74#
+ fine_freq_track_1/sky130_fd_sc_hs__inv_2_3/A fine_freq_track_1/sky130_fd_sc_hs__nand4_1_5/A
+ fine_freq_track_1/sky130_fd_sc_hs__o21a_1_37/a_83_244# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_31/a_313_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_9/a_812_138# fine_freq_track_1/sky130_fd_sc_hs__nor2_1_7/B
+ fine_freq_track_1/sky130_fd_sc_hs__nand4_1_1/C fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_11/a_856_304#
+ fine_freq_track_1/sky130_fd_sc_hs__inv_4_123/Y fine_freq_track_1/sky130_fd_sc_hs__o21a_1_71/B1
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_11/a_850_127# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_83/a_1627_493#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_31/a_125_78# fine_freq_track_1/sky130_fd_sc_hs__nor2b_1_19/Y
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_17/a_1647_81# fine_freq_track_1/sky130_fd_sc_hs__fa_2_5/a_1119_79#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_13/a_1827_81# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_9/a_1547_508#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_19/a_714_127# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_57/a_1647_81#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_17/a_1224_74# fine_freq_track_1/sky130_fd_sc_hs__inv_4_19/A
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_1/Q_N fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_9/a_2010_409#
+ fine_freq_track_1/sky130_fd_sc_hs__nor2_1_57/Y fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_3/a_817_508#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_11/a_796_463# fine_freq_track_1/sky130_fd_sc_hs__fa_2_9/SUM
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_43/a_789_463# fine_freq_track_1/sky130_fd_sc_hs__o22ai_1_9/Y
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_91/a_1827_81# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_37/a_498_360#
+ fine_freq_track_1/sky130_fd_sc_hs__nor2b_2_1/Y fine_freq_track_1/sky130_fd_sc_hs__nor3_1_3/Y
+ fine_freq_track_1/sky130_fd_sc_hs__xor2_1_7/a_158_392# fine_freq_track_1/sky130_fd_sc_hs__a22oi_1_7/a_159_74#
+ fine_freq_track_1/sky130_fd_sc_hs__nand2_2_5/a_27_74# fine_freq_track_1/sky130_fd_sc_hs__nor2_1_69/B
+ fine_freq_track_1/sky130_fd_sc_hs__o21ai_1_3/Y fine_freq_track_1/sky130_fd_sc_hs__nor2_1_5/B
+ fine_freq_track_1/sky130_fd_sc_hs__nand3_1_1/B fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_41/D
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_21/a_1350_392# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_75/a_124_78#
+ fine_freq_track_1/sky130_fd_sc_hs__inv_4_41/A fine_freq_track_1/sky130_fd_sc_hs__fa_2_5/SUM
+ fine_freq_track_1/sky130_fd_sc_hs__o21a_1_27/A1 fine_freq_track_1/sky130_fd_sc_hs__nor2_1_99/A
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_7/a_1598_93# fine_freq_track_1/sky130_fd_sc_hs__o21a_1_65/a_320_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_9/a_841_401# fine_freq_track_1/sky130_fd_sc_hs__a22oi_1_1/a_339_74#
+ fine_freq_track_1/sky130_fd_sc_hs__fa_2_23/B fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_1/a_1624_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfxtp_4_2/a_206_368# fine_freq_track_1/sky130_fd_sc_hs__sdlclkp_4_1/a_1292_74#
+ fine_freq_track_1/sky130_fd_sc_hs__o21a_1_17/a_376_387# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_21/a_1465_471#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_17/a_890_138# fine_freq_track_1/sky130_fd_sc_hs__a21oi_1_65/a_29_368#
+ fine_freq_track_1/sky130_fd_sc_hs__or2_1_1/X fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_39/a_1465_471#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_57/a_890_138# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_47/a_37_78#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_9/a_507_368# fine_freq_track_1/sky130_fd_sc_hs__fa_2_3/a_336_347#
+ fine_freq_track_1/sky130_fd_sc_hs__inv_4_29/A fine_freq_track_1/sky130_fd_sc_hs__nand2_2_5/B
+ fine_freq_track_1/sky130_fd_sc_hs__o21a_1_3/A1 fine_freq_track_1/sky130_fd_sc_hs__dfstp_2_5/a_1566_92#
+ fine_freq_track_1/sky130_fd_sc_hs__nor4_1_1/A fine_freq_track_1/sky130_fd_sc_hs__nand4_2_1/a_304_74#
+ fine_freq_track_1/sky130_fd_sc_hs__nor2_1_21/Y fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_31/a_910_118#
+ fine_freq_track_1/sky130_fd_sc_hs__a32oi_1_1/a_391_74# fine_freq_track_1/sky130_fd_sc_hs__maj3_1_3/C
+ fine_freq_track_1/sky130_fd_sc_hs__nor2_1_63/Y fine_freq_track_1/sky130_fd_sc_hs__inv_4_91/A
+ fine_freq_track_1/sky130_fd_sc_hs__nor2_1_61/a_116_368# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_33/a_1550_119#
+ fine_freq_track_1/sky130_fd_sc_hs__nor2b_1_3/a_278_368# fine_freq_track_1/sky130_fd_sc_hs__fa_2_9/B
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_3/a_498_360# fine_freq_track_1/sky130_fd_sc_hs__nor3_1_9/C
+ fine_freq_track_1/sky130_fd_sc_hs__nor2_1_73/Y fine_freq_track_1/sky130_fd_sc_hs__o31ai_1_3/a_114_74#
+ fine_freq_track_1/sky130_fd_sc_hs__inv_4_109/A fine_freq_track_1/sky130_fd_sc_hs__a22o_1_23/a_132_392#
+ fine_freq_track_1/sky130_fd_sc_hs__fa_2_5/CIN fine_freq_track_1/sky130_fd_sc_hs__inv_4_39/Y
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_29/a_1934_94# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_25/a_1624_74#
+ fine_freq_track_1/sky130_fd_sc_hs__fa_2_15/a_992_347# fine_freq_track_1/sky130_fd_sc_hs__nor2b_1_37/a_278_368#
+ fine_freq_track_1/sky130_fd_sc_hs__dfxtp_2_7/a_708_101# fine_freq_track_1/sky130_fd_sc_hs__a21oi_1_95/a_117_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfxtp_4_5/D fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_7/a_1547_508#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_67/a_313_74# fine_freq_track_1/sky130_fd_sc_hs__xnor2_1_5/Y
+ fine_freq_track_1/sky130_fd_sc_hs__nand2_1_89/Y fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_43/a_120_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_49/a_714_127# fine_freq_track_1/sky130_fd_sc_hs__o31ai_1_3/Y
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_43/a_1547_508# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_35/a_313_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_9/a_2026_424# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_33/a_789_463#
+ fine_freq_track_1/sky130_fd_sc_hs__o21a_1_1/A1 fine_freq_track_1/sky130_fd_sc_hs__nand4_1_1/D
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_81/a_1827_81# fine_freq_track_1/sky130_fd_sc_hs__xor2_1_5/a_355_368#
+ fine_freq_track_1/sky130_fd_sc_hs__inv_2_5/A fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_31/a_1627_493#
+ fine_freq_track_1/sky130_fd_sc_hs__inv_4_99/A fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_7/a_910_118#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_35/a_125_78# fine_freq_track_1/sky130_fd_sc_hs__o21a_1_25/X
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_23/a_706_463# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_87/a_1678_395#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_49/a_1627_493# fine_freq_track_1/sky130_fd_sc_hs__a21oi_1_111/a_29_368#
+ fine_freq_track_1/sky130_fd_sc_hs__inv_4_89/Y fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_19/a_1736_119#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_39/a_494_366# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_19/a_1266_119#
+ fine_freq_track_1/sky130_fd_sc_hs__o21a_1_53/a_83_244# fine_freq_track_1/sky130_fd_sc_hs__inv_4_23/A
+ fine_freq_track_1/sky130_fd_sc_hs__o21a_1_61/A2 fine_freq_track_1/sky130_fd_sc_hs__o21a_1_59/A2
+ fine_freq_track_1/sky130_fd_sc_hs__inv_4_117/Y fine_freq_track_1/sky130_fd_sc_hs__o21ai_1_11/Y
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_33/a_1434_74# fine_freq_track_1/sky130_fd_sc_hs__nor2_1_49/Y
+ fine_freq_track_1/sky130_fd_sc_hs__fa_2_17/a_27_79# fine_freq_track_1/sky130_fd_sc_hs__nor3_1_13/B
+ fine_freq_track_1/sky130_fd_sc_hs__nand3_1_1/C fine_freq_track_1/sky130_fd_sc_hs__xnor2_1_9/Y
+ fine_freq_track_1/sky130_fd_sc_hs__dfxtp_4_2/a_437_503# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_51/a_2010_409#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_41/a_832_118# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_79/a_124_78#
+ fine_freq_track_1/sky130_fd_sc_hs__nor2b_1_21/a_27_112# fine_freq_track_1/sky130_fd_sc_hs__nor2_1_99/B
+ fine_freq_track_1/sky130_fd_sc_hs__o21a_1_75/A2 fine_freq_track_1/sky130_fd_sc_hs__nand2_1_53/a_117_74#
+ fine_freq_track_1/sky130_fd_sc_hs__o21a_1_69/a_320_74# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_27/a_38_78#
+ fine_freq_track_1/sky130_fd_sc_hs__o21a_1_9/X fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_21/a_910_118#
+ fine_freq_track_1/sky130_fd_sc_hs__inv_4_69/Y fine_freq_track_1/sky130_fd_sc_hs__nor3_1_5/a_114_368#
+ fine_freq_track_1/sky130_fd_sc_hs__o21a_1_35/a_320_74# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_11/a_699_463#
+ fine_freq_track_1/sky130_fd_sc_hs__nor2_1_51/a_116_368# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_31/a_1550_119#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_13/a_124_78# fine_freq_track_1/sky130_fd_sc_hs__fa_2_19/a_27_378#
+ fine_freq_track_1/sky130_fd_sc_hs__a21oi_1_69/a_29_368# fine_freq_track_1/sky130_fd_sc_hs__inv_4_133/A
+ fine_freq_track_1/sky130_fd_sc_hs__a22oi_1_21/a_71_368# fine_freq_track_1/sky130_fd_sc_hs__nand2b_1_3/a_27_112#
+ fine_freq_track_1/sky130_fd_sc_hs__o21a_1_7/X fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_19/a_2010_409#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_19/a_1934_94# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_15/a_1624_74#
+ fine_freq_track_1/sky130_fd_sc_hs__a21oi_1_35/a_29_368# fine_freq_track_1/sky130_fd_sc_hs__nor2b_1_27/a_278_368#
+ fine_freq_track_1/sky130_fd_sc_hs__nor2_1_1/Y fine_freq_track_1/sky130_fd_sc_hs__nor4_1_1/B
+ fine_freq_track_1/sky130_fd_sc_hs__a32oi_1_5/a_391_74# fine_freq_track_1/sky130_fd_sc_hs__fa_2_15/SUM
+ fine_freq_track_1/sky130_fd_sc_hs__nand2_1_71/Y fine_freq_track_1/sky130_fd_sc_hs__o21a_1_71/X
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_81/a_1627_493# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_9/a_1434_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_29/a_33_74# fine_freq_track_1/sky130_fd_sc_hs__inv_4_71/A
+ fine_freq_track_1/sky130_fd_sc_hs__nor2_1_101/Y fine_freq_track_1/sky130_fd_sc_hs__o21a_1_9/B1
+ fine_freq_track_1/sky130_fd_sc_hs__sdlclkp_1_1/a_1166_94# fine_freq_track_1/sky130_fd_sc_hs__inv_2_3/Y
+ fine_freq_track_1/sky130_fd_sc_hs__o31ai_1_7/a_114_74# fine_freq_track_1/sky130_fd_sc_hs__a32oi_1_1/a_27_368#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_71/a_1350_392# fine_freq_track_1/sky130_fd_sc_hs__o31ai_1_1/Y
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_7/a_1827_81# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_7/a_2010_409#
+ fine_freq_track_1/sky130_fd_sc_hs__o21a_1_19/X fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_37/a_1224_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_41/a_1547_508# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_23/a_789_463#
+ fine_freq_track_1/sky130_fd_sc_hs__fa_2_19/a_701_79# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_71/a_1827_81#
+ fine_freq_track_1/sky130_fd_sc_hs__o31ai_1_7/Y fine_freq_track_1/sky130_fd_sc_hs__a22oi_1_23/Y
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_7/a_313_74# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_13/a_706_463#
+ fine_freq_track_1/sky130_fd_sc_hs__a22o_1_25/a_222_392# fine_freq_track_1/sky130_fd_sc_hs__a21oi_1_99/a_117_74#
+ fine_freq_track_1/sky130_fd_sc_hs__inv_4_89/A fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_29/a_300_74#
+ fine_freq_track_1/sky130_fd_sc_hs__inv_4_7/Y fine_freq_track_1/sky130_fd_sc_hs__inv_4_51/Y
+ fine_freq_track_1/sky130_fd_sc_hs__nand2_1_91/A fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_43/a_319_360#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_29/a_494_366# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_43/a_834_355#
+ fine_freq_track_1/sky130_fd_sc_hs__o21a_1_7/A2 fine_freq_track_1/sky130_fd_sc_hs__xor2_1_9/a_194_125#
+ fine_freq_track_1/sky130_fd_sc_hs__nor3_1_15/a_198_368# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_67/a_494_366#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_39/a_1350_392# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_39/a_313_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfstp_2_1/a_781_74# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_13/a_120_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_47/a_922_127# fine_freq_track_1/sky130_fd_sc_hs__o21a_1_75/A1
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_45/a_33_74# fine_freq_track_1/sky130_fd_sc_hs__inv_4_97/A
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_9/a_856_304# fine_freq_track_1/sky130_fd_sc_hs__fa_2_5/B
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_35/a_1678_395# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_9/a_850_127#
+ fine_freq_track_1/sky130_fd_sc_hs__inv_4_99/Y fine_freq_track_1/sky130_fd_sc_hs__inv_4_1/A
+ fine_freq_track_1/sky130_fd_sc_hs__xnor2_1_11/Y fine_freq_track_1/sky130_fd_sc_hs__o21a_1_35/a_376_387#
+ fine_freq_track_1/sky130_fd_sc_hs__a21oi_1_115/a_29_368# fine_freq_track_1/sky130_fd_sc_hs__inv_4_75/Y
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_83/a_313_74# fine_freq_track_1/sky130_fd_sc_hs__inv_4_15/Y
+ fine_freq_track_1/sky130_fd_sc_hs__o31ai_1_1/A3 fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_19/D
+ fine_freq_track_1/sky130_fd_sc_hs__o21a_1_75/a_376_387# fine_freq_track_1/sky130_fd_sc_hs__o21a_1_57/a_83_244#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_69/a_2010_409# fine_freq_track_1/sky130_fd_sc_hs__nand2_2_7/Y
+ fine_freq_track_1/sky130_fd_sc_hs__xnor2_1_7/B fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_11/a_910_118#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_45/a_817_508# fine_freq_track_1/sky130_fd_sc_hs__fa_2_15/a_487_79#
+ fine_freq_track_1/sky130_fd_sc_hs__inv_4_13/Y fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_3/a_1224_74#
+ fine_freq_track_1/sky130_fd_sc_hs__o21a_1_57/X fine_freq_track_1/sky130_fd_sc_hs__dfstp_2_7/a_1356_74#
+ fine_freq_track_1/sky130_fd_sc_hs__nor2b_1_25/a_27_112# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_17/a_2010_409#
+ fine_freq_track_1/sky130_fd_sc_hs__inv_4_107/Y fine_freq_track_1/sky130_fd_sc_hs__nor2b_1_17/a_278_368#
+ fine_freq_track_1/sky130_fd_sc_hs__nand2_1_57/a_117_74# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_41/a_841_401#
+ fine_freq_track_1/sky130_fd_sc_hs__nand2_2_13/Y fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_49/a_124_78#
+ fine_freq_track_1/sky130_fd_sc_hs__a22o_1_1/a_222_392# fine_freq_track_1/sky130_fd_sc_hs__a22oi_1_9/a_339_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_49/a_1934_94# fine_freq_track_1/sky130_fd_sc_hs__o21a_1_1/X
+ fine_freq_track_1/sky130_fd_sc_hs__fa_2_1/SUM fine_freq_track_1/sky130_fd_sc_hs__nand3_1_1/a_233_74#
+ fine_freq_track_1/sky130_fd_sc_hs__o21a_1_49/X fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_43/a_812_138#
+ fine_freq_track_1/sky130_fd_sc_hs__dfxtp_2_3/a_431_508# fine_freq_track_1/sky130_fd_sc_hs__o21a_1_67/A2
+ fine_freq_track_1/sky130_fd_sc_hs__o211ai_1_9/C1 fine_freq_track_1/sky130_fd_sc_hs__a22oi_1_25/a_71_368#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_27/a_1647_81# fine_freq_track_1/sky130_fd_sc_hs__nand2b_1_7/a_27_112#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_57/a_37_78# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_21/a_1827_81#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_61/a_124_78# fine_freq_track_1/sky130_fd_sc_hs__dfxtp_2_1/a_695_459#
+ fine_freq_track_1/sky130_fd_sc_hs__xor2_1_1/X fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_13/a_789_463#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_7/a_2026_424# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_61/a_1827_81#
+ fine_freq_track_1/sky130_fd_sc_hs__a32oi_1_9/a_391_74# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_89/a_1350_392#
+ fine_freq_track_1/sky130_fd_sc_hs__o21a_1_51/a_320_74# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_45/a_498_360#
+ fine_freq_track_1/sky130_fd_sc_hs__a22o_1_15/a_222_392# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_91/a_789_463#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_85/a_1678_395# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_47/a_1627_493#
+ fine_freq_track_1/sky130_fd_sc_hs__conb_1_1/HI fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_3/a_33_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_17/a_1736_119# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_33/a_834_355#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_19/a_494_366# fine_freq_track_1/sky130_fd_sc_hs__o21a_1_31/X
+ fine_freq_track_1/sky130_fd_sc_hs__a32oi_1_5/a_27_368# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_17/a_1266_119#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_37/a_1350_392# fine_freq_track_1/sky130_fd_sc_hs__o21a_1_57/B1
+ fine_freq_track_1/sky130_fd_sc_hs__inv_4_135/A fine_freq_track_1/sky130_fd_sc_hs__inv_4_113/A
+ fine_freq_track_1/sky130_fd_sc_hs__o22ai_1_5/a_27_74# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_27/a_890_138#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_37/a_1465_471# fine_freq_track_1/sky130_fd_sc_hs__inv_4_31/Y
+ fine_freq_track_1/sky130_fd_sc_hs__o211ai_1_1/a_31_74# fine_freq_track_1/sky130_fd_sc_hs__o22ai_1_1/A2
+ fine_freq_track_1/sky130_fd_sc_hs__dfxtp_4_3/a_651_503# fine_freq_track_1/sky130_fd_sc_hs__o21a_1_65/a_376_387#
+ fine_freq_track_1/sky130_fd_sc_hs__o21a_1_77/B1 fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_67/a_2010_409#
+ fine_freq_track_1/sky130_fd_sc_hs__o21a_1_9/A1 fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_5/Q_N
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_17/a_120_74# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_35/a_817_508#
+ fine_freq_track_1/sky130_fd_sc_hs__nor2b_1_33/Y fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_13/a_33_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfxtp_2_9/a_27_74# fine_freq_track_1/sky130_fd_sc_hs__nor2_1_31/a_116_368#
+ fine_freq_track_1/sky130_fd_sc_hs__o21a_1_1/a_83_244# fine_freq_track_1/sky130_fd_sc_hs__o21a_1_21/X
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_45/a_300_74# fine_freq_track_1/sky130_fd_sc_hs__nor2_1_75/B
+ fine_freq_track_1/sky130_fd_sc_hs__nand2_1_91/B fine_freq_track_1/sky130_fd_sc_hs__o21a_1_61/X
+ fine_freq_track_1/sky130_fd_sc_hs__nor2_2_1/a_35_368# fine_freq_track_1/sky130_fd_sc_hs__a21oi_1_119/a_29_368#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_5/a_699_463# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_7/a_300_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_87/a_313_74# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_49/a_1550_119#
+ fine_freq_track_1/sky130_fd_sc_hs__nor2b_1_41/A fine_freq_track_1/sky130_fd_sc_hs__inv_4_5/Y
+ fine_freq_track_1/sky130_fd_sc_hs__fa_2_9/a_484_347# fine_freq_track_1/sky130_fd_sc_hs__a21oi_1_82/a_117_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_11/a_300_74# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_53/a_313_74#
+ fine_freq_track_1/sky130_fd_sc_hs__fa_2_23/a_336_347# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_35/a_1624_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_5/a_922_127# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_39/a_1598_93#
+ fine_freq_track_1/sky130_fd_sc_hs__o21a_1_27/a_83_244# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_33/a_812_138#
+ fine_freq_track_1/sky130_fd_sc_hs__fa_2_3/a_27_79# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_21/a_125_78#
+ fine_freq_track_1/sky130_fd_sc_hs__fa_2_19/a_484_347# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_5/a_1547_508#
+ fine_freq_track_1/sky130_fd_sc_hs__nor2b_1_29/a_27_112# fine_freq_track_1/sky130_fd_sc_hs__nor2b_1_1/a_27_112#
+ fine_freq_track_1/sky130_fd_sc_hs__a22o_1_25/a_230_79# fine_freq_track_1/sky130_fd_sc_hs__nor4_1_3/C
+ fine_freq_track_1/sky130_fd_sc_hs__nor2_2_3/Y fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_5/a_1482_48#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_5/a_2010_409# fine_freq_track_1/sky130_fd_sc_hs__o2bb2ai_1_1/a_114_74#
+ fine_freq_track_1/sky130_fd_sc_hs__fa_2_7/CIN fine_freq_track_1/sky130_fd_sc_hs__o21ai_1_1/Y
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_37/a_38_78# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_51/a_1827_81#
+ fine_freq_track_1/sky130_fd_sc_hs__nand2_4_5/Y fine_freq_track_1/sky130_fd_sc_hs__inv_4_37/Y
+ fine_freq_track_1/sky130_fd_sc_hs__inv_4_17/A fine_freq_track_1/sky130_fd_sc_hs__o21ai_1_5/B1
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_1/a_817_508# fine_freq_track_1/sky130_fd_sc_hs__inv_4_35/A
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_1/a_124_78# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_31/D
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_81/a_789_463# fine_freq_track_1/sky130_fd_sc_hs__fa_2_13/SUM
+ fine_freq_track_1/sky130_fd_sc_hs__a222oi_1_1/Y fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_33/a_706_463#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_23/a_319_360# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_23/a_834_355#
+ fine_freq_track_1/sky130_fd_sc_hs__fa_2_15/a_1119_79# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_25/a_37_78#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_65/a_124_78# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_47/a_494_366#
+ fine_freq_track_1/sky130_fd_sc_hs__dfxtp_4_5/a_27_74# fine_freq_track_1/sky130_fd_sc_hs__dfxtp_4_9/a_1178_124#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_27/a_922_127# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_87/a_494_366#
+ fine_freq_track_1/sky130_fd_sc_hs__o211ai_1_7/a_116_368# fine_freq_track_1/sky130_fd_sc_hs__o21a_1_55/a_320_74#
+ fine_freq_track_1/sky130_fd_sc_hs__a222o_1_1/X fine_freq_track_1/sky130_fd_sc_hs__a32oi_1_1/a_119_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_41/a_1434_74# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_33/a_1678_395#
+ fine_freq_track_1/sky130_fd_sc_hs__o21a_1_21/A1 fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_29/a_1482_48#
+ fine_freq_track_1/sky130_fd_sc_hs__inv_4_127/A fine_freq_track_1/sky130_fd_sc_hs__xnor2_1_1/a_112_119#
+ fine_freq_track_1/sky130_fd_sc_hs__nor2b_1_21/Y fine_freq_track_1/sky130_fd_sc_hs__a22oi_1_5/a_71_368#
+ fine_freq_track_1/sky130_fd_sc_hs__o21a_1_55/a_376_387# fine_freq_track_1/sky130_fd_sc_hs__a21oi_1_55/a_29_368#
+ fine_freq_track_1/sky130_fd_sc_hs__a32oi_1_9/a_27_368# fine_freq_track_1/sky130_fd_sc_hs__nor2_1_61/Y
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_7/a_507_368# fine_freq_track_1/sky130_fd_sc_hs__fa_2_3/a_992_347#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_25/a_817_508# fine_freq_track_1/sky130_fd_sc_hs__dfstp_2_4/a_1566_92#
+ fine_freq_track_1/sky130_fd_sc_hs__nor2_1_95/A fine_freq_track_1/sky130_fd_sc_hs__nor2_1_65/A
+ fine_freq_track_1/sky130_fd_sc_hs__nor2_1_21/a_116_368# fine_freq_track_1/sky130_fd_sc_hs__o21a_1_1/a_376_387#
+ fine_freq_track_1/sky130_fd_sc_hs__nor2_1_3/Y fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_41/a_37_78#
+ fine_freq_track_1/sky130_fd_sc_hs__nor2_1_21/B fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_1/a_498_360#
+ fine_freq_track_1/sky130_fd_sc_hs__nand2_2_9/a_27_74# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_47/a_1550_119#
+ fine_freq_track_1/sky130_fd_sc_hs__sdlclkp_4_1/a_116_395# fine_freq_track_1/sky130_fd_sc_hs__a22oi_1_1/Y
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_15/a_2010_409# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_9/a_706_463#
+ fine_freq_track_1/sky130_fd_sc_hs__a22o_1_21/a_132_392# fine_freq_track_1/sky130_fd_sc_hs__fa_2_13/a_336_347#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_29/a_1598_93# fine_freq_track_1/sky130_fd_sc_hs__nor2b_1_35/a_278_368#
+ fine_freq_track_1/sky130_fd_sc_hs__inv_2_7/A fine_freq_track_1/sky130_fd_sc_hs__xnor2_1_1/a_293_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_23/a_812_138# fine_freq_track_1/sky130_fd_sc_hs__o21a_1_5/a_83_244#
+ fine_freq_track_1/sky130_fd_sc_hs__dfstp_2_5/a_716_456# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_49/a_300_74#
+ fine_freq_track_1/sky130_fd_sc_hs__o21a_1_53/X fine_freq_track_1/sky130_fd_sc_hs__nor2_1_49/B
+ fine_freq_track_1/sky130_fd_sc_hs__and2_2_1/a_31_74# fine_freq_track_1/sky130_fd_sc_hs__inv_4_1/Y
+ fine_freq_track_1/sky130_fd_sc_hs__nand2_1_67/Y fine_freq_track_1/sky130_fd_sc_hs__a21oi_1_85/a_117_74#
+ fine_freq_track_1/sky130_fd_sc_hs__fa_2_15/CIN fine_freq_track_1/sky130_fd_sc_hs__inv_2_9/A
+ fine_freq_track_1/sky130_fd_sc_hs__fa_2_5/a_683_347# fine_freq_track_1/sky130_fd_sc_hs__fa_2_23/CIN
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_33/a_120_74# fine_freq_track_1/sky130_fd_sc_hs__inv_4_51/A
+ fine_freq_track_1/sky130_fd_sc_hs__a21oi_1_51/a_117_74# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_41/a_1827_81#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_47/a_714_127# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_87/a_1350_392#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_85/a_1647_81# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_45/a_1224_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_7/a_789_463# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_25/a_498_360#
+ fine_freq_track_1/sky130_fd_sc_hs__fa_2_13/CIN fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_71/a_789_463#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_83/a_1678_395# fine_freq_track_1/sky130_fd_sc_hs__a222oi_1_1/a_116_392#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_31/Q_N fine_freq_track_1/sky130_fd_sc_hs__dfxtp_2_9/a_644_504#
+ fine_freq_track_1/sky130_fd_sc_hs__a22o_1_27/X fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_13/a_319_360#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_13/a_834_355# fine_freq_track_1/sky130_fd_sc_hs__a21oi_1_101/a_29_368#
+ fine_freq_track_1/sky130_fd_sc_hs__a22o_1_29/a_230_79# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_37/a_494_366#
+ fine_freq_track_1/sky130_fd_sc_hs__nand2_1_111/a_117_74# fine_freq_track_1/sky130_fd_sc_hs__a21oi_1_1/a_117_74#
+ fine_freq_track_1/sky130_fd_sc_hs__sdlclkp_4_1/a_792_48# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_3/a_494_366#
+ fine_freq_track_1/sky130_fd_sc_hs__inv_4_53/A fine_freq_track_1/sky130_fd_sc_hs__o21ai_1_5/a_162_368#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_17/a_922_127# fine_freq_track_1/sky130_fd_sc_hs__o21a_1_43/a_83_244#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_77/a_494_366# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_91/a_834_355#
+ fine_freq_track_1/sky130_fd_sc_hs__dfxtp_2_11/a_206_368# fine_freq_track_1/sky130_fd_sc_hs__nor2_1_91/Y
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_33/D fine_freq_track_1/sky130_fd_sc_hs__a21oi_1_19/Y
+ fine_freq_track_1/sky130_fd_sc_hs__nand2_4_5/a_27_74# fine_freq_track_1/sky130_fd_sc_hs__a22o_1_9/a_132_392#
+ fine_freq_track_1/sky130_fd_sc_hs__dfxtp_2_11/a_1125_508# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_19/a_1482_48#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_35/a_1465_471# fine_freq_track_1/sky130_fd_sc_hs__o21a_1_45/a_376_387#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_69/a_124_78# fine_freq_track_1/sky130_fd_sc_hs__nor2b_1_11/a_27_112#
+ fine_freq_track_1/sky130_fd_sc_hs__nor2b_1_29/Y fine_freq_track_1/sky130_fd_sc_hs__nor2_1_51/B
+ fine_freq_track_1/sky130_fd_sc_hs__nand2_4_7/A fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_85/a_890_138#
+ fine_freq_track_1/sky130_fd_sc_hs__o21a_1_59/a_320_74# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_15/a_817_508#
+ fine_freq_track_1/sky130_fd_sc_hs__a32oi_1_5/a_119_74# fine_freq_track_1/sky130_fd_sc_hs__dfxtp_4_9/a_735_102#
+ fine_freq_track_1/sky130_fd_sc_hs__nor2_1_11/a_116_368# fine_freq_track_1/sky130_fd_sc_hs__o21a_1_71/A2
+ fine_freq_track_1/sky130_fd_sc_hs__o211ai_1_5/a_311_74# fine_freq_track_1/sky130_fd_sc_hs__conb_1_1/LO
+ fine_freq_track_1/sky130_fd_sc_hs__fa_2_21/SUM fine_freq_track_1/sky130_fd_sc_hs__nor2b_1_13/Y
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_19/a_2026_424# fine_freq_track_1/sky130_fd_sc_hs__a21oi_1_59/a_29_368#
+ fine_freq_track_1/sky130_fd_sc_hs__nor2_1_23/Y fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_21/a_38_78#
+ fine_freq_track_1/sky130_fd_sc_hs__a22oi_1_11/a_71_368# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_19/a_1598_93#
+ fine_freq_track_1/sky130_fd_sc_hs__inv_4_67/A fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_13/a_812_138#
+ fine_freq_track_1/sky130_fd_sc_hs__inv_4_3/Y fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_29/D
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_81/a_37_78# fine_freq_track_1/sky130_fd_sc_hs__fa_2_21/a_27_378#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_3/a_1547_508# fine_freq_track_1/sky130_fd_sc_hs__xnor2_1_9/B
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_91/a_812_138# fine_freq_track_1/sky130_fd_sc_hs__fa_2_9/a_1205_79#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_1/a_1647_81# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_5/a_2026_424#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_31/a_1827_81# fine_freq_track_1/sky130_fd_sc_hs__xnor2_1_5/a_293_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_75/a_1647_81# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_21/a_789_463#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_23/a_33_74# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_15/a_498_360#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_39/a_796_463# fine_freq_track_1/sky130_fd_sc_hs__fa_2_1/A
+ fine_freq_track_1/sky130_fd_sc_hs__a22o_1_25/a_52_123# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_61/a_789_463#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_45/a_1627_493# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_15/a_1736_119#
+ fine_freq_track_1/sky130_fd_sc_hs__maj3_1_1/X fine_freq_track_1/sky130_fd_sc_hs__a21oi_1_89/a_117_74#
+ fine_freq_track_1/sky130_fd_sc_hs__xor2_1_11/a_355_368# fine_freq_track_1/sky130_fd_sc_hs__a222oi_1_3/a_461_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_19/a_300_74# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_15/a_1266_119#
+ fine_freq_track_1/sky130_fd_sc_hs__fa_2_19/a_1205_79# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_1/Q
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_35/a_1350_392# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_37/a_120_74#
+ fine_freq_track_1/sky130_fd_sc_hs__inv_4_81/A fine_freq_track_1/sky130_fd_sc_hs__xor2_1_7/a_194_125#
+ fine_freq_track_1/sky130_fd_sc_hs__dfxtp_4_7/a_1178_124# fine_freq_track_1/sky130_fd_sc_hs__nor2_1_15/Y
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_81/a_834_355# fine_freq_track_1/sky130_fd_sc_hs__o21a_1_23/X
+ fine_freq_track_1/sky130_fd_sc_hs__fa_2_21/a_701_79# fine_freq_track_1/sky130_fd_sc_hs__inv_4_97/Y
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_29/a_313_74# fine_freq_track_1/sky130_fd_sc_hs__xnor2_1_7/A
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_31/a_1678_395# fine_freq_track_1/sky130_fd_sc_hs__a21oi_1_23/a_117_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_7/a_856_304# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_29/a_125_78#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_7/a_850_127# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_49/a_1678_395#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_47/a_1482_48# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_3/a_125_78#
+ fine_freq_track_1/sky130_fd_sc_hs__o21ai_1_9/a_27_74# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_31/a_832_118#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_65/a_2010_409# fine_freq_track_1/sky130_fd_sc_hs__a21oi_1_5/a_117_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_1/a_890_138# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_45/a_38_78#
+ fine_freq_track_1/sky130_fd_sc_hs__sdlclkp_4_1/a_324_79# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_5/a_714_127#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_75/a_890_138# fine_freq_track_1/sky130_fd_sc_hs__fa_2_17/CIN
+ fine_freq_track_1/sky130_fd_sc_hs__o21a_1_47/a_83_244# fine_freq_track_1/sky130_fd_sc_hs__a22o_1_1/a_230_79#
+ fine_freq_track_1/sky130_fd_sc_hs__o21a_1_13/a_83_244# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_1/a_1224_74#
+ fine_freq_track_1/sky130_fd_sc_hs__o21a_1_3/a_320_74# fine_freq_track_1/sky130_fd_sc_hs__nor2_1_43/B
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_17/a_2026_424# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_49/a_699_463#
+ fine_freq_track_1/sky130_fd_sc_hs__or3b_2_1/C_N fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_35/a_37_78#
+ fine_freq_track_1/sky130_fd_sc_hs__and2_2_1/a_118_74# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_89/a_699_463#
+ fine_freq_track_1/sky130_fd_sc_hs__nor2b_1_15/a_27_112# fine_freq_track_1/sky130_fd_sc_hs__inv_4_35/Y
+ fine_freq_track_1/sky130_fd_sc_hs__o21a_1_47/X fine_freq_track_1/sky130_fd_sc_hs__a22o_1_11/a_230_79#
+ fine_freq_track_1/sky130_fd_sc_hs__nor3_1_9/a_198_368# fine_freq_track_1/sky130_fd_sc_hs__nand2_1_47/a_117_74#
+ fine_freq_track_1/sky130_fd_sc_hs__inv_4_47/Y fine_freq_track_1/sky130_fd_sc_hs__inv_4_9/A
+ fine_freq_track_1/sky130_fd_sc_hs__nand2_4_11/a_27_74# fine_freq_track_1/sky130_fd_sc_hs__a32oi_1_9/a_119_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_47/a_1934_94# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_43/a_1624_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_49/a_1598_93# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_47/a_33_74#
+ fine_freq_track_1/sky130_fd_sc_hs__sdlclkp_4_1/a_354_105# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_1/a_1547_508#
+ fine_freq_track_1/sky130_fd_sc_hs__nand2_1_91/a_117_74# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_81/a_812_138#
+ fine_freq_track_1/sky130_fd_sc_hs__a32oi_1_7/Y fine_freq_track_1/sky130_fd_sc_hs__a21oi_1_9/Y
+ fine_freq_track_1/sky130_fd_sc_hs__nand2_1_99/A fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_3/a_2010_409#
+ fine_freq_track_1/sky130_fd_sc_hs__a22oi_1_15/a_71_368# fine_freq_track_1/sky130_fd_sc_hs__xnor2_1_1/a_138_385#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_25/a_1647_81# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_27/a_714_127#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_85/a_1350_392# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_7/a_832_118#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_51/a_124_78# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_65/a_1647_81#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_25/a_1224_74# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_7/Q_N
+ fine_freq_track_1/sky130_fd_sc_hs__nor2_1_3/B fine_freq_track_1/sky130_fd_sc_hs__maj3_1_1/a_84_74#
+ fine_freq_track_1/sky130_fd_sc_hs__o21a_1_41/a_320_74# fine_freq_track_1/sky130_fd_sc_hs__inv_4_31/A
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_81/a_1678_395# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_85/D
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_51/a_789_463# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_13/a_1736_119#
+ fine_freq_track_1/sky130_fd_sc_hs__xor2_1_7/a_455_87# fine_freq_track_1/sky130_fd_sc_hs__a22o_1_13/a_222_392#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_13/a_1266_119# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_41/a_706_463#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_7/a_834_355# fine_freq_track_1/sky130_fd_sc_hs__o21a_1_19/A1
+ fine_freq_track_1/sky130_fd_sc_hs__o21a_1_5/A1 fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_33/a_319_360#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_17/a_494_366# fine_freq_track_1/sky130_fd_sc_hs__a21oi_1_41/a_29_368#
+ fine_freq_track_1/sky130_fd_sc_hs__inv_4_111/A fine_freq_track_1/sky130_fd_sc_hs__inv_4_9/Y
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_57/a_494_366# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_71/a_834_355#
+ fine_freq_track_1/sky130_fd_sc_hs__xnor2_1_9/a_293_74# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_37/a_922_127#
+ fine_freq_track_1/sky130_fd_sc_hs__nand2_2_1/A fine_freq_track_1/sky130_fd_sc_hs__a22o_1_29/a_52_123#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_33/a_1465_471# fine_freq_track_1/sky130_fd_sc_hs__o21a_1_25/a_376_387#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_25/a_890_138# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_21/a_832_118#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_63/a_2010_409# fine_freq_track_1/sky130_fd_sc_hs__dfxtp_4_2/a_651_503#
+ fine_freq_track_1/sky130_fd_sc_hs__nor2_1_7/A fine_freq_track_1/sky130_fd_sc_hs__inv_4_121/Y
+ fine_freq_track_1/sky130_fd_sc_hs__o31ai_1_3/B1 fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_65/a_890_138#
+ fine_freq_track_1/sky130_fd_sc_hs__nor2b_1_11/Y fine_freq_track_1/sky130_fd_sc_hs__nor2_1_73/B
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_31/D fine_freq_track_1/sky130_fd_sc_hs__o21a_1_77/X
+ fine_freq_track_1/sky130_fd_sc_hs__a21oi_1_27/a_117_74# fine_freq_track_1/sky130_fd_sc_hs__fa_2_19/a_1094_347#
+ fine_freq_track_1/sky130_fd_sc_hs__nor2_1_89/A fine_freq_track_1/sky130_fd_sc_hs__inv_4_61/Y
+ fine_freq_track_1/sky130_fd_sc_hs__nor2_1_75/Y fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_45/a_1550_119#
+ fine_freq_track_1/sky130_fd_sc_hs__nand4_2_1/D fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_35/a_300_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfxtp_2_9/a_538_429# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_13/a_2010_409#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_77/a_313_74# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_79/a_699_463#
+ fine_freq_track_1/sky130_fd_sc_hs__a21oi_1_71/a_117_74# fine_freq_track_1/sky130_fd_sc_hs__a21oi_1_9/a_117_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfxtp_2_11/a_708_101# fine_freq_track_1/sky130_fd_sc_hs__nor2_1_115/a_116_368#
+ fine_freq_track_1/sky130_fd_sc_hs__dfxtp_2_1/a_27_74# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_9/a_319_360#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_31/a_841_401# fine_freq_track_1/sky130_fd_sc_hs__nor2_1_77/Y
+ fine_freq_track_1/sky130_fd_sc_hs__fa_2_23/a_992_347# fine_freq_track_1/sky130_fd_sc_hs__a22o_1_5/a_230_79#
+ fine_freq_track_1/sky130_fd_sc_hs__nor2b_1_45/a_278_368# fine_freq_track_1/sky130_fd_sc_hs__inv_4_137/Y
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_11/a_313_74# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_7/a_812_138#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_43/a_125_78# fine_freq_track_1/sky130_fd_sc_hs__nor4_1_3/A
+ fine_freq_track_1/sky130_fd_sc_hs__o21a_1_7/a_320_74# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_71/a_812_138#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_75/a_37_78# fine_freq_track_1/sky130_fd_sc_hs__o21a_1_75/X
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_11/a_125_78# fine_freq_track_1/sky130_fd_sc_hs__and2_2_5/a_118_74#
+ fine_freq_track_1/sky130_fd_sc_hs__nor2b_1_19/a_27_112# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_15/a_1647_81#
+ fine_freq_track_1/sky130_fd_sc_hs__o21a_1_29/X fine_freq_track_1/sky130_fd_sc_hs__a22o_1_15/a_230_79#
+ fine_freq_track_1/sky130_fd_sc_hs__fa_2_3/a_1119_79# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_3/a_2026_424#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_11/a_1827_81# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_17/a_714_127#
+ fine_freq_track_1/sky130_fd_sc_hs__o22ai_1_1/A1 fine_freq_track_1/sky130_fd_sc_hs__and2_2_1/X
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_55/a_1647_81# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_15/a_1224_74#
+ fine_freq_track_1/sky130_fd_sc_hs__fa_2_17/B fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_39/a_507_368#
+ fine_freq_track_1/sky130_fd_sc_hs__dfxtp_2_5/D fine_freq_track_1/sky130_fd_sc_hs__nand2b_4_1/a_243_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_41/a_789_463# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_43/a_1627_493#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_35/a_498_360# fine_freq_track_1/sky130_fd_sc_hs__a22oi_1_21/a_159_74#
+ fine_freq_track_1/sky130_fd_sc_hs__nand2_1_95/a_117_74# fine_freq_track_1/sky130_fd_sc_hs__a32oi_1_5/Y
+ fine_freq_track_1/sky130_fd_sc_hs__fa_2_5/A fine_freq_track_1/sky130_fd_sc_hs__a22oi_1_19/a_71_368#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_21/a_834_355# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_33/a_1350_392#
+ fine_freq_track_1/sky130_fd_sc_hs__inv_4_71/Y fine_freq_track_1/sky130_fd_sc_hs__dfxtp_4_5/a_1178_124#
+ fine_freq_track_1/sky130_fd_sc_hs__a21oi_1_105/a_117_74# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_55/a_124_78#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_61/a_834_355# fine_freq_track_1/sky130_fd_sc_hs__sdlclkp_1_1/a_722_492#
+ fine_freq_track_1/sky130_fd_sc_hs__a222oi_1_3/a_369_392# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_5/a_1934_94#
+ fine_freq_track_1/sky130_fd_sc_hs__o211ai_1_5/a_116_368# fine_freq_track_1/sky130_fd_sc_hs__o21a_1_45/a_320_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_7/a_841_401# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_21/a_124_78#
+ fine_freq_track_1/sky130_fd_sc_hs__inv_4_101/A fine_freq_track_1/sky130_fd_sc_hs__a21oi_1_77/a_29_368#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_47/a_1678_395# fine_freq_track_1/sky130_fd_sc_hs__o21a_1_11/a_320_74#
+ fine_freq_track_1/sky130_fd_sc_hs__o21a_1_15/a_376_387# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_27/a_1482_48#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_15/a_890_138# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_11/a_832_118#
+ fine_freq_track_1/sky130_fd_sc_hs__a21oi_1_45/a_29_368# fine_freq_track_1/sky130_fd_sc_hs__inv_4_85/A
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_55/a_890_138# fine_freq_track_1/sky130_fd_sc_hs__a21oi_1_11/a_29_368#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_39/a_38_78# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_9/a_1550_119#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_31/a_33_74# fine_freq_track_1/sky130_fd_sc_hs__fa_2_1/a_336_347#
+ fine_freq_track_1/sky130_fd_sc_hs__dfxtp_4_3/a_696_458# fine_freq_track_1/sky130_fd_sc_hs__dfstp_2_1/a_1566_92#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_39/a_910_118# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_35/D
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_15/a_2026_424# fine_freq_track_1/sky130_fd_sc_hs__nor2b_1_1/a_278_368#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_69/a_699_463# fine_freq_track_1/sky130_fd_sc_hs__a22o_1_1/a_52_123#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_29/a_37_78# fine_freq_track_1/sky130_fd_sc_hs__nor2_1_105/a_116_368#
+ fine_freq_track_1/sky130_fd_sc_hs__dfxtp_4_2/D fine_freq_track_1/sky130_fd_sc_hs__fa_2_1/a_487_79#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_21/a_841_401# fine_freq_track_1/sky130_fd_sc_hs__o21a_1_51/X
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_23/a_1624_74# fine_freq_track_1/sky130_fd_sc_hs__fa_2_11/a_336_347#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_27/a_1934_94# fine_freq_track_1/sky130_fd_sc_hs__fa_2_13/a_992_347#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_15/Q_N fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_11/D
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_21/a_812_138# fine_freq_track_1/sky130_fd_sc_hs__a22o_1_11/a_52_123#
+ fine_freq_track_1/sky130_fd_sc_hs__dfstp_2_4/a_716_456# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_61/a_812_138#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_1/a_2010_409# fine_freq_track_1/sky130_fd_sc_hs__a21oi_1_75/a_117_74#
+ fine_freq_track_1/sky130_fd_sc_hs__o22ai_1_9/a_340_368# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_1/a_2026_424#
+ fine_freq_track_1/sky130_fd_sc_hs__dfstp_2_4/a_27_74# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_83/a_1350_392#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_47/a_313_74# fine_freq_track_1/sky130_fd_sc_hs__nand2_1_85/Y
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_45/a_1647_81# fine_freq_track_1/sky130_fd_sc_hs__a222o_1_1/a_27_390#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_23/a_120_74# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_29/a_507_368#
+ fine_freq_track_1/sky130_fd_sc_hs__nor2b_1_3/Y fine_freq_track_1/sky130_fd_sc_hs__a22o_1_9/a_230_79#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_31/a_789_463# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_47/a_125_78#
+ fine_freq_track_1/sky130_fd_sc_hs__xor2_1_3/a_355_368# fine_freq_track_1/sky130_fd_sc_hs__inv_4_109/Y
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_11/a_1736_119# fine_freq_track_1/sky130_fd_sc_hs__a21oi_1_123/a_29_368#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_11/a_1266_119# fine_freq_track_1/sky130_fd_sc_hs__dfxtp_2_7/a_644_504#
+ fine_freq_track_1/sky130_fd_sc_hs__or2_1_3/a_63_368# fine_freq_track_1/sky130_fd_sc_hs__a22o_1_19/a_230_79#
+ fine_freq_track_1/sky130_fd_sc_hs__fa_2_15/a_683_347# fine_freq_track_1/sky130_fd_sc_hs__a31oi_1_1/a_145_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_51/a_834_355# fine_freq_track_1/sky130_fd_sc_hs__maj3_1_3/X
+ fine_freq_track_1/sky130_fd_sc_hs__o21a_1_33/a_83_244# fine_freq_track_1/sky130_fd_sc_hs__dfstp_2_7/D
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_31/a_1434_74# fine_freq_track_1/sky130_fd_sc_hs__o21a_1_3/X
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_31/a_1465_471# fine_freq_track_1/sky130_fd_sc_hs__a22oi_1_25/a_159_74#
+ fine_freq_track_1/sky130_fd_sc_hs__nand2b_1_3/Y fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_17/a_1482_48#
+ fine_freq_track_1/sky130_fd_sc_hs__nand3b_2_1/a_403_54# fine_freq_track_1/sky130_fd_sc_hs__o22ai_1_3/Y
+ fine_freq_track_1/sky130_fd_sc_hs__a21oi_1_109/a_117_74# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_45/a_890_138#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_59/a_124_78# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_7/a_1550_119#
+ fine_freq_track_1/sky130_fd_sc_hs__nand2_1_33/a_117_74# fine_freq_track_1/sky130_fd_sc_hs__o21a_1_49/a_320_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_13/a_817_508# fine_freq_track_1/sky130_fd_sc_hs__fa_2_17/a_1094_347#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_25/a_124_78# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_43/a_1550_119#
+ fine_freq_track_1/sky130_fd_sc_hs__nor3_1_3/a_114_368# fine_freq_track_1/sky130_fd_sc_hs__xnor2_1_11/a_293_74#
+ fine_freq_track_1/sky130_fd_sc_hs__o22ai_1_9/A1 fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_11/a_2010_409#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_59/a_699_463# fine_freq_track_1/sky130_fd_sc_hs__nor2_1_99/a_116_368#
+ fine_freq_track_1/sky130_fd_sc_hs__nor2_1_59/A fine_freq_track_1/sky130_fd_sc_hs__a21oi_1_121/a_117_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_11/a_841_401# fine_freq_track_1/sky130_fd_sc_hs__a22o_1_11/a_132_392#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_17/a_1934_94# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_13/a_1624_74#
+ fine_freq_track_1/sky130_fd_sc_hs__clkbuf_2_1/a_43_192# fine_freq_track_1/sky130_fd_sc_hs__nor2b_1_25/a_278_368#
+ fine_freq_track_1/sky130_fd_sc_hs__o21a_1_15/X fine_freq_track_1/sky130_fd_sc_hs__a21oi_1_93/a_29_368#
+ fine_freq_track_1/sky130_fd_sc_hs__nand2_4_7/a_27_74# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_51/a_812_138#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_39/a_856_304# fine_freq_track_1/sky130_fd_sc_hs__nor3_1_1/C
+ fine_freq_track_1/sky130_fd_sc_hs__nor2_1_9/B fine_freq_track_1/sky130_fd_sc_hs__maj3_1_3/a_226_384#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_7/a_1434_74# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_39/a_850_127#
+ fine_freq_track_1/sky130_fd_sc_hs__a22o_1_5/a_52_123# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_69/a_37_78#
+ fine_freq_track_1/sky130_fd_sc_hs__fa_2_5/a_487_79# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_35/a_1647_81#
+ fine_freq_track_1/sky130_fd_sc_hs__nor2_1_83/Y fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_19/a_507_368#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_5/a_1827_81# fine_freq_track_1/sky130_fd_sc_hs__nand4_1_1/Y
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_37/a_714_127# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_73/a_1647_81#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_35/a_1224_74# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_41/a_1627_493#
+ fine_freq_track_1/sky130_fd_sc_hs__a22o_1_15/a_52_123# fine_freq_track_1/sky130_fd_sc_hs__o22ai_1_9/a_142_368#
+ fine_freq_track_1/sky130_fd_sc_hs__dfstp_2_5/a_1278_74# fine_freq_track_1/sky130_fd_sc_hs__a22o_1_23/a_222_392#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_29/a_1736_119# fine_freq_track_1/sky130_fd_sc_hs__inv_4_95/Y
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_31/a_1350_392# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_23/a_38_78#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_41/a_319_360# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_27/a_494_366#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_41/a_834_355# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_29/a_1266_119#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_49/a_1350_392# fine_freq_track_1/sky130_fd_sc_hs__a21oi_1_82/Y
+ fine_freq_track_1/sky130_fd_sc_hs__nor3_1_13/a_198_368# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_19/a_313_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_21/a_1434_74# fine_freq_track_1/sky130_fd_sc_hs__a21oi_1_13/a_117_74#
+ fine_freq_track_1/sky130_fd_sc_hs__o2bb2ai_1_1/a_131_383# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_19/a_125_78#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_13/a_37_78# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_61/a_2010_409#
+ fine_freq_track_1/sky130_fd_sc_hs__nand4_1_1/a_259_74# fine_freq_track_1/sky130_fd_sc_hs__dfxtp_2_5/a_206_368#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_35/a_890_138# fine_freq_track_1/sky130_fd_sc_hs__a31oi_1_1/A2
+ fine_freq_track_1/sky130_fd_sc_hs__o21a_1_73/a_376_387# fine_freq_track_1/sky130_fd_sc_hs__nor4_1_3/D
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_73/a_890_138# fine_freq_track_1/sky130_fd_sc_hs__nor3_1_9/A
+ fine_freq_track_1/sky130_fd_sc_hs__nor2b_1_1/Y fine_freq_track_1/sky130_fd_sc_hs__dfsbp_2_1/Q
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_43/a_817_508# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_41/a_1550_119#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_13/a_2026_424# fine_freq_track_1/sky130_fd_sc_hs__nor2_1_41/B
+ fine_freq_track_1/sky130_fd_sc_hs__o21a_1_45/X fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_5/a_796_463#
+ fine_freq_track_1/sky130_fd_sc_hs__nor2_1_89/a_116_368# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_29/a_2010_409#
+ fine_freq_track_1/sky130_fd_sc_hs__nor2b_1_15/a_278_368# fine_freq_track_1/sky130_fd_sc_hs__nand2_1_37/a_117_74#
+ fine_freq_track_1/sky130_fd_sc_hs__a22oi_1_23/a_339_74# fine_freq_track_1/sky130_fd_sc_hs__dfsbp_2_1/a_1501_92#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_47/a_1598_93# fine_freq_track_1/sky130_fd_sc_hs__dfsbp_2_1/a_1521_508#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_91/a_1627_493# fine_freq_track_1/sky130_fd_sc_hs__a22oi_1_5/a_159_74#
+ fine_freq_track_1/sky130_fd_sc_hs__xnor2_1_15/a_293_74# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_41/a_812_138#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_29/a_856_304# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_29/a_850_127#
+ fine_freq_track_1/sky130_fd_sc_hs__dfxtp_2_1/a_431_508# fine_freq_track_1/sky130_fd_sc_hs__nand2_1_81/a_117_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_73/a_124_78# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_81/a_1350_392#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_83/D fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_41/a_124_78#
+ fine_freq_track_1/sky130_fd_sc_hs__o21a_1_13/A1 fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_63/a_1647_81#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_11/a_789_463# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_49/a_507_368#
+ fine_freq_track_1/sky130_fd_sc_hs__a21oi_1_97/a_29_368# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_29/a_796_463#
+ fine_freq_track_1/sky130_fd_sc_hs__o21a_1_31/a_320_74# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_43/a_498_360#
+ fine_freq_track_1/sky130_fd_sc_hs__dfstp_2_5/a_398_74# fine_freq_track_1/sky130_fd_sc_hs__a2bb2oi_1_1/Y
+ fine_freq_track_1/sky130_fd_sc_hs__fa_2_15/a_27_378# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_59/a_1627_493#
+ fine_freq_track_1/sky130_fd_sc_hs__a22o_1_9/a_52_123# fine_freq_track_1/sky130_fd_sc_hs__dfxtp_4_3/a_1178_124#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_37/a_37_78# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_31/a_834_355#
+ fine_freq_track_1/sky130_fd_sc_hs__fa_2_9/a_487_79# fine_freq_track_1/sky130_fd_sc_hs__a21oi_1_31/a_29_368#
+ fine_freq_track_1/sky130_fd_sc_hs__fa_2_23/a_1119_79# fine_freq_track_1/sky130_fd_sc_hs__o211ai_1_5/Y
+ fine_freq_track_1/sky130_fd_sc_hs__nand2_1_23/Y fine_freq_track_1/sky130_fd_sc_hs__nand2_4_15/a_27_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_19/a_1547_508# fine_freq_track_1/sky130_fd_sc_hs__nor2_1_13/Y
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_11/a_1434_74# fine_freq_track_1/sky130_fd_sc_hs__a22o_1_19/a_52_123#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_45/a_1678_395# fine_freq_track_1/sky130_fd_sc_hs__o21ai_1_9/Y
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_37/a_1482_48# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_47/a_1465_471#
+ fine_freq_track_1/sky130_fd_sc_hs__o21a_1_63/a_376_387# fine_freq_track_1/sky130_fd_sc_hs__nor2_2_1/A
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_79/a_2010_409# fine_freq_track_1/sky130_fd_sc_hs__a21oi_1_49/a_117_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_63/a_890_138# fine_freq_track_1/sky130_fd_sc_hs__dfxtp_4_3/a_544_485#
+ fine_freq_track_1/sky130_fd_sc_hs__fa_2_15/a_701_79# fine_freq_track_1/sky130_fd_sc_hs__a21oi_1_17/a_117_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_3/a_313_74# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_33/a_817_508#
+ fine_freq_track_1/sky130_fd_sc_hs__nor2_1_79/a_116_368# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_39/a_699_463#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_25/a_300_74# fine_freq_track_1/sky130_fd_sc_hs__dfxtp_2_7/a_538_429#
+ fine_freq_track_1/sky130_fd_sc_hs__nand4_1_5/a_259_74# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_41/a_120_74#
+ fine_freq_track_1/sky130_fd_sc_hs__fa_2_7/a_484_347# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_5/D
+ fine_freq_track_1/sky130_fd_sc_hs__a21oi_1_61/a_117_74# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_5/a_120_74#
+ fine_freq_track_1/sky130_fd_sc_hs__xnor2_1_9/a_376_368# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_37/a_1934_94#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_33/a_1624_74# fine_freq_track_1/sky130_fd_sc_hs__inv_2_1/Y
+ fine_freq_track_1/sky130_fd_sc_hs__fa_2_21/a_336_347# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_3/a_922_127#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_19/a_856_304# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_31/a_812_138#
+ fine_freq_track_1/sky130_fd_sc_hs__a32oi_1_5/A1 fine_freq_track_1/sky130_fd_sc_hs__o21a_1_37/X
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_19/a_850_127# fine_freq_track_1/sky130_fd_sc_hs__nand2_1_121/a_117_74#
+ fine_freq_track_1/sky130_fd_sc_hs__fa_2_17/a_484_347# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_3/a_1482_48#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_53/a_1647_81# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_19/a_796_463#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_45/Q_N fine_freq_track_1/sky130_fd_sc_hs__o22ai_1_1/a_27_74#
+ fine_freq_track_1/sky130_fd_sc_hs__a22oi_1_11/a_159_74# fine_freq_track_1/sky130_fd_sc_hs__dfxtp_2_9/a_1125_508#
+ fine_freq_track_1/sky130_fd_sc_hs__xor2_1_5/a_158_392# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_27/a_1736_119#
+ fine_freq_track_1/sky130_fd_sc_hs__nand2_1_85/a_117_74# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_37/Q_N
+ fine_freq_track_1/sky130_fd_sc_hs__nand3b_2_1/a_206_74# fine_freq_track_1/sky130_fd_sc_hs__dfxtp_4_2/a_1178_124#
+ fine_freq_track_1/sky130_fd_sc_hs__conb_1_1/a_21_290# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_9/a_33_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_31/a_706_463# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_27/a_1266_119#
+ fine_freq_track_1/sky130_fd_sc_hs__fa_2_13/a_1119_79# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_27/Q_N
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_47/a_1350_392# fine_freq_track_1/sky130_fd_sc_hs__sdlclkp_4_1/a_119_143#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_17/a_38_78# fine_freq_track_1/sky130_fd_sc_hs__nor2_1_11/Y
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_45/a_124_78# fine_freq_track_1/sky130_fd_sc_hs__dfxtp_2_5/a_27_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_5/a_1598_93# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_19/Q_N
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_85/a_494_366# fine_freq_track_1/sky130_fd_sc_hs__o31ai_1_5/Y
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_9/a_1624_74# fine_freq_track_1/sky130_fd_sc_hs__dfstp_2_7/a_398_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfxtp_4_9/a_206_368# fine_freq_track_1/sky130_fd_sc_hs__o21a_1_13/a_376_387#
+ fine_freq_track_1/sky130_fd_sc_hs__sdlclkp_4_1/a_1289_368# fine_freq_track_1/sky130_fd_sc_hs__nand2_2_3/Y
+ fine_freq_track_1/sky130_fd_sc_hs__o21a_1_53/a_376_387# fine_freq_track_1/sky130_fd_sc_hs__o211ai_1_7/a_31_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_5/a_1550_119# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_53/a_890_138#
+ fine_freq_track_1/sky130_fd_sc_hs__fa_2_15/a_1094_347# fine_freq_track_1/sky130_fd_sc_hs__fa_2_23/a_27_79#
+ fine_freq_track_1/sky130_fd_sc_hs__fa_2_1/a_992_347# fine_freq_track_1/sky130_fd_sc_hs__dfxtp_4_2/a_696_458#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_23/a_817_508# fine_freq_track_1/sky130_fd_sc_hs__o21a_1_9/a_376_387#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_19/a_33_74# fine_freq_track_1/sky130_fd_sc_hs__o31ai_1_5/a_114_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_29/a_699_463# fine_freq_track_1/sky130_fd_sc_hs__nor2_1_69/a_116_368#
+ fine_freq_track_1/sky130_fd_sc_hs__inv_4_73/Y fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_27/a_2010_409#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_33/a_38_78# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_67/a_699_463#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_15/D fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_7/a_706_463#
+ fine_freq_track_1/sky130_fd_sc_hs__fa_2_11/a_992_347# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_27/a_1598_93#
+ fine_freq_track_1/sky130_fd_sc_hs__o21ai_1_1/B1 fine_freq_track_1/sky130_fd_sc_hs__dfxtp_2_5/a_708_101#
+ fine_freq_track_1/sky130_fd_sc_hs__fa_2_9/a_27_79# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_21/a_37_78#
+ fine_freq_track_1/sky130_fd_sc_hs__dfstp_2_1/a_716_456# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_49/a_856_304#
+ fine_freq_track_1/sky130_fd_sc_hs__dfxtp_4_2/a_27_74# fine_freq_track_1/sky130_fd_sc_hs__dfxtp_4_7/Q
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_49/a_850_127# fine_freq_track_1/sky130_fd_sc_hs__a21oi_1_65/a_117_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_9/a_120_74# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_37/a_313_74#
+ fine_freq_track_1/sky130_fd_sc_hs__fa_2_3/a_683_347# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_49/a_1827_81#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_35/a_33_74# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_83/a_1647_81#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_43/a_1224_74# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_89/a_1827_81#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_5/a_789_463# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_23/a_498_360#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_47/a_796_463# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_57/a_1627_493#
+ fine_freq_track_1/sky130_fd_sc_hs__a21oi_1_113/a_29_368# fine_freq_track_1/sky130_fd_sc_hs__dfxtp_2_7/a_1125_508#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_3/a_300_74# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_5/a_910_118#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_21/a_706_463# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_11/a_834_355#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_17/a_1547_508# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_1/a_494_366#
+ fine_freq_track_1/sky130_fd_sc_hs__nand2_2_15/a_27_74# fine_freq_track_1/sky130_fd_sc_hs__o21ai_1_3/a_162_368#
+ fine_freq_track_1/sky130_fd_sc_hs__o21a_1_23/a_83_244# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_75/a_494_366#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_43/a_1678_395# fine_freq_track_1/sky130_fd_sc_hs__fa_2_9/A
+ fine_freq_track_1/sky130_fd_sc_hs__a222oi_1_3/a_697_74# fine_freq_track_1/sky130_fd_sc_hs__a22oi_1_15/a_159_74#
+ fine_freq_track_1/sky130_fd_sc_hs__a22o_1_7/a_132_392# fine_freq_track_1/sky130_fd_sc_hs__nand2_1_89/a_117_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_45/a_1465_471# fine_freq_track_1/sky130_fd_sc_hs__dfxtp_4_9/a_437_503#
+ fine_freq_track_1/sky130_fd_sc_hs__o21a_1_43/a_376_387# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_77/a_2010_409#
+ fine_freq_track_1/sky130_fd_sc_hs__xnor2_1_1/Y fine_freq_track_1/sky130_fd_sc_hs__nor2_1_95/B
+ fine_freq_track_1/sky130_fd_sc_hs__nand2b_1_3/a_269_74# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_83/a_890_138#
+ fine_freq_track_1/sky130_fd_sc_hs__nand2_1_23/a_117_74# fine_freq_track_1/sky130_fd_sc_hs__o21a_1_39/a_320_74#
+ fine_freq_track_1/sky130_fd_sc_hs__fa_2_7/B fine_freq_track_1/sky130_fd_sc_hs__nor2_1_47/Y
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_11/a_2026_424# fine_freq_track_1/sky130_fd_sc_hs__dfsbp_2_1/a_1531_118#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_29/a_910_118# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_15/a_124_78#
+ fine_freq_track_1/sky130_fd_sc_hs__nor3_1_3/B fine_freq_track_1/sky130_fd_sc_hs__dfxtp_4_7/a_735_102#
+ fine_freq_track_1/sky130_fd_sc_hs__nor2_1_91/B fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_19/a_699_463#
+ fine_freq_track_1/sky130_fd_sc_hs__nor2_1_59/a_116_368# fine_freq_track_1/sky130_fd_sc_hs__fa_2_9/a_1094_347#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_25/a_2010_409# fine_freq_track_1/sky130_fd_sc_hs__a21oi_1_39/a_29_368#
+ fine_freq_track_1/sky130_fd_sc_hs__a21oi_1_111/a_117_74# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_25/D
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_17/a_1598_93# fine_freq_track_1/sky130_fd_sc_hs__fa_2_1/B
+ fine_freq_track_1/sky130_fd_sc_hs__dfxtp_4_9/a_1034_424# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_11/a_812_138#
+ fine_freq_track_1/sky130_fd_sc_hs__a22oi_1_13/Y fine_freq_track_1/sky130_fd_sc_hs__inv_4_83/A
+ fine_freq_track_1/sky130_fd_sc_hs__nand4_1_3/a_181_74# fine_freq_track_1/sky130_fd_sc_hs__maj3_1_1/a_226_384#
+ fine_freq_track_1/sky130_fd_sc_hs__a22oi_1_1/a_71_368# fine_freq_track_1/sky130_fd_sc_hs__fa_2_7/a_1205_79#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_9/a_1647_81# fine_freq_track_1/sky130_fd_sc_hs__nand2_4_1/a_27_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_79/a_1827_81# fine_freq_track_1/sky130_fd_sc_hs__o21a_1_13/X
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_13/a_498_360# fine_freq_track_1/sky130_fd_sc_hs__sdlclkp_1_1/a_1238_94#
+ fine_freq_track_1/sky130_fd_sc_hs__nor2_1_9/a_116_368# fine_freq_track_1/sky130_fd_sc_hs__dfstp_2_4/a_1278_74#
+ fine_freq_track_1/sky130_fd_sc_hs__inv_4_5/A fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_11/a_706_463#
+ fine_freq_track_1/sky130_fd_sc_hs__a22o_1_21/a_222_392# fine_freq_track_1/sky130_fd_sc_hs__a21oi_1_69/a_117_74#
+ fine_freq_track_1/sky130_fd_sc_hs__nor2_1_43/Y fine_freq_track_1/sky130_fd_sc_hs__fa_2_17/a_1205_79#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_25/a_494_366# fine_freq_track_1/sky130_fd_sc_hs__a211oi_4_1/a_901_368#
+ fine_freq_track_1/sky130_fd_sc_hs__a21oi_1_35/a_117_74# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_65/a_494_366#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_45/a_922_127# fine_freq_track_1/sky130_fd_sc_hs__nand4_2_1/a_515_74#
+ fine_freq_track_1/sky130_fd_sc_hs__nor3_1_7/A fine_freq_track_1/sky130_fd_sc_hs__o21a_1_33/a_376_387#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_45/a_1482_48# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_39/a_832_118#
+ fine_freq_track_1/sky130_fd_sc_hs__fa_2_21/B fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_3/a_1550_119#
+ fine_freq_track_1/sky130_fd_sc_hs__dfxtp_2_3/a_206_368# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_9/a_890_138#
+ fine_freq_track_1/sky130_fd_sc_hs__fa_2_13/a_1094_347# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_3/a_714_127#
+ fine_freq_track_1/sky130_fd_sc_hs__o21a_1_43/X fine_freq_track_1/sky130_fd_sc_hs__fa_2_17/a_487_79#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_19/a_910_118# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_41/a_817_508#
+ fine_freq_track_1/sky130_fd_sc_hs__a22oi_1_19/a_159_74# fine_freq_track_1/sky130_fd_sc_hs__nor2_1_49/a_116_368#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_29/a_2026_424# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_47/a_699_463#
+ fine_freq_track_1/sky130_fd_sc_hs__o21a_1_71/a_83_244# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_5/D
+ fine_freq_track_1/sky130_fd_sc_hs__nand2b_1_7/a_269_74# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_87/a_699_463#
+ fine_freq_track_1/sky130_fd_sc_hs__nor2_1_123/a_116_368# fine_freq_track_1/sky130_fd_sc_hs__a222oi_1_3/a_119_74#
+ fine_freq_track_1/sky130_fd_sc_hs__nor2b_1_13/a_278_368# fine_freq_track_1/sky130_fd_sc_hs__nand2_1_27/a_117_74#
+ fine_freq_track_1/sky130_fd_sc_hs__a22oi_1_13/a_339_74# fine_freq_track_1/sky130_fd_sc_hs__nor3_1_7/a_198_368#
+ fine_freq_track_1/sky130_fd_sc_hs__a22o_1_9/a_222_392# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_41/a_1624_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfstp_2_7/a_1521_508# fine_freq_track_1/sky130_fd_sc_hs__o31ai_1_7/a_119_368#
+ fine_freq_track_1/sky130_fd_sc_hs__inv_4_19/Y fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_87/a_37_78#
+ fine_freq_track_1/sky130_fd_sc_hs__nand2_1_71/a_117_74# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_15/a_37_78#
+ fine_freq_track_1/sky130_fd_sc_hs__a21oi_1_115/a_117_74# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_63/a_124_78#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_31/a_124_78# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_23/a_1224_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_69/a_1827_81# fine_freq_track_1/sky130_fd_sc_hs__o211ai_1_1/a_311_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_47/a_507_368# fine_freq_track_1/sky130_fd_sc_hs__a21oi_1_87/a_29_368#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_27/a_796_463# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_55/a_1627_493#
+ fine_freq_track_1/sky130_fd_sc_hs__o21a_1_21/a_320_74# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_25/a_1736_119#
+ fine_freq_track_1/sky130_fd_sc_hs__o21ai_1_5/a_27_74# fine_freq_track_1/sky130_fd_sc_hs__dfstp_2_7/a_767_384#
+ fine_freq_track_1/sky130_fd_sc_hs__a21oi_1_53/a_29_368# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_25/a_1266_119#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_41/a_38_78# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_45/a_1350_392#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_31/a_319_360# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_15/a_494_366#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_5/a_834_355# fine_freq_track_1/sky130_fd_sc_hs__a21oi_1_21/a_29_368#
+ fine_freq_track_1/sky130_fd_sc_hs__inv_4_93/A fine_freq_track_1/sky130_fd_sc_hs__o21ai_1_7/Y
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_55/a_494_366# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_41/a_1678_395#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_35/a_922_127# fine_freq_track_1/sky130_fd_sc_hs__o21a_1_73/X
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_31/a_37_78# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_43/a_1465_471#
+ fine_freq_track_1/sky130_fd_sc_hs__a21oi_1_3/a_29_368# fine_freq_track_1/sky130_fd_sc_hs__o21a_1_23/a_376_387#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_75/a_2010_409# fine_freq_track_1/sky130_fd_sc_hs__fa_2_19/a_1202_368#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_1/a_1550_119# fine_freq_track_1/sky130_fd_sc_hs__fa_2_11/a_1094_347#
+ fine_freq_track_1/sky130_fd_sc_hs__dfxtp_4_2/a_544_485# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_47/a_300_74#
+ fine_freq_track_1/sky130_fd_sc_hs__nor2_2_3/a_35_368# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_31/a_817_508#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_47/a_910_118# fine_freq_track_1/sky130_fd_sc_hs__nor2_1_39/a_116_368#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_27/a_2026_424# fine_freq_track_1/sky130_fd_sc_hs__o21a_1_5/B1
+ fine_freq_track_1/sky130_fd_sc_hs__fa_2_7/a_1094_347# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_39/Q_N
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_37/a_699_463# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_15/a_300_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_3/a_699_463# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_57/a_313_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_77/a_699_463# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_31/a_120_74#
+ fine_freq_track_1/sky130_fd_sc_hs__nor2_1_113/a_116_368# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_39/a_841_401#
+ fine_freq_track_1/sky130_fd_sc_hs__a222o_1_1/a_386_74# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_7/a_319_360#
+ fine_freq_track_1/sky130_fd_sc_hs__dfxtp_4_7/a_1034_424# fine_freq_track_1/sky130_fd_sc_hs__fa_2_21/a_992_347#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_1/a_922_127# fine_freq_track_1/sky130_fd_sc_hs__nor2b_1_43/a_278_368#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_37/a_1598_93# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_23/a_125_78#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_5/a_812_138# fine_freq_track_1/sky130_fd_sc_hs__nor2b_1_5/a_27_112#
+ fine_freq_track_1/sky130_fd_sc_hs__o21a_1_75/a_83_244# fine_freq_track_1/sky130_fd_sc_hs__inv_4_115/Y
+ fine_freq_track_1/sky130_fd_sc_hs__a211oi_1_3/a_71_368# fine_freq_track_1/sky130_fd_sc_hs__nand2_1_51/Y
+ fine_freq_track_1/sky130_fd_sc_hs__o21a_1_69/A2 fine_freq_track_1/sky130_fd_sc_hs__fa_2_1/a_1119_79#
+ fine_freq_track_1/sky130_fd_sc_hs__dfstp_2_5/D fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_1/a_1482_48#
+ fine_freq_track_1/sky130_fd_sc_hs__a22oi_1_17/a_339_74# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_13/a_1224_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_59/a_1827_81# fine_freq_track_1/sky130_fd_sc_hs__dfxtp_2_11/a_644_504#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_17/a_796_463# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_91/a_1678_395#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_53/a_1627_493# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_49/a_789_463#
+ fine_freq_track_1/sky130_fd_sc_hs__dfxtp_2_5/a_1125_508# fine_freq_track_1/sky130_fd_sc_hs__nor2b_1_43/a_27_112#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_33/a_498_360# fine_freq_track_1/sky130_fd_sc_hs__nand2b_4_1/a_31_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_89/a_789_463# fine_freq_track_1/sky130_fd_sc_hs__dfsbp_2_1/a_757_401#
+ fine_freq_track_1/sky130_fd_sc_hs__nand2_1_75/a_117_74# fine_freq_track_1/sky130_fd_sc_hs__a21oi_1_119/a_117_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_67/a_124_78# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_21/a_319_360#
+ fine_freq_track_1/sky130_fd_sc_hs__fa_2_11/a_1119_79# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_15/a_1547_508#
+ fine_freq_track_1/sky130_fd_sc_hs__dfstp_2_5/a_225_74# fine_freq_track_1/sky130_fd_sc_hs__nand2_1_41/a_117_74#
+ fine_freq_track_1/sky130_fd_sc_hs__fa_2_23/a_683_347# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_45/a_494_366#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_35/a_124_78# fine_freq_track_1/sky130_fd_sc_hs__a222oi_1_1/a_369_392#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_3/a_1934_94# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_25/a_922_127#
+ fine_freq_track_1/sky130_fd_sc_hs__o21a_1_25/a_320_74# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_1/a_33_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_59/a_1678_395# fine_freq_track_1/sky130_fd_sc_hs__a22oi_1_9/a_71_368#
+ fine_freq_track_1/sky130_fd_sc_hs__o21a_1_67/X fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_7/a_37_78#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_11/a_38_78# fine_freq_track_1/sky130_fd_sc_hs__xnor2_1_9/a_112_119#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_25/a_1482_48# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_73/a_2010_409#
+ fine_freq_track_1/sky130_fd_sc_hs__inv_4_7/A fine_freq_track_1/sky130_fd_sc_hs__nand2_1_3/a_117_74#
+ fine_freq_track_1/sky130_fd_sc_hs__a21oi_1_25/a_29_368# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_5/a_507_368#
+ fine_freq_track_1/sky130_fd_sc_hs__xnor2_1_9/A fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_21/a_817_508#
+ fine_freq_track_1/sky130_fd_sc_hs__nor2_1_29/a_116_368# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_71/a_37_78#
+ fine_freq_track_1/sky130_fd_sc_hs__xor2_1_3/a_455_87# fine_freq_track_1/sky130_fd_sc_hs__a21oi_1_7/a_29_368#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_17/D fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_23/a_2010_409#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_9/a_498_360# fine_freq_track_1/sky130_fd_sc_hs__nand2_2_9/B
+ fine_freq_track_1/sky130_fd_sc_hs__nor2_1_103/a_116_368# fine_freq_track_1/sky130_fd_sc_hs__dfxtp_2_7/a_27_74#
+ fine_freq_track_1/sky130_fd_sc_hs__nor2b_1_33/a_278_368# fine_freq_track_1/sky130_fd_sc_hs__sdlclkp_1_1/a_709_54#
+ fine_freq_track_1/sky130_fd_sc_hs__inv_4_95/A fine_freq_track_1/sky130_fd_sc_hs__nand2_2_11/Y
+ fine_freq_track_1/sky130_fd_sc_hs__dfxtp_2_3/a_708_101# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_47/a_856_304#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_47/a_850_127# fine_freq_track_1/sky130_fd_sc_hs__a21oi_1_55/a_117_74#
+ fine_freq_track_1/sky130_fd_sc_hs__inv_4_29/Y fine_freq_track_1/sky130_fd_sc_hs__o22ai_1_7/a_340_368#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_43/a_1647_81# fine_freq_track_1/sky130_fd_sc_hs__a21oi_1_15/Y
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_27/a_507_368# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_45/a_714_127#
+ fine_freq_track_1/sky130_fd_sc_hs__dfxtp_2_3/a_1125_508# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_23/a_1736_119#
+ fine_freq_track_1/sky130_fd_sc_hs__a31oi_1_1/a_136_368# fine_freq_track_1/sky130_fd_sc_hs__o21a_1_77/A2
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_27/a_125_78# fine_freq_track_1/sky130_fd_sc_hs__xor2_1_1/a_355_368#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_79/a_789_463# fine_freq_track_1/sky130_fd_sc_hs__nor2b_1_9/a_27_112#
+ fine_freq_track_1/sky130_fd_sc_hs__a21oi_1_103/a_29_368# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_1/a_125_78#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_23/a_1266_119# fine_freq_track_1/sky130_fd_sc_hs__nand2_1_115/a_117_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_43/a_1350_392# fine_freq_track_1/sky130_fd_sc_hs__nor2_1_29/B
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_11/a_319_360# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_13/a_1547_508#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_9/a_38_78# fine_freq_track_1/sky130_fd_sc_hs__nand2_2_3/B
+ fine_freq_track_1/sky130_fd_sc_hs__nor2_1_19/B fine_freq_track_1/sky130_fd_sc_hs__fa_2_13/a_683_347#
+ fine_freq_track_1/sky130_fd_sc_hs__xor2_1_11/a_158_392# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_35/a_494_366#
+ fine_freq_track_1/sky130_fd_sc_hs__fa_2_1/a_27_378# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_15/a_922_127#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_73/a_494_366# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_7/a_124_78#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_39/a_1434_74# fine_freq_track_1/sky130_fd_sc_hs__nor2b_1_47/a_27_112#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_41/a_1465_471# fine_freq_track_1/sky130_fd_sc_hs__nor3_1_13/Y
+ fine_freq_track_1/sky130_fd_sc_hs__nand2_1_79/a_117_74# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_15/a_1482_48#
+ fine_freq_track_1/sky130_fd_sc_hs__fa_2_17/a_1202_368# fine_freq_track_1/sky130_fd_sc_hs__nor2b_1_13/a_27_112#
+ fine_freq_track_1/sky130_fd_sc_hs__o31ai_1_7/A1 fine_freq_track_1/sky130_fd_sc_hs__dfstp_2_7/a_225_74#
+ fine_freq_track_1/sky130_fd_sc_hs__nand2_1_45/a_117_74# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_43/a_890_138#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_39/a_124_78# fine_freq_track_1/sky130_fd_sc_hs__o211ai_1_9/a_311_74#
+ fine_freq_track_1/sky130_fd_sc_hs__nand2_1_13/a_117_74# fine_freq_track_1/sky130_fd_sc_hs__o21a_1_29/a_320_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_11/a_817_508# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_27/a_910_118#
+ fine_freq_track_1/sky130_fd_sc_hs__nor2_1_19/a_116_368# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_25/a_2026_424#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_9/a_1627_493# fine_freq_track_1/sky130_fd_sc_hs__a22oi_1_11/Y
+ fine_freq_track_1/sky130_fd_sc_hs__fa_2_5/a_1094_347# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_21/a_2010_409#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_17/a_699_463# fine_freq_track_1/sky130_fd_sc_hs__nor3_1_1/a_114_368#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_83/a_124_78# fine_freq_track_1/sky130_fd_sc_hs__fa_2_1/a_701_79#
+ fine_freq_track_1/sky130_fd_sc_hs__nand2_1_7/a_117_74# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_57/a_699_463#
+ fine_freq_track_1/sky130_fd_sc_hs__nor2_1_97/a_116_368# fine_freq_track_1/sky130_fd_sc_hs__o21a_1_73/a_320_74#
+ fine_freq_track_1/sky130_fd_sc_hs__a21oi_1_29/a_29_368# fine_freq_track_1/sky130_fd_sc_hs__a21oi_1_101/a_117_74#
+ fine_freq_track_1/sky130_fd_sc_hs__or2_1_1/B fine_freq_track_1/sky130_fd_sc_hs__o31ai_1_7/a_203_368#
+ fine_freq_track_1/sky130_fd_sc_hs__dfxtp_4_5/a_1034_424# fine_freq_track_1/sky130_fd_sc_hs__nor2b_1_23/a_278_368#
+ fine_freq_track_1/sky130_fd_sc_hs__a31oi_1_1/a_223_74# fine_freq_track_1/sky130_fd_sc_hs__a21oi_1_73/a_29_368#
+ fine_freq_track_1/sky130_fd_sc_hs__nor3_1_15/Y fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_33/a_1647_81#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_39/a_1827_81# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_17/a_507_368#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_35/a_714_127# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_33/a_1224_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_21/a_1736_119# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_37/a_796_463#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_69/a_789_463# fine_freq_track_1/sky130_fd_sc_hs__dfstp_2_7/a_2022_94#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_21/a_1266_119# fine_freq_track_1/sky130_fd_sc_hs__o22ai_1_7/a_142_368#
+ fine_freq_track_1/sky130_fd_sc_hs__nor2_1_7/a_116_368# fine_freq_track_1/sky130_fd_sc_hs__dfstp_2_1/a_1278_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_39/a_120_74# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_49/a_37_78#
+ fine_freq_track_1/sky130_fd_sc_hs__a21oi_1_59/a_117_74# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_49/a_834_355#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_89/a_834_355# fine_freq_track_1/sky130_fd_sc_hs__xor2_1_5/a_194_125#
+ fine_freq_track_1/sky130_fd_sc_hs__nor3_1_11/a_198_368# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_63/a_494_366#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_57/a_1678_395# fine_freq_track_1/sky130_fd_sc_hs__a21oi_1_107/a_29_368#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_5/a_856_304# fine_freq_track_1/sky130_fd_sc_hs__nand2_1_119/a_117_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_5/a_850_127# fine_freq_track_1/sky130_fd_sc_hs__o21a_1_41/X
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_43/a_313_74# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_33/a_890_138#
+ fine_freq_track_1/sky130_fd_sc_hs__a31oi_2_1/a_114_74# fine_freq_track_1/sky130_fd_sc_hs__o21a_1_71/a_376_387#
+ fine_freq_track_1/sky130_fd_sc_hs__nand2_4_3/a_27_74# fine_freq_track_1/sky130_fd_sc_hs__dfxtp_2_11/a_538_429#
+ fine_freq_track_1/sky130_fd_sc_hs__fa_2_5/a_27_378# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_1/a_714_127#
+ fine_freq_track_1/sky130_fd_sc_hs__o21a_1_17/a_83_244# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_17/a_910_118#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_3/D fine_freq_track_1/sky130_fd_sc_hs__nor2_1_47/a_116_368#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_9/a_1224_74# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_65/a_37_78#
+ fine_freq_track_1/sky130_fd_sc_hs__o21a_1_61/a_83_244# fine_freq_track_1/sky130_fd_sc_hs__a22o_1_13/a_230_79#
+ fine_freq_track_1/sky130_fd_sc_hs__nor2_1_87/a_116_368# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_3/a_796_463#
+ fine_freq_track_1/sky130_fd_sc_hs__nand4_1_1/a_373_74# fine_freq_track_1/sky130_fd_sc_hs__dfstp_2_5/a_1356_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_21/Q_N fine_freq_track_1/sky130_fd_sc_hs__nand2_1_17/a_117_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfstp_2_5/a_1521_508# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_45/a_1934_94#
+ fine_freq_track_1/sky130_fd_sc_hs__nor2_1_89/Y fine_freq_track_1/sky130_fd_sc_hs__dfxtp_2_11/a_1019_424#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_49/a_812_138# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_87/a_124_78#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_27/a_856_304# fine_freq_track_1/sky130_fd_sc_hs__o31ai_1_5/a_119_368#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_27/a_850_127# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_89/a_812_138#
+ fine_freq_track_1/sky130_fd_sc_hs__fa_2_5/a_701_79# fine_freq_track_1/sky130_fd_sc_hs__nand2_1_61/a_117_74#
+ fine_freq_track_1/sky130_fd_sc_hs__o21a_1_77/a_320_74# fine_freq_track_1/sky130_fd_sc_hs__nor3_1_3/C
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_53/a_124_78# fine_freq_track_1/sky130_fd_sc_hs__xnor2_1_9/a_138_385#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_23/a_1647_81# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_29/a_1827_81#
+ fine_freq_track_1/sky130_fd_sc_hs__dfxtp_2_9/a_695_459# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_25/a_714_127#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_5/a_832_118# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_51/a_1627_493#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_67/a_1827_81# fine_freq_track_1/sky130_fd_sc_hs__dfxtp_2_1/a_1125_508#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_59/a_789_463# fine_freq_track_1/sky130_fd_sc_hs__fa_2_19/a_27_79#
+ fine_freq_track_1/sky130_fd_sc_hs__sdlclkp_1_1/a_566_74# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_41/a_498_360#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_39/a_1736_119# fine_freq_track_1/sky130_fd_sc_hs__sdlclkp_1_1/a_318_74#
+ fine_freq_track_1/sky130_fd_sc_hs__o21ai_1_5/Y fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_41/a_1350_392#
+ fine_freq_track_1/sky130_fd_sc_hs__a22o_1_11/a_222_392# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_39/a_1266_119#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_11/a_1547_508# fine_freq_track_1/sky130_fd_sc_hs__clkbuf_8_1/a_125_368#
+ fine_freq_track_1/sky130_fd_sc_hs__fa_2_21/a_1119_79# fine_freq_track_1/sky130_fd_sc_hs__dfsbp_2_1/a_595_97#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_21/a_33_74# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_79/a_834_355#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_53/a_494_366# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_19/a_1627_493#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_71/a_2010_409# fine_freq_track_1/sky130_fd_sc_hs__dfxtp_2_11/a_27_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_19/a_37_78# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_35/a_1482_48#
+ fine_freq_track_1/sky130_fd_sc_hs__dfsbp_2_1/a_1453_118# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_29/a_832_118#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_23/a_890_138# fine_freq_track_1/sky130_fd_sc_hs__dfxtp_4_9/a_651_503#
+ fine_freq_track_1/sky130_fd_sc_hs__a21oi_1_93/Y fine_freq_track_1/sky130_fd_sc_hs__o21a_1_61/a_376_387#
+ fine_freq_track_1/sky130_fd_sc_hs__nor3_1_5/B fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_23/a_2026_424#
+ fine_freq_track_1/sky130_fd_sc_hs__dfsbp_2_1/a_731_97# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_7/a_1627_493#
+ fine_freq_track_1/sky130_fd_sc_hs__fa_2_3/a_1094_347# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_9/a_125_78#
+ fine_freq_track_1/sky130_fd_sc_hs__nor2_1_81/Y fine_freq_track_1/sky130_fd_sc_hs__nor2_1_77/a_116_368#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_39/a_2010_409# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_21/a_120_74#
+ fine_freq_track_1/sky130_fd_sc_hs__a21oi_1_41/a_117_74# fine_freq_track_1/sky130_fd_sc_hs__fa_2_5/a_484_347#
+ fine_freq_track_1/sky130_fd_sc_hs__a211oi_1_3/a_354_368# fine_freq_track_1/sky130_fd_sc_hs__fa_2_9/a_27_378#
+ fine_freq_track_1/sky130_fd_sc_hs__a32oi_1_1/a_469_74# fine_freq_track_1/sky130_fd_sc_hs__o21ai_2_1/a_27_74#
+ fine_freq_track_1/sky130_fd_sc_hs__xnor2_1_7/a_376_368# fine_freq_track_1/sky130_fd_sc_hs__dfstp_2_4/a_1521_508#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_31/a_1624_74# fine_freq_track_1/sky130_fd_sc_hs__o21a_1_9/a_320_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_35/a_1934_94# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_91/a_313_74#
+ fine_freq_track_1/sky130_fd_sc_hs__fa_2_3/SUM fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_19/a_1550_119#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_17/a_856_304# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_13/a_125_78#
+ fine_freq_track_1/sky130_fd_sc_hs__a222o_1_1/a_32_74# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_17/a_850_127#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_79/a_812_138# fine_freq_track_1/sky130_fd_sc_hs__o21a_1_65/a_83_244#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_91/a_1350_392# fine_freq_track_1/sky130_fd_sc_hs__nand2_1_101/a_117_74#
+ fine_freq_track_1/sky130_fd_sc_hs__nand4_1_5/a_373_74# fine_freq_track_1/sky130_fd_sc_hs__o211ai_1_11/a_116_368#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_13/a_1647_81# fine_freq_track_1/sky130_fd_sc_hs__dfsbp_2_1/a_27_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_19/a_1827_81# fine_freq_track_1/sky130_fd_sc_hs__fa_2_23/a_487_79#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_15/a_714_127# fine_freq_track_1/sky130_fd_sc_hs__dfstp_2_7/a_1266_341#
+ fine_freq_track_1/sky130_fd_sc_hs__dfstp_2_5/a_612_74# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_37/a_507_368#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_9/a_817_508# fine_freq_track_1/sky130_fd_sc_hs__nand2_1_97/a_117_74#
+ fine_freq_track_1/sky130_fd_sc_hs__conb_1_3/a_165_290# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_91/a_1647_81#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_69/a_1627_493# fine_freq_track_1/sky130_fd_sc_hs__dfsbp_2_1/a_1001_74#
+ fine_freq_track_1/sky130_fd_sc_hs__nor2b_1_33/a_27_112# fine_freq_track_1/sky130_fd_sc_hs__nor2_4_1/a_27_368#
+ fine_freq_track_1/sky130_fd_sc_hs__fa_2_9/a_701_79# fine_freq_track_1/sky130_fd_sc_hs__nand2_1_65/a_117_74#
+ fine_freq_track_1/sky130_fd_sc_hs__xor2_1_3/a_158_392# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_39/a_706_463#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_59/a_1350_392# fine_freq_track_1/sky130_fd_sc_hs__or3b_2_1/a_27_368#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_69/a_834_355# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_29/a_1547_508#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_1/a_1934_94# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_55/a_1678_395#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_3/a_1598_93# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_17/a_1627_493#
+ fine_freq_track_1/sky130_fd_sc_hs__a22oi_1_1/a_159_74# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_83/a_494_366#
+ fine_freq_track_1/sky130_fd_sc_hs__o211ai_1_3/a_116_368# fine_freq_track_1/sky130_fd_sc_hs__o21a_1_15/a_320_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_5/a_841_401# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_7/a_1624_74#
+ fine_freq_track_1/sky130_fd_sc_hs__fa_2_15/a_1202_368# fine_freq_track_1/sky130_fd_sc_hs__dfxtp_4_7/a_206_368#
+ fine_freq_track_1/sky130_fd_sc_hs__o21a_1_11/a_376_387# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_19/a_832_118#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_89/a_2010_409# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_13/a_890_138#
+ fine_freq_track_1/sky130_fd_sc_hs__a21oi_1_15/a_29_368# fine_freq_track_1/sky130_fd_sc_hs__o21a_1_51/a_376_387#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_15/D fine_freq_track_1/sky130_fd_sc_hs__xnor2_1_15/a_376_368#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_1/a_37_78# fine_freq_track_1/sky130_fd_sc_hs__fa_2_9/a_336_347#
+ fine_freq_track_1/sky130_fd_sc_hs__o211ai_1_11/a_31_74# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_91/a_890_138#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_37/a_910_118# fine_freq_track_1/sky130_fd_sc_hs__nor2_1_27/a_116_368#
+ fine_freq_track_1/sky130_fd_sc_hs__nand2_2_7/B fine_freq_track_1/sky130_fd_sc_hs__nor2_1_67/a_116_368#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_27/a_699_463# fine_freq_track_1/sky130_fd_sc_hs__fa_2_7/COUT
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_59/a_37_78# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_37/a_2010_409#
+ fine_freq_track_1/sky130_fd_sc_hs__dfxtp_4_3/a_1034_424# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_29/a_841_401#
+ fine_freq_track_1/sky130_fd_sc_hs__a22o_1_29/a_132_392# fine_freq_track_1/sky130_fd_sc_hs__nor3_1_5/C
+ fine_freq_track_1/sky130_fd_sc_hs__fa_2_19/a_336_347# fine_freq_track_1/sky130_fd_sc_hs__dfstp_2_1/a_1521_508#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_25/a_1934_94# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_21/a_1624_74#
+ fine_freq_track_1/sky130_fd_sc_hs__a22o_1_13/a_52_123# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_5/a_33_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_69/a_812_138# fine_freq_track_1/sky130_fd_sc_hs__a21oi_1_77/a_117_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_13/a_38_78# fine_freq_track_1/sky130_fd_sc_hs__a21oi_1_45/a_117_74#
+ fine_freq_track_1/sky130_fd_sc_hs__a32oi_1_5/a_469_74# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_17/a_313_74#
+ fine_freq_track_1/sky130_fd_sc_hs__fa_2_1/a_683_347# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_47/a_1827_81#
+ fine_freq_track_1/sky130_fd_sc_hs__a21oi_1_11/a_117_74# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_81/a_1647_81#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_39/a_789_463# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_41/a_1224_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_87/a_1827_81# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_67/a_1627_493#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_17/a_125_78# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_73/a_37_78#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_45/a_796_463# fine_freq_track_1/sky130_fd_sc_hs__o22ai_1_7/a_27_74#
+ fine_freq_track_1/sky130_fd_sc_hs__o21a_1_69/a_83_244# fine_freq_track_1/sky130_fd_sc_hs__o211ai_1_3/a_31_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_3/a_910_118# fine_freq_track_1/sky130_fd_sc_hs__nand2_1_105/a_117_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfxtp_2_5/a_644_504# fine_freq_track_1/sky130_fd_sc_hs__o21a_1_35/a_83_244#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_59/a_834_355# fine_freq_track_1/sky130_fd_sc_hs__fa_2_11/a_683_347#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_9/a_494_366# fine_freq_track_1/sky130_fd_sc_hs__dfstp_2_7/a_612_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_53/a_1678_395# fine_freq_track_1/sky130_fd_sc_hs__o21ai_1_1/a_162_368#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_13/a_922_127# fine_freq_track_1/sky130_fd_sc_hs__nor2b_1_9/Y
+ fine_freq_track_1/sky130_fd_sc_hs__nor2b_1_37/a_27_112# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_3/a_38_78#
+ fine_freq_track_1/sky130_fd_sc_hs__a22o_1_5/a_132_392# fine_freq_track_1/sky130_fd_sc_hs__nand2_1_69/a_117_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfxtp_4_7/a_437_503# fine_freq_track_1/sky130_fd_sc_hs__o21a_1_41/a_376_387#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_47/a_832_118# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_29/a_124_78#
+ fine_freq_track_1/sky130_fd_sc_hs__fa_2_9/a_1202_368# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_81/a_890_138#
+ fine_freq_track_1/sky130_fd_sc_hs__fa_2_5/a_27_79# fine_freq_track_1/sky130_fd_sc_hs__fa_2_1/a_1094_347#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_5/a_1627_493# fine_freq_track_1/sky130_fd_sc_hs__o21a_1_19/a_320_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfxtp_4_5/a_735_102# fine_freq_track_1/sky130_fd_sc_hs__a21oi_1_123/a_117_74#
+ fine_freq_track_1/sky130_fd_sc_hs__nor2_1_57/a_116_368# fine_freq_track_1/sky130_fd_sc_hs__a21oi_1_19/a_29_368#
+ fine_freq_track_1/sky130_fd_sc_hs__o21a_1_63/a_320_74# fine_freq_track_1/sky130_fd_sc_hs__dfxtp_4_2/a_1034_424#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_19/a_841_401# fine_freq_track_1/sky130_fd_sc_hs__a22o_1_19/a_132_392#
+ fine_freq_track_1/sky130_fd_sc_hs__o31ai_1_5/a_203_368# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_15/a_1934_94#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_11/a_1624_74# fine_freq_track_1/sky130_fd_sc_hs__dfstp_2_4/a_398_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_17/a_1550_119# fine_freq_track_1/sky130_fd_sc_hs__nor2b_1_17/Y
+ fine_freq_track_1/sky130_fd_sc_hs__a21oi_1_63/a_29_368# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_59/a_812_138#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_37/a_856_304# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_5/a_1434_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_37/a_850_127# fine_freq_track_1/sky130_fd_sc_hs__dfxtp_4_7/a_27_74#
+ fine_freq_track_1/sky130_fd_sc_hs__nand2_2_11/a_27_74# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_7/a_1647_81#
+ fine_freq_track_1/sky130_fd_sc_hs__nand2_2_1/a_27_74# fine_freq_track_1/sky130_fd_sc_hs__fa_2_5/a_1205_79#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_37/a_1827_81# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_3/a_1827_81#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_39/D fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_29/a_789_463#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_71/a_1647_81# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_77/a_1827_81#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_37/a_1736_119# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_41/Q_N
+ fine_freq_track_1/sky130_fd_sc_hs__o31ai_1_1/a_114_74# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_67/a_789_463#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_37/a_1266_119# fine_freq_track_1/sky130_fd_sc_hs__dfstp_2_1/a_27_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_33/Q_N fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_29/a_120_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_57/a_1350_392# fine_freq_track_1/sky130_fd_sc_hs__a32oi_1_9/a_469_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_27/a_1547_508# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_23/Q_N
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_15/a_1627_493# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_29/a_1434_74#
+ fine_freq_track_1/sky130_fd_sc_hs__a21oi_1_93/a_117_74# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_43/a_37_78#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_43/a_922_127# fine_freq_track_1/sky130_fd_sc_hs__fa_2_13/a_1202_368#
+ fine_freq_track_1/sky130_fd_sc_hs__a211oi_1_3/a_159_74# fine_freq_track_1/sky130_fd_sc_hs__nand2_1_109/a_117_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_87/a_2010_409# fine_freq_track_1/sky130_fd_sc_hs__o21a_1_31/a_376_387#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_43/a_1482_48# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_33/a_313_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfxtp_2_1/a_206_368# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_7/a_890_138#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_21/a_2026_424# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_71/a_890_138#
+ fine_freq_track_1/sky130_fd_sc_hs__xnor2_1_3/Y fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_33/a_125_78#
+ fine_freq_track_1/sky130_fd_sc_hs__and2_2_3/a_31_74# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_39/a_2026_424#
+ fine_freq_track_1/sky130_fd_sc_hs__nor3_1_1/A fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_1/a_796_463#
+ fine_freq_track_1/sky130_fd_sc_hs__o21a_1_51/a_83_244# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_85/a_699_463#
+ fine_freq_track_1/sky130_fd_sc_hs__dfstp_2_4/a_1356_74# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_47/a_841_401#
+ fine_freq_track_1/sky130_fd_sc_hs__nor2_1_121/a_116_368# fine_freq_track_1/sky130_fd_sc_hs__nor3_1_5/a_198_368#
+ fine_freq_track_1/sky130_fd_sc_hs__a22oi_1_9/a_159_74# fine_freq_track_1/sky130_fd_sc_hs__a22o_1_7/a_222_392#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_9/a_1678_395# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_45/a_1598_93#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_77/a_124_78# fine_freq_track_1/sky130_fd_sc_hs__nand2_1_51/a_117_74#
+ fine_freq_track_1/sky130_fd_sc_hs__o21a_1_67/a_320_74# fine_freq_track_1/sky130_fd_sc_hs__a22oi_1_3/a_339_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_21/a_1647_81# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_9/a_1465_471#
+ fine_freq_track_1/sky130_fd_sc_hs__dfxtp_2_7/a_695_459# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_11/a_124_78#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_19/a_789_463# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_61/a_1647_81#
+ fine_freq_track_1/sky130_fd_sc_hs__fa_2_17/a_27_378# fine_freq_track_1/sky130_fd_sc_hs__a21oi_1_67/a_29_368#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_25/a_796_463# fine_freq_track_1/sky130_fd_sc_hs__nor2_1_57/B
+ fine_freq_track_1/sky130_fd_sc_hs__nand2b_1_1/a_27_112# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_67/a_37_78#
+ fine_freq_track_1/sky130_fd_sc_hs__a21oi_1_33/a_29_368# fine_freq_track_1/sky130_fd_sc_hs__sdlclkp_4_1/a_744_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_39/a_834_355# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_39/a_319_360#
+ fine_freq_track_1/sky130_fd_sc_hs__a32oi_1_3/a_391_74# fine_freq_track_1/sky130_fd_sc_hs__fa_2_13/a_27_79#
+ fine_freq_track_1/sky130_fd_sc_hs__nand4_1_5/D fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_19/a_1434_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_33/a_922_127# fine_freq_track_1/sky130_fd_sc_hs__fa_2_11/a_1202_368#
+ fine_freq_track_1/sky130_fd_sc_hs__fa_2_7/SUM fine_freq_track_1/sky130_fd_sc_hs__xor2_1_11/a_194_125#
+ fine_freq_track_1/sky130_fd_sc_hs__o21a_1_21/a_376_387# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_27/a_832_118#
+ fine_freq_track_1/sky130_fd_sc_hs__dfsbp_2_1/a_706_463# fine_freq_track_1/sky130_fd_sc_hs__fa_2_23/a_1094_347#
+ fine_freq_track_1/sky130_fd_sc_hs__fa_2_17/a_701_79# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_21/a_890_138#
+ fine_freq_track_1/sky130_fd_sc_hs__fa_2_7/a_1202_368# fine_freq_track_1/sky130_fd_sc_hs__dfsbp_2_1/a_1261_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfxtp_2_11/a_1172_124# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_61/a_890_138#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_5/a_313_74# fine_freq_track_1/sky130_fd_sc_hs__nand2_4_9/A
+ fine_freq_track_1/sky130_fd_sc_hs__nor3_1_7/Y fine_freq_track_1/sky130_fd_sc_hs__a21oi_1_97/a_117_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_83/a_37_78# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_57/D
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_27/a_300_74# fine_freq_track_1/sky130_fd_sc_hs__nor2_1_37/a_116_368#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_45/a_910_118# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_35/a_2010_409#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_45/a_120_74# fine_freq_track_1/sky130_fd_sc_hs__nor2_1_75/a_116_368#
+ fine_freq_track_1/sky130_fd_sc_hs__dfxtp_2_5/a_538_429# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_7/a_120_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_1/a_699_463# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_11/a_120_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_75/a_699_463# fine_freq_track_1/sky130_fd_sc_hs__a21oi_1_31/a_117_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_25/a_33_74# fine_freq_track_1/sky130_fd_sc_hs__nor2_1_111/a_116_368#
+ fine_freq_track_1/sky130_fd_sc_hs__o21ai_1_1/a_27_74# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_37/a_125_78#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_35/a_1598_93# fine_freq_track_1/sky130_fd_sc_hs__nor2b_1_41/a_278_368#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_81/a_313_74# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_39/a_812_138#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_1/a_300_74# fine_freq_track_1/sky130_fd_sc_hs__o21a_1_55/a_83_244#
+ fine_freq_track_1/sky130_fd_sc_hs__fa_2_15/a_484_347# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_17/a_1827_81#
+ fine_freq_track_1/sky130_fd_sc_hs__dfstp_2_5/a_1266_341# fine_freq_track_1/sky130_fd_sc_hs__fa_2_13/a_487_79#
+ fine_freq_track_1/sky130_fd_sc_hs__dfxtp_4_9/a_1226_296# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_13/a_714_127#
+ fine_freq_track_1/sky130_fd_sc_hs__nor2_1_15/B fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_51/a_1647_81#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_57/a_1827_81# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_65/a_1627_493#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_9/Q_N fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_7/a_817_508#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_15/a_796_463# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_35/a_1736_119#
+ fine_freq_track_1/sky130_fd_sc_hs__nor3_1_15/B fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_47/a_789_463#
+ fine_freq_track_1/sky130_fd_sc_hs__nor2b_1_23/a_27_112# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_31/a_498_360#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_35/a_1266_119# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_87/a_789_463#
+ fine_freq_track_1/sky130_fd_sc_hs__inv_4_27/Y fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_55/a_1350_392#
+ fine_freq_track_1/sky130_fd_sc_hs__nand2_1_55/a_117_74# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_47/a_38_78#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_29/a_834_355# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_47/a_124_78#
+ fine_freq_track_1/sky130_fd_sc_hs__a22oi_1_7/a_339_74# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_67/a_834_355#
+ fine_freq_track_1/sky130_fd_sc_hs__fa_2_21/a_683_347# fine_freq_track_1/sky130_fd_sc_hs__o21a_1_37/a_320_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_51/a_1678_395# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_43/a_494_366#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_23/a_922_127# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_1/a_1598_93#
+ fine_freq_track_1/sky130_fd_sc_hs__a22oi_1_23/a_71_368# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_47/a_1434_74#
+ fine_freq_track_1/sky130_fd_sc_hs__nand2b_1_5/a_27_112# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_85/a_2010_409#
+ fine_freq_track_1/sky130_fd_sc_hs__a21oi_1_37/a_29_368# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_23/a_1482_48#
+ fine_freq_track_1/sky130_fd_sc_hs__xnor2_1_7/a_112_119# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_17/a_832_118#
+ fine_freq_track_1/sky130_fd_sc_hs__a32oi_1_7/a_391_74# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_51/a_890_138#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_3/a_1627_493# fine_freq_track_1/sky130_fd_sc_hs__a21oi_1_83/a_29_368#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_19/a_1678_395# fine_freq_track_1/sky130_fd_sc_hs__nand3b_2_1/a_27_94#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_3/a_507_368# fine_freq_track_1/sky130_fd_sc_hs__fa_2_9/a_992_347#
+ fine_freq_track_1/sky130_fd_sc_hs__dfxtp_4_9/a_696_458# fine_freq_track_1/sky130_fd_sc_hs__o21a_1_7/a_376_387#
+ fine_freq_track_1/sky130_fd_sc_hs__dfxtp_4_2/Q fine_freq_track_1/sky130_fd_sc_hs__a32oi_1_3/a_27_368#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_25/a_699_463# fine_freq_track_1/sky130_fd_sc_hs__nor2b_1_9/a_278_368#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_7/a_498_360# fine_freq_track_1/sky130_fd_sc_hs__or3b_2_1/a_190_260#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_65/a_699_463# fine_freq_track_1/sky130_fd_sc_hs__nor2_1_101/a_116_368#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_27/a_841_401# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_9/a_313_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_5/a_706_463# fine_freq_track_1/sky130_fd_sc_hs__fa_2_19/a_992_347#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_15/a_1550_119# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_7/a_1678_395#
+ fine_freq_track_1/sky130_fd_sc_hs__nor2b_1_31/a_278_368# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_25/a_1598_93#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_29/a_812_138# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_49/a_120_74#
+ fine_freq_track_1/sky130_fd_sc_hs__maj3_1_3/a_403_136# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_67/a_812_138#
+ fine_freq_track_1/sky130_fd_sc_hs__dfxtp_2_1/a_708_101# fine_freq_track_1/sky130_fd_sc_hs__dfstp_2_5/a_781_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_7/a_1465_471# fine_freq_track_1/sky130_fd_sc_hs__dfstp_2_4/a_1266_341#
+ fine_freq_track_1/sky130_fd_sc_hs__o22ai_1_5/a_340_368# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_41/a_1647_81#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_63/a_1627_493# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_43/a_300_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_43/a_714_127# fine_freq_track_1/sky130_fd_sc_hs__a21oi_1_117/a_29_368#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_37/a_789_463# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_85/a_313_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_3/a_789_463# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_21/a_498_360#
+ fine_freq_track_1/sky130_fd_sc_hs__nor3_1_15/a_114_368# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_77/a_789_463#
+ fine_freq_track_1/sky130_fd_sc_hs__xnor2_1_15/a_112_119# fine_freq_track_1/sky130_fd_sc_hs__o21a_1_59/a_83_244#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_53/a_1350_392# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_29/a_706_463#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_19/a_834_355# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_1/a_910_118#
+ fine_freq_track_1/sky130_fd_sc_hs__dfxtp_2_3/a_644_504# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_25/a_1547_508#
+ fine_freq_track_1/sky130_fd_sc_hs__a21oi_1_91/Y fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_13/a_1627_493#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_33/a_494_366# fine_freq_track_1/sky130_fd_sc_hs__dfstp_2_7/a_1489_118#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_69/a_1678_395# fine_freq_track_1/sky130_fd_sc_hs__nor2b_1_27/a_27_112#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_7/a_33_74# fine_freq_track_1/sky130_fd_sc_hs__a22o_1_23/a_230_79#
+ fine_freq_track_1/sky130_fd_sc_hs__inv_4_25/Y fine_freq_track_1/sky130_fd_sc_hs__nand2_1_59/a_117_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_13/a_1482_48# fine_freq_track_1/sky130_fd_sc_hs__dfxtp_2_3/a_27_74#
+ fine_freq_track_1/sky130_fd_sc_hs__fa_2_21/a_1094_347# fine_freq_track_1/sky130_fd_sc_hs__inv_4_57/Y
+ fine_freq_track_1/sky130_fd_sc_hs__fa_2_5/a_1202_368# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_41/a_890_138#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_19/a_124_78# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_17/a_1678_395#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_37/a_2026_424# fine_freq_track_1/sky130_fd_sc_hs__or2_1_3/a_152_368#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_25/a_910_118# fine_freq_track_1/sky130_fd_sc_hs__o21a_1_55/X
+ fine_freq_track_1/sky130_fd_sc_hs__nor2_1_17/a_116_368# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_33/a_2010_409#
+ fine_freq_track_1/sky130_fd_sc_hs__dfxtp_2_9/a_1019_424# fine_freq_track_1/sky130_fd_sc_hs__nand2b_1_9/a_27_112#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_77/a_37_78# fine_freq_track_1/sky130_fd_sc_hs__nor2b_1_5/Y
+ fine_freq_track_1/sky130_fd_sc_hs__a21oi_1_113/a_117_74# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_15/a_699_463#
+ fine_freq_track_1/sky130_fd_sc_hs__o211ai_1_5/a_31_74# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_55/a_699_463#
+ fine_freq_track_1/sky130_fd_sc_hs__nor2_1_95/a_116_368# fine_freq_track_1/sky130_fd_sc_hs__o21a_1_53/a_320_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_17/a_841_401# fine_freq_track_1/sky130_fd_sc_hs__nor2b_1_15/Y
+ fine_freq_track_1/sky130_fd_sc_hs__dfstp_2_7/a_1057_118# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_13/a_1550_119#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_13/a_1934_94# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_15/a_1598_93#
+ fine_freq_track_1/sky130_fd_sc_hs__nor2b_1_21/a_278_368# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_17/Q_N
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_19/a_812_138# fine_freq_track_1/sky130_fd_sc_hs__a32oi_1_7/a_27_368#
+ fine_freq_track_1/sky130_fd_sc_hs__dfstp_2_1/a_1266_341# fine_freq_track_1/sky130_fd_sc_hs__dfxtp_4_7/a_1226_296#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_31/a_1647_81# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_33/a_1736_119#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_33/a_714_127# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_31/a_1224_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_11/a_498_360# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_33/a_1266_119#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_35/a_796_463# fine_freq_track_1/sky130_fd_sc_hs__o22ai_1_5/a_142_368#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_19/a_706_463# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_19/a_120_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfstp_2_7/a_781_74# fine_freq_track_1/sky130_fd_sc_hs__a21oi_1_39/a_117_74#
+ fine_freq_track_1/sky130_fd_sc_hs__a2bb2oi_1_1/a_399_368# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_47/a_834_355#
+ fine_freq_track_1/sky130_fd_sc_hs__o21ai_1_11/a_162_368# fine_freq_track_1/sky130_fd_sc_hs__fa_2_15/a_1205_79#
+ fine_freq_track_1/sky130_fd_sc_hs__o21a_1_3/a_83_244# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_23/a_494_366#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_87/a_834_355# fine_freq_track_1/sky130_fd_sc_hs__xor2_1_3/a_194_125#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_67/a_1678_395# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_89/a_313_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_27/a_1434_74# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_41/a_922_127#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_13/a_300_74# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_83/a_2010_409#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_3/a_856_304# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_3/a_850_127#
+ fine_freq_track_1/sky130_fd_sc_hs__nand2_2_13/a_27_74# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_37/a_832_118#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_23/a_313_74# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_31/a_890_138#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_1/a_1627_493# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_15/a_910_118#
+ fine_freq_track_1/sky130_fd_sc_hs__dfxtp_2_7/a_1019_424# fine_freq_track_1/sky130_fd_sc_hs__nor2b_1_3/a_27_112#
+ fine_freq_track_1/sky130_fd_sc_hs__a22o_1_27/a_230_79# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_7/a_1224_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_45/a_699_463# fine_freq_track_1/sky130_fd_sc_hs__o21a_1_41/a_83_244#
+ fine_freq_track_1/sky130_fd_sc_hs__nor2_1_85/a_116_368# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_9/a_1350_392#
+ fine_freq_track_1/sky130_fd_sc_hs__dfxtp_2_11/a_1217_314# fine_freq_track_1/sky130_fd_sc_hs__dfstp_2_1/a_1356_74#
+ fine_freq_track_1/sky130_fd_sc_hs__nand4_2_1/a_27_74# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_3/a_124_78#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_5/a_1678_395# fine_freq_track_1/sky130_fd_sc_hs__nor2b_1_11/a_278_368#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_43/a_1934_94# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_77/D
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_47/a_812_138# fine_freq_track_1/sky130_fd_sc_hs__dfxtp_2_9/a_431_508#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_87/a_812_138# fine_freq_track_1/sky130_fd_sc_hs__dfstp_2_4/a_225_74#
+ fine_freq_track_1/sky130_fd_sc_hs__o21a_1_57/a_320_74# fine_freq_track_1/sky130_fd_sc_hs__a32oi_1_3/a_119_74#
+ fine_freq_track_1/sky130_fd_sc_hs__xnor2_1_7/a_138_385# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_27/a_1827_81#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_23/a_714_127# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_31/a_1736_119#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_3/a_832_118# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_17/a_789_463#
+ fine_freq_track_1/sky130_fd_sc_hs__a2bb2oi_1_1/a_488_74# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_21/a_1224_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_45/a_507_368# fine_freq_track_1/sky130_fd_sc_hs__a21oi_1_57/a_29_368#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_31/a_1266_119# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_57/a_789_463#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_23/a_1547_508# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_47/a_706_463#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_37/a_834_355# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_11/a_1627_493#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_13/a_494_366# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_3/a_834_355#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_77/a_834_355# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_61/a_37_78#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_17/a_1434_74# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_31/a_922_127#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_91/a_494_366# fine_freq_track_1/sky130_fd_sc_hs__a2bb2oi_1_1/a_126_112#
+ fine_freq_track_1/sky130_fd_sc_hs__xnor2_1_3/a_293_74# fine_freq_track_1/sky130_fd_sc_hs__fa_2_3/a_1202_368#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_33/a_1482_48# fine_freq_track_1/sky130_fd_sc_hs__dfxtp_4_7/a_651_503#
+ fine_freq_track_1/sky130_fd_sc_hs__o21a_1_7/a_83_244# fine_freq_track_1/sky130_fd_sc_hs__a22o_1_23/a_52_123#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_15/a_1678_395# fine_freq_track_1/sky130_fd_sc_hs__dfxtp_4_9/a_544_485#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_35/a_2026_424# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_31/a_2010_409#
+ fine_freq_track_1/sky130_fd_sc_hs__a21oi_1_87/a_117_74# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_39/a_817_508#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_19/a_1465_471# fine_freq_track_1/sky130_fd_sc_hs__a222oi_1_1/a_461_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_17/a_300_74# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_35/a_120_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_49/a_2010_409# fine_freq_track_1/sky130_fd_sc_hs__a21oi_1_53/a_117_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_35/a_699_463# fine_freq_track_1/sky130_fd_sc_hs__dfxtp_2_3/a_538_429#
+ fine_freq_track_1/sky130_fd_sc_hs__xnor2_1_15/a_138_385# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_27/a_313_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_73/a_699_463# fine_freq_track_1/sky130_fd_sc_hs__fa_2_3/a_484_347#
+ fine_freq_track_1/sky130_fd_sc_hs__a21oi_1_21/a_117_74# fine_freq_track_1/sky130_fd_sc_hs__a211oi_1_1/a_354_368#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_11/a_1550_119# fine_freq_track_1/sky130_fd_sc_hs__o2bb2ai_1_1/a_397_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_37/a_841_401# fine_freq_track_1/sky130_fd_sc_hs__o21ai_2_1/a_116_368#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_39/a_1624_74# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_5/a_319_360#
+ fine_freq_track_1/sky130_fd_sc_hs__xnor2_1_5/a_376_368# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_33/a_1934_94#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_71/a_313_74# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_37/a_812_138#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_19/D fine_freq_track_1/sky130_fd_sc_hs__a21oi_1_3/a_117_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_3/a_812_138# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_25/a_38_78#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_77/a_812_138# fine_freq_track_1/sky130_fd_sc_hs__o21a_1_45/a_83_244#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_5/a_1465_471# fine_freq_track_1/sky130_fd_sc_hs__dfxtp_4_5/a_1226_296#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_11/a_1647_81# fine_freq_track_1/sky130_fd_sc_hs__fa_2_9/a_1119_79#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_61/a_1627_493# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_9/a_1482_48#
+ fine_freq_track_1/sky130_fd_sc_hs__o21a_1_11/a_83_244# fine_freq_track_1/sky130_fd_sc_hs__nor2b_2_1/a_27_392#
+ fine_freq_track_1/sky130_fd_sc_hs__o21a_1_1/a_320_74# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_11/a_1224_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_35/a_507_368# fine_freq_track_1/sky130_fd_sc_hs__conb_1_1/a_165_290#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_51/a_1350_392# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_21/a_1547_508#
+ fine_freq_track_1/sky130_fd_sc_hs__xor2_1_1/a_158_392# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_37/a_124_78#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_29/a_319_360# fine_freq_track_1/sky130_fd_sc_hs__a32oi_1_7/a_119_74#
+ fine_freq_track_1/sky130_fd_sc_hs__fa_2_19/a_1119_79# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_27/a_33_74#
+ fine_freq_track_1/sky130_fd_sc_hs__o21a_1_27/a_320_74# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_29/a_1627_493#
+ fine_freq_track_1/sky130_fd_sc_hs__dfstp_2_7/a_1596_118# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_21/a_922_127#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_81/a_494_366# fine_freq_track_1/sky130_fd_sc_hs__o211ai_1_1/a_116_368#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_81/a_2010_409# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_3/a_841_401#
+ fine_freq_track_1/sky130_fd_sc_hs__a22oi_1_13/a_71_368# fine_freq_track_1/sky130_fd_sc_hs__dfxtp_4_5/a_206_368#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_19/a_1350_392# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_79/D
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_11/a_890_138# fine_freq_track_1/sky130_fd_sc_hs__xnor2_1_13/a_376_368#
+ fine_freq_track_1/sky130_fd_sc_hs__fa_2_23/a_27_378# fine_freq_track_1/sky130_fd_sc_hs__fa_2_7/a_336_347#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_1/a_507_368# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_17/a_1465_471#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_29/a_817_508# fine_freq_track_1/sky130_fd_sc_hs__dfstp_2_7/a_1566_92#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_35/a_910_118# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_7/a_1350_392#
+ fine_freq_track_1/sky130_fd_sc_hs__nor2_1_65/a_116_368# fine_freq_track_1/sky130_fd_sc_hs__xnor2_1_7/a_293_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_43/a_33_74# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_63/a_699_463#
+ fine_freq_track_1/sky130_fd_sc_hs__a22o_1_27/a_52_123# fine_freq_track_1/sky130_fd_sc_hs__maj3_1_3/a_406_384#
+ fine_freq_track_1/sky130_fd_sc_hs__a22o_1_27/a_132_392# fine_freq_track_1/sky130_fd_sc_hs__fa_2_17/a_336_347#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_23/a_1934_94# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_29/a_1550_119#
+ fine_freq_track_1/sky130_fd_sc_hs__maj3_1_1/a_403_136# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_45/a_856_304#
+ fine_freq_track_1/sky130_fd_sc_hs__fa_2_23/a_701_79# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_45/a_850_127#
+ fine_freq_track_1/sky130_fd_sc_hs__a21oi_1_25/a_117_74# fine_freq_track_1/sky130_fd_sc_hs__sdlclkp_1_1/a_667_80#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_33/a_300_74# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_25/a_507_368#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_79/a_1627_493# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_41/a_714_127#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_5/a_125_78# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_49/a_1736_119#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_75/a_313_74# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_47/Q_N
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_85/a_1827_81# fine_freq_track_1/sky130_fd_sc_hs__xor2_1_9/a_355_368#
+ fine_freq_track_1/sky130_fd_sc_hs__a21oi_1_7/a_117_74# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_43/a_796_463#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_49/a_1266_119# fine_freq_track_1/sky130_fd_sc_hs__o21a_1_49/a_83_244#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_69/a_1350_392# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_27/a_706_463#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_17/a_834_355# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_19/a_319_360#
+ fine_freq_track_1/sky130_fd_sc_hs__a22o_1_3/a_230_79# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_39/a_1547_508#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_57/a_834_355# fine_freq_track_1/sky130_fd_sc_hs__dfstp_2_5/a_1489_118#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_41/a_125_78# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_65/a_1678_395#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_7/a_494_366# fine_freq_track_1/sky130_fd_sc_hs__o21a_1_5/a_320_74#
+ fine_freq_track_1/sky130_fd_sc_hs__nor2b_1_49/a_27_112# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_11/a_922_127#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_71/a_494_366# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_55/a_37_78#
+ fine_freq_track_1/sky130_fd_sc_hs__and2_2_3/a_118_74# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_37/a_1434_74#
+ fine_freq_track_1/sky130_fd_sc_hs__nor2b_1_17/a_27_112# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_17/a_1350_392#
+ fine_freq_track_1/sky130_fd_sc_hs__a22o_1_3/a_132_392# fine_freq_track_1/sky130_fd_sc_hs__nand2_1_49/a_117_74#
+ fine_freq_track_1/sky130_fd_sc_hs__fa_2_1/a_1202_368# fine_freq_track_1/sky130_fd_sc_hs__a222o_1_1/a_119_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfxtp_4_5/a_437_503# fine_freq_track_1/sky130_fd_sc_hs__conb_1_3/LO
+ fine_freq_track_1/sky130_fd_sc_hs__nor2b_2_1/a_228_368# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_45/a_832_118#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_33/a_2026_424# fine_freq_track_1/sky130_fd_sc_hs__nand2_1_93/a_117_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfxtp_2_5/a_1019_424# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_19/a_817_508#
+ fine_freq_track_1/sky130_fd_sc_hs__a22oi_1_17/a_71_368# fine_freq_track_1/sky130_fd_sc_hs__sdlclkp_1_1/a_116_424#
+ fine_freq_track_1/sky130_fd_sc_hs__nand2_1_9/a_117_74# fine_freq_track_1/sky130_fd_sc_hs__nor3_1_9/a_114_368#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_47/a_2010_409# fine_freq_track_1/sky130_fd_sc_hs__a21oi_1_103/a_117_74#
+ fine_freq_track_1/sky130_fd_sc_hs__nor2_1_55/a_116_368# fine_freq_track_1/sky130_fd_sc_hs__a2bb2oi_1_1/a_117_392#
+ fine_freq_track_1/sky130_fd_sc_hs__nor2_1_53/Y fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_53/a_699_463#
+ fine_freq_track_1/sky130_fd_sc_hs__dfstp_2_5/a_1057_118# fine_freq_track_1/sky130_fd_sc_hs__o21a_1_43/a_320_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_3/a_1678_395# fine_freq_track_1/sky130_fd_sc_hs__a22o_1_17/a_132_392#
+ fine_freq_track_1/sky130_fd_sc_hs__o22ai_1_3/a_27_74# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_13/a_1598_93#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_17/a_812_138# fine_freq_track_1/sky130_fd_sc_hs__nor2b_1_27/Y
+ fine_freq_track_1/sky130_fd_sc_hs__a21oi_1_43/a_29_368# fine_freq_track_1/sky130_fd_sc_hs__nor2_1_13/B
+ fine_freq_track_1/sky130_fd_sc_hs__nor4_1_1/Y fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_57/a_812_138#
+ fine_freq_track_1/sky130_fd_sc_hs__dfxtp_2_11/a_695_459# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_3/a_1465_471#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_35/a_856_304# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_35/a_850_127#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_3/a_1434_74# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_11/a_33_74#
+ fine_freq_track_1/sky130_fd_sc_hs__fa_2_3/a_1205_79# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_5/a_1647_81#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_15/a_507_368# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_31/a_714_127#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_1/a_1827_81# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_27/a_789_463#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_47/a_1736_119# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_75/a_1827_81#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_47/a_1266_119# fine_freq_track_1/sky130_fd_sc_hs__o211ai_1_9/a_31_74#
+ fine_freq_track_1/sky130_fd_sc_hs__nor2_1_5/a_116_368# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_67/a_1350_392#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_17/a_706_463# fine_freq_track_1/sky130_fd_sc_hs__a22o_1_29/a_222_392#
+ fine_freq_track_1/sky130_fd_sc_hs__a21oi_1_29/a_117_74# fine_freq_track_1/sky130_fd_sc_hs__fa_2_1/a_27_79#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_47/a_319_360# fine_freq_track_1/sky130_fd_sc_hs__dfstp_2_4/a_1489_118#
+ fine_freq_track_1/sky130_fd_sc_hs__a211oi_4_1/a_77_368# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_21/a_494_366#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_63/a_1678_395# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_27/a_1627_493#
+ fine_freq_track_1/sky130_fd_sc_hs__dfxtp_2_9/a_1172_124# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_37/a_300_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_61/a_494_366# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_79/a_313_74#
+ fine_freq_track_1/sky130_fd_sc_hs__nor2_2_3/A fine_freq_track_1/sky130_fd_sc_hs__a21oi_1_73/a_117_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_35/a_38_78# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_1/a_856_304#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_1/a_850_127# fine_freq_track_1/sky130_fd_sc_hs__a22o_1_7/a_230_79#
+ fine_freq_track_1/sky130_fd_sc_hs__nor2b_1_43/Y fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_41/a_1482_48#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_13/a_1678_395# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_13/a_313_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_45/a_125_78# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_5/a_890_138#
+ fine_freq_track_1/sky130_fd_sc_hs__dfxtp_2_3/a_1019_424# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_15/a_1465_471#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_3/Q_N fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_49/a_817_508#
+ fine_freq_track_1/sky130_fd_sc_hs__a22o_1_17/a_230_79# fine_freq_track_1/sky130_fd_sc_hs__or2_1_1/a_63_368#
+ fine_freq_track_1/sky130_fd_sc_hs__nor2_1_45/a_116_368# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_5/a_1350_392#
+ fine_freq_track_1/sky130_fd_sc_hs__o21a_1_31/a_83_244# fine_freq_track_1/sky130_fd_sc_hs__dfstp_2_4/a_1057_118#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_37/a_33_74# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_83/a_699_463#
+ fine_freq_track_1/sky130_fd_sc_hs__dfstp_2_4/a_612_74# fine_freq_track_1/sky130_fd_sc_hs__a22oi_1_23/a_159_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_45/a_841_401# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_27/a_1550_119#
+ fine_freq_track_1/sky130_fd_sc_hs__nor3_1_3/a_198_368# fine_freq_track_1/sky130_fd_sc_hs__dfxtp_4_9/a_1141_508#
+ fine_freq_track_1/sky130_fd_sc_hs__a22o_1_5/a_222_392# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_41/a_1934_94#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_43/a_1598_93# fine_freq_track_1/sky130_fd_sc_hs__nand2_1_63/a_117_74#
+ fine_freq_track_1/sky130_fd_sc_hs__a21oi_1_107/a_117_74# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_57/a_124_78#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_1/a_1465_471# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_25/a_856_304#
+ fine_freq_track_1/sky130_fd_sc_hs__o31ai_1_3/a_119_368# fine_freq_track_1/sky130_fd_sc_hs__dfxtp_2_7/a_431_508#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_25/a_850_127# fine_freq_track_1/sky130_fd_sc_hs__dfxtp_4_3/a_1226_296#
+ fine_freq_track_1/sky130_fd_sc_hs__nand2_1_31/a_117_74# fine_freq_track_1/sky130_fd_sc_hs__o21a_1_47/a_320_74#
+ fine_freq_track_1/sky130_fd_sc_hs__fa_2_23/a_484_347# fine_freq_track_1/sky130_fd_sc_hs__a21oi_1_79/a_29_368#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_25/a_1827_81# fine_freq_track_1/sky130_fd_sc_hs__nand2_2_7/a_27_74#
+ fine_freq_track_1/sky130_fd_sc_hs__o21a_1_13/a_320_74# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_77/a_1627_493#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_21/a_714_127# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_1/a_832_118#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_65/a_1827_81# fine_freq_track_1/sky130_fd_sc_hs__a21oi_1_47/a_29_368#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_23/a_796_463# fine_freq_track_1/sky130_fd_sc_hs__dfstp_2_5/a_767_384#
+ fine_freq_track_1/sky130_fd_sc_hs__a22o_1_19/a_222_392# fine_freq_track_1/sky130_fd_sc_hs__dfstp_2_7/a_27_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfstp_2_1/a_1489_118# fine_freq_track_1/sky130_fd_sc_hs__a21oi_1_91/a_29_368#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_25/a_1627_493# fine_freq_track_1/sky130_fd_sc_hs__dfxtp_2_7/a_1172_124#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_51/a_494_366# fine_freq_track_1/sky130_fd_sc_hs__fa_2_23/a_1202_368#
+ fine_freq_track_1/sky130_fd_sc_hs__a222o_1_1/a_651_74# fine_freq_track_1/sky130_fd_sc_hs__a22o_1_3/a_52_123#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_15/a_1350_392# fine_freq_track_1/sky130_fd_sc_hs__fa_2_3/a_487_79#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_25/a_832_118# fine_freq_track_1/sky130_fd_sc_hs__o21a_1_69/a_376_387#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_31/a_2026_424# fine_freq_track_1/sky130_fd_sc_hs__nor2_2_3/B
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_43/a_910_118# fine_freq_track_1/sky130_fd_sc_hs__nor2_1_35/a_116_368#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_49/a_313_74# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_25/a_120_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_9/a_699_463# fine_freq_track_1/sky130_fd_sc_hs__nor2_1_73/a_116_368#
+ fine_freq_track_1/sky130_fd_sc_hs__dfstp_2_1/a_1057_118# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_1/a_1678_395#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_17/D fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_63/a_37_78#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_9/a_922_127# fine_freq_track_1/sky130_fd_sc_hs__nor2b_1_49/a_278_368#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_31/a_1934_94# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_33/a_1598_93#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_61/a_313_74# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_15/a_856_304#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_15/a_850_127# fine_freq_track_1/sky130_fd_sc_hs__dfxtp_4_2/a_1226_296#
+ fine_freq_track_1/sky130_fd_sc_hs__o21a_1_39/X fine_freq_track_1/sky130_fd_sc_hs__fa_2_13/a_484_347#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_15/a_1827_81# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_11/a_714_127#
+ fine_freq_track_1/sky130_fd_sc_hs__nor2b_1_35/a_27_112# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_55/a_1827_81#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_13/a_796_463# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_39/a_498_360#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_85/a_789_463# fine_freq_track_1/sky130_fd_sc_hs__a22oi_1_21/a_339_74#
+ fine_freq_track_1/sky130_fd_sc_hs__nand2_1_35/a_117_74# fine_freq_track_1/sky130_fd_sc_hs__o22ai_1_11/a_27_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_37/a_1547_508# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_37/a_706_463#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_27/a_834_355# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_27/a_319_360#
+ fine_freq_track_1/sky130_fd_sc_hs__xnor2_1_13/a_293_74# fine_freq_track_1/sky130_fd_sc_hs__dfstp_2_5/a_1596_118#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_41/a_494_366# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_11/Q_N
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_1/a_841_401# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_45/a_1434_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_5/a_1624_74# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_29/a_38_78#
+ fine_freq_track_1/sky130_fd_sc_hs__xnor2_1_5/a_112_119# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_15/a_832_118#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_11/a_1678_395# fine_freq_track_1/sky130_fd_sc_hs__a21oi_1_95/a_29_368#
+ fine_freq_track_1/sky130_fd_sc_hs__o21a_1_59/a_376_387# fine_freq_track_1/sky130_fd_sc_hs__dfxtp_2_1/a_1019_424#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_13/a_1465_471# fine_freq_track_1/sky130_fd_sc_hs__dfstp_2_1/a_398_74#
+ fine_freq_track_1/sky130_fd_sc_hs__fa_2_13/a_27_378# fine_freq_track_1/sky130_fd_sc_hs__fa_2_7/a_992_347#
+ fine_freq_track_1/sky130_fd_sc_hs__o21a_1_69/X fine_freq_track_1/sky130_fd_sc_hs__dfxtp_4_7/a_696_458#
+ fine_freq_track_1/sky130_fd_sc_hs__a22o_1_7/a_52_123# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_45/a_2010_409#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_89/a_37_78# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_17/a_37_78#
+ fine_freq_track_1/sky130_fd_sc_hs__nor2_1_25/a_116_368# fine_freq_track_1/sky130_fd_sc_hs__o21a_1_5/a_376_387#
+ fine_freq_track_1/sky130_fd_sc_hs__fa_2_7/a_487_79# fine_freq_track_1/sky130_fd_sc_hs__fa_2_17/SUM
+ fine_freq_track_1/sky130_fd_sc_hs__nor2b_1_7/a_278_368# fine_freq_track_1/sky130_fd_sc_hs__nor2_1_109/a_116_368#
+ fine_freq_track_1/sky130_fd_sc_hs__a22o_1_17/a_52_123# fine_freq_track_1/sky130_fd_sc_hs__maj3_1_1/a_406_384#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_25/a_841_401# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_3/a_706_463#
+ fine_freq_track_1/sky130_fd_sc_hs__dfxtp_4_7/a_1141_508# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_29/a_1624_74#
+ fine_freq_track_1/sky130_fd_sc_hs__fa_2_17/a_992_347# fine_freq_track_1/sky130_fd_sc_hs__nor2b_1_39/a_278_368#
+ fine_freq_track_1/sky130_fd_sc_hs__o21ai_1_7/a_27_74# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_21/a_1934_94#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_23/a_1598_93# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_27/a_812_138#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_43/a_38_78# fine_freq_track_1/sky130_fd_sc_hs__dfstp_2_7/a_716_456#
+ fine_freq_track_1/sky130_fd_sc_hs__fa_2_13/a_701_79# fine_freq_track_1/sky130_fd_sc_hs__a21oi_1_15/a_117_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_1/a_313_74# fine_freq_track_1/sky130_fd_sc_hs__fa_2_9/a_683_347#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_75/a_1627_493# fine_freq_track_1/sky130_fd_sc_hs__o22ai_1_3/a_340_368#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_49/a_1647_81# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_45/a_1736_119#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_45/a_1827_81# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_33/a_37_78#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_23/a_300_74# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_89/a_1647_81#
+ fine_freq_track_1/sky130_fd_sc_hs__nand4_1_3/a_259_74# fine_freq_track_1/sky130_fd_sc_hs__conb_1_3/HI
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_45/a_1266_119# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_65/a_313_74#
+ fine_freq_track_1/sky130_fd_sc_hs__xor2_1_7/a_355_368# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_1/a_789_463#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_65/a_1350_392# fine_freq_track_1/sky130_fd_sc_hs__nor3_1_13/a_114_368#
+ fine_freq_track_1/sky130_fd_sc_hs__sdlclkp_4_1/a_785_455# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_3/a_120_74#
+ fine_freq_track_1/sky130_fd_sc_hs__xnor2_1_13/a_112_119# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_75/a_789_463#
+ fine_freq_track_1/sky130_fd_sc_hs__o21a_1_39/a_83_244# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_17/a_319_360#
+ fine_freq_track_1/sky130_fd_sc_hs__dfxtp_2_1/a_644_504# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_61/a_1678_395#
+ fine_freq_track_1/sky130_fd_sc_hs__fa_2_19/a_683_347# fine_freq_track_1/sky130_fd_sc_hs__dfstp_2_4/a_1596_118#
+ fine_freq_track_1/sky130_fd_sc_hs__fa_2_23/a_1205_79# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_31/a_494_366#
+ fine_freq_track_1/sky130_fd_sc_hs__fa_2_21/a_1202_368# fine_freq_track_1/sky130_fd_sc_hs__nor2b_1_39/a_27_112#
+ fine_freq_track_1/sky130_fd_sc_hs__o21ai_1_9/a_162_368# fine_freq_track_1/sky130_fd_sc_hs__o21a_1_11/X
+ fine_freq_track_1/sky130_fd_sc_hs__a22oi_1_25/a_339_74# fine_freq_track_1/sky130_fd_sc_hs__nand2_1_39/a_117_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfsbp_2_1/a_398_74# fine_freq_track_1/sky130_fd_sc_hs__o21a_1_49/a_376_387#
+ fine_freq_track_1/sky130_fd_sc_hs__dfxtp_2_9/a_1217_314# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_49/a_890_138#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_29/a_1678_395# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_47/a_2026_424#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_89/a_890_138# fine_freq_track_1/sky130_fd_sc_hs__nand2_1_83/a_117_74#
+ fine_freq_track_1/sky130_fd_sc_hs__or2_1_1/a_152_368# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_23/a_910_118#
+ fine_freq_track_1/sky130_fd_sc_hs__nor2_1_15/a_116_368# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_3/a_1350_392#
+ fine_freq_track_1/sky130_fd_sc_hs__dfxtp_4_3/a_735_102# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_43/a_124_78#
+ fine_freq_track_1/sky130_fd_sc_hs__a21oi_1_99/a_29_368# fine_freq_track_1/sky130_fd_sc_hs__nor2_1_93/a_116_368#
+ fine_freq_track_1/sky130_fd_sc_hs__o21a_1_33/a_320_74# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_15/a_841_401#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_25/a_1550_119# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_19/a_1624_74#
+ fine_freq_track_1/sky130_fd_sc_hs__o31ai_1_3/a_203_368# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_11/a_1934_94#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_9/a_1736_119# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_1/a_1434_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_9/a_1266_119# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_73/a_1627_493#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_35/a_1827_81# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_13/a_507_368#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_79/a_1647_81# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_39/a_1224_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_9/a_37_78# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_25/a_789_463#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_73/a_1827_81# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_63/a_1350_392#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_33/a_796_463# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_65/a_789_463#
+ fine_freq_track_1/sky130_fd_sc_hs__dfstp_2_5/a_2022_94# fine_freq_track_1/sky130_fd_sc_hs__inv_2_9/Y
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_35/a_1547_508# fine_freq_track_1/sky130_fd_sc_hs__o22ai_1_3/a_142_368#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_23/a_1627_493# fine_freq_track_1/sky130_fd_sc_hs__a21oi_1_19/a_117_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfxtp_2_5/a_1172_124# fine_freq_track_1/sky130_fd_sc_hs__dfstp_2_1/a_1596_118#
+ fine_freq_track_1/sky130_fd_sc_hs__fa_2_13/a_1205_79# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_79/a_1678_395#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_85/a_834_355# fine_freq_track_1/sky130_fd_sc_hs__xor2_1_1/a_194_125#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_13/a_1350_392# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_69/a_313_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_25/a_1434_74# fine_freq_track_1/sky130_fd_sc_hs__a21oi_1_63/a_117_74#
+ fine_freq_track_1/sky130_fd_sc_hs__o21a_1_39/a_376_387# fine_freq_track_1/sky130_fd_sc_hs__dfsbp_2_1/a_1258_341#
+ fine_freq_track_1/sky130_fd_sc_hs__dfxtp_2_7/a_1217_314# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_15/a_33_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_35/a_832_118# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_9/a_714_127#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_79/a_890_138# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_1/a_38_78#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_43/a_2010_409# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_13/a_910_118#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_47/a_817_508# fine_freq_track_1/sky130_fd_sc_hs__fa_2_23/SUM
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_9/a_796_463# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_43/a_699_463#
+ fine_freq_track_1/sky130_fd_sc_hs__fa_2_11/a_487_79# fine_freq_track_1/sky130_fd_sc_hs__o21a_1_21/a_83_244#
+ fine_freq_track_1/sky130_fd_sc_hs__nor2_1_83/a_116_368# fine_freq_track_1/sky130_fd_sc_hs__a222oi_1_1/a_697_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfxtp_4_5/a_1141_508# fine_freq_track_1/sky130_fd_sc_hs__a22oi_1_13/a_159_74#
+ fine_freq_track_1/sky130_fd_sc_hs__nand2_1_87/a_117_74# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_47/a_1624_74#
+ fine_freq_track_1/sky130_fd_sc_hs__conb_1_3/a_21_290# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_41/a_1598_93#
+ fine_freq_track_1/sky130_fd_sc_hs__nand2b_1_1/a_269_74# fine_freq_track_1/sky130_fd_sc_hs__a22oi_1_5/a_339_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_7/a_1736_119# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_85/a_812_138#
+ fine_freq_track_1/sky130_fd_sc_hs__nand2_1_21/a_117_74# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_7/a_1266_119#
+ fine_freq_track_1/sky130_fd_sc_hs__xnor2_1_5/a_138_385# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_43/a_1736_119#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_91/a_124_78# fine_freq_track_1/sky130_fd_sc_hs__dfxtp_2_5/a_695_459#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_69/a_1647_81# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_43/a_1266_119#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_15/a_789_463# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_63/a_1827_81#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_27/a_37_78# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_43/a_507_368#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_55/a_789_463# fine_freq_track_1/sky130_fd_sc_hs__dfstp_2_4/a_767_384#
+ fine_freq_track_1/sky130_fd_sc_hs__inv_4_15/A fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_21/a_1627_493#
+ fine_freq_track_1/sky130_fd_sc_hs__dfxtp_2_3/a_1172_124# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_45/a_706_463#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_37/a_319_360# fine_freq_track_1/sky130_fd_sc_hs__a21oi_1_82/a_29_368#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_11/a_494_366# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_39/a_33_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_1/a_834_355# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_75/a_834_355#
+ fine_freq_track_1/sky130_fd_sc_hs__nand4_1_1/a_181_74# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_15/a_1434_74#
+ fine_freq_track_1/sky130_fd_sc_hs__o21a_1_29/a_376_387# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_31/a_1482_48#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_11/a_1465_471# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_27/a_1678_395#
+ fine_freq_track_1/sky130_fd_sc_hs__dfxtp_4_5/a_651_503# fine_freq_track_1/sky130_fd_sc_hs__maj3_1_3/a_595_136#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_45/a_2026_424# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_69/a_890_138#
+ fine_freq_track_1/sky130_fd_sc_hs__dfxtp_4_7/a_544_485# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_47/a_120_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_1/a_1350_392# fine_freq_track_1/sky130_fd_sc_hs__a21oi_1_67/a_117_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_15/a_120_74# fine_freq_track_1/sky130_fd_sc_hs__dfstp_2_4/a_781_74#
+ fine_freq_track_1/sky130_fd_sc_hs__a21oi_1_33/a_117_74# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_33/a_699_463#
+ fine_freq_track_1/sky130_fd_sc_hs__xnor2_1_13/a_138_385# fine_freq_track_1/sky130_fd_sc_hs__dfxtp_2_1/a_538_429#
+ fine_freq_track_1/sky130_fd_sc_hs__nand4_2_1/Y fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_23/a_1550_119#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_39/a_125_78# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_41/a_300_74#
+ fine_freq_track_1/sky130_fd_sc_hs__fa_2_1/a_484_347# fine_freq_track_1/sky130_fd_sc_hs__nor2_1_119/a_116_368#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_35/a_841_401# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_5/a_300_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_3/a_319_360# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_7/a_922_127#
+ fine_freq_track_1/sky130_fd_sc_hs__xnor2_1_3/a_376_368# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_13/Q_N
+ fine_freq_track_1/sky130_fd_sc_hs__o211ai_1_11/a_311_74# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_31/a_1598_93#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_51/a_313_74# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_13/a_856_304#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_1/a_812_138# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_75/a_812_138#
+ fine_freq_track_1/sky130_fd_sc_hs__o2bb2ai_1_1/a_490_368# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_13/a_850_127#
+ fine_freq_track_1/sky130_fd_sc_hs__o21a_1_25/a_83_244# fine_freq_track_1/sky130_fd_sc_hs__fa_2_11/a_484_347#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_41/a_1736_119# fine_freq_track_1/sky130_fd_sc_hs__fa_2_7/a_1119_79#
+ fine_freq_track_1/sky130_fd_sc_hs__a22oi_1_17/a_159_74# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_7/a_1482_48#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_59/a_1647_81# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_41/a_1266_119#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_53/a_1827_81# fine_freq_track_1/sky130_fd_sc_hs__a22o_1_21/a_230_79#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_33/a_507_368# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_5/a_817_508#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_45/a_789_463# fine_freq_track_1/sky130_fd_sc_hs__nor4_1_3/a_342_368#
+ fine_freq_track_1/sky130_fd_sc_hs__nand2b_1_5/a_269_74# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_33/a_1547_508#
+ fine_freq_track_1/sky130_fd_sc_hs__a222oi_1_1/a_119_74# fine_freq_track_1/sky130_fd_sc_hs__a22oi_1_11/a_339_74#
+ fine_freq_track_1/sky130_fd_sc_hs__nand2_1_25/a_117_74# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_25/a_834_355#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_17/a_124_78# fine_freq_track_1/sky130_fd_sc_hs__fa_2_17/a_1119_79#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_77/a_1678_395# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_65/a_834_355#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_9/a_1934_94# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_11/a_1350_392#
+ fine_freq_track_1/sky130_fd_sc_hs__o21a_1_19/a_376_387# fine_freq_track_1/sky130_fd_sc_hs__fa_2_11/a_27_79#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_21/a_1482_48# fine_freq_track_1/sky130_fd_sc_hs__nand2_1_15/Y
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_25/a_1678_395# fine_freq_track_1/sky130_fd_sc_hs__a21oi_1_85/a_29_368#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_59/a_890_138# fine_freq_track_1/sky130_fd_sc_hs__xnor2_1_11/a_376_368#
+ fine_freq_track_1/sky130_fd_sc_hs__nand4_1_5/a_181_74# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_41/a_2010_409#
+ fine_freq_track_1/sky130_fd_sc_hs__a22oi_1_3/a_71_368# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_29/a_1465_471#
+ fine_freq_track_1/sky130_fd_sc_hs__a21oi_1_51/a_29_368# fine_freq_track_1/sky130_fd_sc_hs__fa_2_5/a_336_347#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_27/a_817_508# fine_freq_track_1/sky130_fd_sc_hs__a211oi_4_1/a_92_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_33/a_910_118# fine_freq_track_1/sky130_fd_sc_hs__sdlclkp_1_1/a_288_48#
+ fine_freq_track_1/sky130_fd_sc_hs__a31oi_2_1/a_27_368# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_23/a_699_463#
+ fine_freq_track_1/sky130_fd_sc_hs__nor2_1_63/a_116_368# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_5/a_498_360#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_21/a_1550_119# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_11/a_37_78#
+ fine_freq_track_1/sky130_fd_sc_hs__a21oi_1_1/a_29_368# fine_freq_track_1/sky130_fd_sc_hs__a22o_1_25/a_132_392#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_1/a_706_463# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_27/a_1624_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_21/a_1598_93# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_25/a_812_138#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_65/a_812_138# fine_freq_track_1/sky130_fd_sc_hs__a21oi_1_37/a_117_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_43/a_856_304# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_71/a_1627_493#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_43/a_850_127# fine_freq_track_1/sky130_fd_sc_hs__o21ai_1_11/a_27_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_9/a_300_74# fine_freq_track_1/sky130_fd_sc_hs__a21oi_1_83/a_117_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_23/a_507_368# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_61/a_1350_392#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_35/a_789_463# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_55/a_313_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_29/a_498_360# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_83/a_1827_81#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_31/a_1547_508# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_41/a_796_463#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_73/a_789_463# fine_freq_track_1/sky130_fd_sc_hs__o21a_1_29/a_83_244#
+ fine_freq_track_1/sky130_fd_sc_hs__fa_2_19/a_487_79# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_9/a_910_118#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_21/a_313_74# fine_freq_track_1/sky130_fd_sc_hs__dfxtp_2_1/a_1172_124#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_25/a_706_463# fine_freq_track_1/sky130_fd_sc_hs__a222o_1_1/a_337_390#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_15/a_834_355# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_39/a_1627_493#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_55/a_834_355# fine_freq_track_1/sky130_fd_sc_hs__nor4_1_3/a_144_368#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_5/a_494_366# fine_freq_track_1/sky130_fd_sc_hs__o21a_1_73/a_83_244#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_91/a_2010_409# fine_freq_track_1/sky130_fd_sc_hs__maj3_1_3/a_223_120#
+ fine_freq_track_1/sky130_fd_sc_hs__nand2b_1_9/a_269_74# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_29/a_1350_392#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_35/a_1434_74# fine_freq_track_1/sky130_fd_sc_hs__a211oi_1_1/a_71_368#
+ fine_freq_track_1/sky130_fd_sc_hs__a22o_1_1/a_132_392# fine_freq_track_1/sky130_fd_sc_hs__dfxtp_2_5/a_1217_314#
+ fine_freq_track_1/sky130_fd_sc_hs__a22oi_1_15/a_339_74# fine_freq_track_1/sky130_fd_sc_hs__nand2_1_29/a_117_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_11/a_1482_48# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_43/a_2026_424#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_43/a_832_118# fine_freq_track_1/sky130_fd_sc_hs__nor2b_1_41/a_27_112#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_27/a_1465_471# fine_freq_track_1/sky130_fd_sc_hs__nand2_1_73/a_117_74#
+ fine_freq_track_1/sky130_fd_sc_hs__a21oi_1_117/a_117_74# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_17/a_817_508#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_59/a_2010_409# fine_freq_track_1/sky130_fd_sc_hs__nor3_1_7/a_114_368#
+ fine_freq_track_1/sky130_fd_sc_hs__dfxtp_4_2/a_735_102# fine_freq_track_1/sky130_fd_sc_hs__dfstp_2_1/a_225_74#
+ fine_freq_track_1/sky130_fd_sc_hs__nand2_4_13/a_27_74# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_13/a_699_463#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_33/a_124_78# fine_freq_track_1/sky130_fd_sc_hs__nor2_1_53/a_116_368#
+ fine_freq_track_1/sky130_fd_sc_hs__o211ai_1_3/a_311_74# fine_freq_track_1/sky130_fd_sc_hs__a21oi_1_89/a_29_368#
+ fine_freq_track_1/sky130_fd_sc_hs__dfxtp_4_3/a_1141_508# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_49/a_33_74#
+ fine_freq_track_1/sky130_fd_sc_hs__o21a_1_23/a_320_74# fine_freq_track_1/sky130_fd_sc_hs__a22o_1_15/a_132_392#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_91/a_699_463# fine_freq_track_1/sky130_fd_sc_hs__dfxtp_2_11/a_431_508#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_17/a_1624_74# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_39/a_1550_119#
+ fine_freq_track_1/sky130_fd_sc_hs__a22oi_1_7/a_71_368# fine_freq_track_1/sky130_fd_sc_hs__nor2b_1_29/a_278_368#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_11/a_1598_93# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_15/a_812_138#
+ fine_freq_track_1/sky130_fd_sc_hs__nand2_1_1/a_117_74# fine_freq_track_1/sky130_fd_sc_hs__a21oi_1_23/a_29_368#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_5/a_1736_119# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_55/a_812_138#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_33/a_856_304# fine_freq_track_1/sky130_fd_sc_hs__maj3_1_3/a_84_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_5/a_1266_119# fine_freq_track_1/sky130_fd_sc_hs__nor4_1_3/a_228_368#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_33/a_850_127# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_51/a_37_78#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_39/a_1647_81# fine_freq_track_1/sky130_fd_sc_hs__xor2_1_1/a_455_87#
+ fine_freq_track_1/sky130_fd_sc_hs__a21oi_1_5/a_29_368# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_89/a_1627_493#
+ fine_freq_track_1/sky130_fd_sc_hs__fa_2_1/a_1205_79# fine_freq_track
Xsky130_fd_sc_hs__einvp_8_11 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__inv_4_39/A sky130_fd_sc_hs__einvp_8_11/TE
+ osc_core_1/inj_out sky130_fd_sc_hs__einvp_8_11/a_802_323# sky130_fd_sc_hs__einvp_8_11/a_27_74#
+ sky130_fd_sc_hs__einvp_8_11/a_27_368# sky130_fd_sc_hs__einvp_8
Xsky130_fd_sc_hs__buf_2_16 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__buf_2_17/A sky130_fd_sc_hs__buf_2_17/X
+ sky130_fd_sc_hs__buf_2_17/a_21_260# sky130_fd_sc_hs__buf_2
Xsky130_fd_sc_hs__buf_2_27 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__buf_2_30/A sky130_fd_sc_hs__buf_2_30/X
+ sky130_fd_sc_hs__buf_2_30/a_21_260# sky130_fd_sc_hs__buf_2
Xsky130_fd_sc_hs__buf_2_38 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__buf_2_39/A sky130_fd_sc_hs__buf_2_39/X
+ sky130_fd_sc_hs__buf_2_39/a_21_260# sky130_fd_sc_hs__buf_2
Xsky130_fd_sc_hs__buf_2_49 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__buf_2_51/X sky130_fd_sc_hs__buf_2_49/X
+ sky130_fd_sc_hs__buf_2_49/a_21_260# sky130_fd_sc_hs__buf_2
Xsky130_fd_sc_hs__o21bai_2_18 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__buf_2_77/A
+ sky130_fd_sc_hs__nand2_2_33/Y sky130_fd_sc_hs__dlrtp_1_79/D sky130_fd_sc_hs__buf_2_79/A
+ sky130_fd_sc_hs__o21bai_2_19/a_27_74# sky130_fd_sc_hs__o21bai_2_19/a_225_74# sky130_fd_sc_hs__o21bai_2_19/a_507_368#
+ sky130_fd_sc_hs__o21bai_2
Xsky130_fd_sc_hs__o21bai_2_29 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__clkinv_4_5/Y
+ sky130_fd_sc_hs__buf_8_3/X sky130_fd_sc_hs__buf_2_103/X sky130_fd_sc_hs__buf_2_109/A
+ sky130_fd_sc_hs__o21bai_2_29/a_27_74# sky130_fd_sc_hs__o21bai_2_29/a_225_74# sky130_fd_sc_hs__o21bai_2_29/a_507_368#
+ sky130_fd_sc_hs__o21bai_2
Xsky130_fd_sc_hs__o21bai_4_7 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__buf_2_151/A
+ sky130_fd_sc_hs__o21bai_4_7/A1 sky130_fd_sc_hs__nand2_2_3/B sky130_fd_sc_hs__dlrtp_1_55/D
+ sky130_fd_sc_hs__o21bai_4_7/a_28_368# sky130_fd_sc_hs__o21bai_4_7/a_27_74# sky130_fd_sc_hs__o21bai_4_7/a_828_48#
+ sky130_fd_sc_hs__o21bai_4
Xsky130_fd_sc_hs__nand2_2_30 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__nand2_2_31/Y
+ sky130_fd_sc_hs__or4_2_1/C sky130_fd_sc_hs__or4_2_1/A sky130_fd_sc_hs__nand2_2_31/a_27_74#
+ sky130_fd_sc_hs__nand2_2
Xsky130_fd_sc_hs__conb_1_205 DVSS: DVDD: DVDD: DVSS: prbs_generator_syn_29/eqn[2]
+ prbs_generator_syn_29/eqn[1] sky130_fd_sc_hs__conb_1_205/a_165_290# sky130_fd_sc_hs__conb_1_205/a_21_290#
+ sky130_fd_sc_hs__conb_1
Xsky130_fd_sc_hs__conb_1_216 DVSS: DVDD: DVDD: DVSS: prbs_generator_syn_25/eqn[22]
+ prbs_generator_syn_25/eqn[20] sky130_fd_sc_hs__conb_1_217/a_165_290# sky130_fd_sc_hs__conb_1_217/a_21_290#
+ sky130_fd_sc_hs__conb_1
Xsky130_fd_sc_hs__conb_1_227 DVSS: DVDD: DVDD: DVSS: prbs_generator_syn_23/eqn[30]
+ sky130_fd_sc_hs__conb_1_227/HI sky130_fd_sc_hs__conb_1_227/a_165_290# sky130_fd_sc_hs__conb_1_227/a_21_290#
+ sky130_fd_sc_hs__conb_1
Xsky130_fd_sc_hs__conb_1_238 DVSS: DVDD: DVDD: DVSS: prbs_generator_syn_29/eqn[31]
+ prbs_generator_syn_29/cke sky130_fd_sc_hs__conb_1_239/a_165_290# sky130_fd_sc_hs__conb_1_239/a_21_290#
+ sky130_fd_sc_hs__conb_1
Xsky130_fd_sc_hs__conb_1_249 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__conb_1_249/LO
+ sky130_fd_sc_hs__conb_1_249/HI sky130_fd_sc_hs__conb_1_249/a_165_290# sky130_fd_sc_hs__conb_1_249/a_21_290#
+ sky130_fd_sc_hs__conb_1
Xsky130_fd_sc_hs__clkbuf_8_19 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__clkbuf_8_19/X
+ sky130_fd_sc_hs__clkbuf_8_19/A sky130_fd_sc_hs__clkbuf_8_19/a_125_368# sky130_fd_sc_hs__clkbuf_8
Xsky130_fd_sc_hs__diode_2_1 hr_16t4_mux_top_1/din[1] DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__diode_2
Xsky130_fd_sc_hs__o21bai_2_4 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__o21bai_2_5/A1
+ sky130_fd_sc_hs__nand2_2_3/B sky130_fd_sc_hs__dlrtp_1_55/D sky130_fd_sc_hs__buf_2_51/A
+ sky130_fd_sc_hs__o21bai_2_5/a_27_74# sky130_fd_sc_hs__o21bai_2_5/a_225_74# sky130_fd_sc_hs__o21bai_2_5/a_507_368#
+ sky130_fd_sc_hs__o21bai_2
Xsky130_fd_sc_hs__o21ai_2_20 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__inv_4_15/Y sky130_fd_sc_hs__or2b_4_5/X
+ sky130_fd_sc_hs__nand2_2_11/B sky130_fd_sc_hs__o21ai_2_21/Y sky130_fd_sc_hs__o21ai_2_21/a_116_368#
+ sky130_fd_sc_hs__o21ai_2_21/a_27_74# sky130_fd_sc_hs__o21ai_2
Xsky130_fd_sc_hs__o21ai_2_31 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__inv_4_19/Y sky130_fd_sc_hs__o21ai_2_31/A2
+ sky130_fd_sc_hs__o21ai_4_1/A1 sky130_fd_sc_hs__buf_2_83/A sky130_fd_sc_hs__o21ai_2_31/a_116_368#
+ sky130_fd_sc_hs__o21ai_2_31/a_27_74# sky130_fd_sc_hs__o21ai_2
Xsky130_fd_sc_hs__o21ai_2_42 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__inv_4_25/Y sky130_fd_sc_hs__or2b_2_3/A
+ sky130_fd_sc_hs__clkinv_4_7/Y sky130_fd_sc_hs__buf_2_129/A sky130_fd_sc_hs__o21ai_2_43/a_116_368#
+ sky130_fd_sc_hs__o21ai_2_43/a_27_74# sky130_fd_sc_hs__o21ai_2
Xsky130_fd_sc_hs__o21ai_2_53 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__nand2_2_27/B
+ sky130_fd_sc_hs__or2b_4_1/X sky130_fd_sc_hs__nand2_2_21/B sky130_fd_sc_hs__buf_2_137/A
+ sky130_fd_sc_hs__o21ai_2_53/a_116_368# sky130_fd_sc_hs__o21ai_2_53/a_27_74# sky130_fd_sc_hs__o21ai_2
Xsky130_fd_sc_hs__clkinv_4_12 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__o21bai_2_5/A1
+ sky130_fd_sc_hs__or4_2_1/C sky130_fd_sc_hs__clkinv_4
Xsky130_fd_sc_hs__einvn_1_1 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__inv_4_49/Y sky130_fd_sc_hs__buf_1_1/A
+ sky130_fd_sc_hs__clkinv_8_15/Y sky130_fd_sc_hs__einvn_1_1/a_281_100# sky130_fd_sc_hs__einvn_1_1/a_278_368#
+ sky130_fd_sc_hs__einvn_1_1/a_22_46# sky130_fd_sc_hs__einvn_1
Xprbs_generator_syn_14 prbs_generator_syn_19/clk prbs_generator_syn_19/rst prbs_generator_syn_15/cke
+ sky130_fd_sc_hs__conb_1_145/LO sky130_fd_sc_hs__conb_1_145/LO sky130_fd_sc_hs__conb_1_145/HI
+ sky130_fd_sc_hs__conb_1_145/HI sky130_fd_sc_hs__conb_1_145/HI sky130_fd_sc_hs__conb_1_145/HI
+ sky130_fd_sc_hs__conb_1_145/HI sky130_fd_sc_hs__conb_1_145/LO sky130_fd_sc_hs__conb_1_145/LO
+ sky130_fd_sc_hs__conb_1_145/LO sky130_fd_sc_hs__conb_1_145/LO prbs_generator_syn_15/eqn[31]
+ sky130_fd_sc_hs__conb_1_147/HI prbs_generator_syn_17/eqn[13] sky130_fd_sc_hs__conb_1_147/HI
+ prbs_generator_syn_17/eqn[13] sky130_fd_sc_hs__conb_1_147/HI prbs_generator_syn_17/eqn[13]
+ prbs_generator_syn_15/eqn[1] prbs_generator_syn_15/eqn[2] prbs_generator_syn_15/eqn[2]
+ prbs_generator_syn_15/eqn[2] prbs_generator_syn_15/eqn[2] prbs_generator_syn_15/eqn[1]
+ sky130_fd_sc_hs__conb_1_151/HI sky130_fd_sc_hs__conb_1_151/LO sky130_fd_sc_hs__conb_1_151/LO
+ sky130_fd_sc_hs__conb_1_151/HI sky130_fd_sc_hs__conb_1_151/LO sky130_fd_sc_hs__conb_1_151/HI
+ sky130_fd_sc_hs__conb_1_151/LO sky130_fd_sc_hs__conb_1_151/HI prbs_generator_syn_15/eqn[31]
+ prbs_generator_syn_15/eqn[30] prbs_generator_syn_15/eqn[30] prbs_generator_syn_15/eqn[30]
+ prbs_generator_syn_15/eqn[30] prbs_generator_syn_15/eqn[30] prbs_generator_syn_15/eqn[30]
+ prbs_generator_syn_15/eqn[30] prbs_generator_syn_15/eqn[30] prbs_generator_syn_15/eqn[22]
+ prbs_generator_syn_15/eqn[22] prbs_generator_syn_15/eqn[20] prbs_generator_syn_15/eqn[22]
+ prbs_generator_syn_15/eqn[22] prbs_generator_syn_15/eqn[22] prbs_generator_syn_15/eqn[22]
+ prbs_generator_syn_15/eqn[22] prbs_generator_syn_15/eqn[22] prbs_generator_syn_15/eqn[13]
+ prbs_generator_syn_15/eqn[13] prbs_generator_syn_15/eqn[13] prbs_generator_syn_15/eqn[9]
+ prbs_generator_syn_15/eqn[9] prbs_generator_syn_15/eqn[9] prbs_generator_syn_15/eqn[9]
+ prbs_generator_syn_15/eqn[9] prbs_generator_syn_15/eqn[9] prbs_generator_syn_15/eqn[9]
+ prbs_generator_syn_15/eqn[9] prbs_generator_syn_15/eqn[2] prbs_generator_syn_15/eqn[1]
+ prbs_generator_syn_15/eqn[2] prbs_generator_syn_19/inj_err prbs_generator_syn_15/eqn[31]
+ prbs_generator_syn_15/eqn[31] hr_16t4_mux_top_1/din[1] DVSS: DVDD: prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_1/a_293_74#
+ prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_15/X prbs_generator_syn_15/sky130_fd_sc_hs__nand2_1_35/B
+ prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_51/Y prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_9/A
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_9/CLK prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_47/a_27_74#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_37/a_1226_296# prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_3/B
+ prbs_generator_syn_15/sky130_fd_sc_hs__nor2b_1_7/a_27_112# prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_29/B
+ prbs_generator_syn_15/sky130_fd_sc_hs__sdlclkp_2_1/a_580_74# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_1/a_1141_508#
+ prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_5/Y prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_41/a_230_79#
+ prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_61/a_138_385# prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_43/a_132_392#
+ prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_3/a_222_392# prbs_generator_syn_15/sky130_fd_sc_hs__nor2b_1_9/a_27_112#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_61/a_27_74# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_35/a_206_368#
+ prbs_generator_syn_15/sky130_fd_sc_hs__nand2_2_3/Y prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_25/B
+ prbs_generator_syn_15/sky130_fd_sc_hs__nand2_1_11/a_117_74# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_67/a_651_503#
+ prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_45/X prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_39/a_696_458#
+ prbs_generator_syn_15/sky130_fd_sc_hs__sdlclkp_2_1/a_1198_74# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_45/a_1034_424#
+ prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_17/a_222_392# prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_55/a_222_392#
+ prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_53/Y prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_35/A
+ prbs_generator_syn_15/m3_13600_1651# prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_59/a_52_123#
+ prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_5/a_293_74# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_35/a_1226_296#
+ prbs_generator_syn_15/sky130_fd_sc_hs__nand2_1_51/B prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_5/a_651_503#
+ prbs_generator_syn_15/sky130_fd_sc_hs__nand2_1_21/B prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_8/a_27_74#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_15/a_27_74# prbs_generator_syn_15/sky130_fd_sc_hs__and2b_2_1/X
+ prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_13/X prbs_generator_syn_15/sky130_fd_sc_hs__nand2_2_3/a_27_74#
+ prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_50/a_138_385# prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_33/a_132_392#
+ prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_1/a_376_368# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_25/a_206_368#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_35/a_437_503# prbs_generator_syn_15/sky130_fd_sc_hs__sdlclkp_2_1/a_708_451#
+ prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_45/a_230_79# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_29/a_696_458#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_32/a_27_74# prbs_generator_syn_15/sky130_fd_sc_hs__nor2b_1_4/Y
+ prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_59/a_293_74# prbs_generator_syn_15/sky130_fd_sc_hs__nand2_1_47/a_117_74#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_73/a_735_102# prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_21/a_112_119#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_23/a_1141_508# prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_25/a_293_74#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_7/Q prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_3/a_112_119#
+ prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_35/B prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_51/X
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_53/a_1178_124# prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_23/a_132_392#
+ prbs_generator_syn_15/sky130_fd_sc_hs__nand2_1_3/B prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_15/a_206_368#
+ prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_63/a_132_392# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_55/a_27_74#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_25/a_437_503# prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_41/a_52_123#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_47/a_651_503# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_73/a_1141_508#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_19/a_696_458# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_57/a_696_458#
+ prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_7/X prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_43/a_1034_424#
+ prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_55/A prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_11/a_112_119#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_21/a_1141_508# prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_35/a_222_392#
+ prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_49/a_230_79# prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_67/Y
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_71/a_27_74# prbs_generator_syn_15/sky130_fd_sc_hs__nand2_1_33/B
+ prbs_generator_syn_15/sky130_fd_sc_hs__conb_1_1/LO prbs_generator_syn_15/sky130_fd_sc_hs__nand2_1_19/a_117_74#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_51/a_1178_124# prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_33/X
+ prbs_generator_syn_15/sky130_fd_sc_hs__nand2_1_29/B prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_41/Y
+ prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_53/a_132_392# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_45/a_206_368#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_15/a_437_503# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_37/a_651_503#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_39/a_544_485# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_53/a_735_102#
+ prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_45/a_52_123# prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_1/B
+ prbs_generator_syn_15/sky130_fd_sc_hs__nand2_2_3/B prbs_generator_syn_15/sky130_fd_sc_hs__clkbuf_16_1/A
+ prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_21/X prbs_generator_syn_15/sky130_fd_sc_hs__nand2_1_25/B
+ prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_39/a_376_368# prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_63/X
+ prbs_generator_syn_15/m3_13600_3481# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_69/a_1178_124#
+ prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_21/a_138_385# prbs_generator_syn_15/sky130_fd_sc_hs__nor2b_1_8/Y
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_19/a_1178_124# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_49/a_27_74#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_45/a_437_503# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_27/a_651_503#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_71/a_1141_508# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_65/a_651_503#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_29/a_544_485# prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_3/a_138_385#
+ prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_55/X prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_43/a_735_102#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_41/a_1034_424# prbs_generator_syn_15/sky130_fd_sc_hs__nand2_1_9/B
+ prbs_generator_syn_15/sky130_fd_sc_hs__nor2b_1_9/Y prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_59/a_1034_424#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_39/a_1141_508# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_33/a_1226_296#
+ prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_49/a_52_123# prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_47/Y
+ prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_43/Y prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_4/a_651_503#
+ prbs_generator_syn_15/sky130_fd_sc_hs__nand2_1_49/B prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_19/A
+ prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_11/a_138_385# prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_5/X
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_63/a_206_368# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_17/a_651_503#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_19/a_544_485# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_55/a_651_503#
+ prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_9/Y prbs_generator_syn_15/sky130_fd_sc_hs__nand2_1_17/B
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_57/a_544_485# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_67/a_696_458#
+ prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_35/X prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_19/a_27_74#
+ prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_45/a_222_392# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_32/a_1226_296#
+ prbs_generator_syn_15/sky130_fd_sc_hs__nand2_1_43/B prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_25/A
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_1/a_206_368# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_49/a_1226_296#
+ prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_1/a_112_119# prbs_generator_syn_15/sky130_fd_sc_hs__or2_1_1/X
+ prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_59/a_376_368# prbs_generator_syn_15/sky130_fd_sc_hs__nand2_1_19/B
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_5/a_696_458# prbs_generator_syn_15/sky130_fd_sc_hs__nor2b_1_1/Y
+ prbs_generator_syn_15/sky130_fd_sc_hs__nor2b_1_5/a_278_368# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_17/a_1178_124#
+ prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_39/X prbs_generator_syn_15/m3_13600_5433#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_63/a_437_503# prbs_generator_syn_15/sky130_fd_sc_hs__nand2_2_5/B
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_23/a_735_102# prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_53/A
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_61/a_735_102# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_57/a_1034_424#
+ prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_63/B prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_37/a_1141_508#
+ prbs_generator_syn_15/sky130_fd_sc_hs__nand2_1_47/B prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_29/X
+ prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_65/Y prbs_generator_syn_15/m3_13600_4701#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_1/a_437_503# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_67/a_1178_124#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_9/a_735_102# prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_13/a_132_392#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_15/a_1178_124# prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_15/A
+ prbs_generator_syn_15/sky130_fd_sc_hs__nand2_1_1/B prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_43/B
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_35/a_651_503# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_8/D
+ prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_29/A prbs_generator_syn_15/sky130_fd_sc_hs__nand2_1_7/B
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_13/a_735_102# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_47/a_696_458#
+ prbs_generator_syn_15/sky130_fd_sc_hs__nand2_1_31/B prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_51/a_735_102#
+ prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_59/X prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_35/a_1141_508#
+ prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_25/a_222_392# prbs_generator_syn_15/sky130_fd_sc_hs__sdlclkp_2_1/a_288_48#
+ prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_55/B prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_17/B
+ prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_43/A prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_7/A
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_65/a_1178_124# prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_59/Y
+ prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_41/X prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_21/a_230_79#
+ prbs_generator_syn_15/sky130_fd_sc_hs__nand2_1_57/a_117_74# prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_1/a_222_392#
+ prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_19/B prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_35/a_293_74#
+ prbs_generator_syn_15/sky130_fd_sc_hs__nand2_1_23/a_117_74# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_73/a_206_368#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_25/a_651_503# prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_1/a_138_385#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_37/a_696_458# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_67/a_544_485#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_43/a_27_74# prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_9/X
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_55/a_1034_424# prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_39/a_112_119#
+ prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_15/a_222_392# prbs_generator_syn_15/sky130_fd_sc_hs__conb_1_1/HI
+ prbs_generator_syn_15/sky130_fd_sc_hs__nand2_1_23/B prbs_generator_syn_15/sky130_fd_sc_hs__nand2_1_53/B
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_9/a_1178_124# prbs_generator_syn_15/sky130_fd_sc_hs__nor2b_1_4/A
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_47/a_1226_296# prbs_generator_syn_15/m3_13600_11045#
+ prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_17/X prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_29/a_376_368#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_5/a_544_485# prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_3/X
+ prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_31/a_132_392# prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_61/A
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_15/a_651_503# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_73/a_437_503#
+ prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_25/a_230_79# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_27/a_696_458#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_65/a_696_458# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_33/a_735_102#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_71/a_735_102# prbs_generator_syn_15/m3_13600_7263#
+ prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_43/a_222_392# prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_50/Y
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_8/a_1178_124# prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_53/B
+ prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_19/a_376_368# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_63/a_1178_124#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_4/a_696_458# prbs_generator_syn_15/sky130_fd_sc_hs__nor2b_1_4/a_278_368#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_13/a_1178_124# prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_61/a_132_392#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_53/a_206_368# prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_21/a_52_123#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_45/a_651_503# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_17/a_696_458#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_47/a_544_485# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_55/a_696_458#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_21/a_735_102# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_37/a_27_74#
+ prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_61/B prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_61/X
+ prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_59/a_112_119# prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_31/A
+ prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_33/a_222_392# prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_29/a_230_79#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_45/a_1226_296# prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_9/a_132_392#
+ prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_5/A prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_57/Y
+ prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_31/X prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_51/a_27_74#
+ prbs_generator_syn_15/sky130_fd_sc_hs__nor2b_1_8/a_27_112# prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_47/a_376_368#
+ prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_53/a_293_74# prbs_generator_syn_15/sky130_fd_sc_hs__nand2_1_43/a_117_74#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_8/a_735_102# prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_21/a_293_74#
+ prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_39/a_138_385# prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_63/Y
+ prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_51/a_132_392# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_43/a_206_368#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_53/a_437_503# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_37/a_544_485#
+ prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_57/X prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_53/a_1034_424#
+ prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_25/a_52_123# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_33/a_1141_508#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_63/Q prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_23/a_222_392#
+ prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_63/a_222_392# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_7/a_1178_124#
+ prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_53/X prbs_generator_syn_15/sky130_fd_sc_hs__nand2_2_5/Y
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_61/a_1178_124# prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_1/a_230_79#
+ prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_43/a_230_79# prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_11/a_230_79#
+ prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_41/a_132_392# prbs_generator_syn_15/sky130_fd_sc_hs__nand2_1_13/a_117_74#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_43/a_437_503# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_27/a_544_485#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_63/a_651_503# prbs_generator_syn_15/sky130_fd_sc_hs__nand2_1_7/a_117_74#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_35/a_696_458# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_65/a_544_485#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_51/a_1034_424# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_41/a_735_102#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_32/a_1141_508# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_49/a_1141_508#
+ prbs_generator_syn_15/sky130_fd_sc_hs__nand2_1_55/B prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_53/a_222_392#
+ prbs_generator_syn_15/sky130_fd_sc_hs__sdlclkp_2_1/a_114_112# prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_9/a_293_74#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_43/a_1226_296# prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_29/a_52_123#
+ prbs_generator_syn_15/sky130_fd_sc_hs__nand2_1_37/B prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_1/a_651_503#
+ prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_27/a_376_368# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_4/a_544_485#
+ prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_67/a_376_368# prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_27/X
+ prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_1/X prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_59/a_138_385#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_29/a_1178_124# prbs_generator_syn_15/m3_13600_2871#
+ prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_5/a_230_79# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_23/a_206_368#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_61/a_206_368# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_17/a_544_485#
+ prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_15/a_230_79# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_25/a_696_458#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_55/a_544_485# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_32/a_735_102#
+ prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_29/a_293_74# prbs_generator_syn_15/sky130_fd_sc_hs__nand2_1_17/a_117_74#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_69/a_1034_424# prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_29/a_112_119#
+ prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_37/X prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_31/B
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_19/a_1034_424# prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_33/A
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_9/a_206_368# prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_57/a_376_368#
+ prbs_generator_syn_15/sky130_fd_sc_hs__sdlclkp_2_1/a_706_317# prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_11/B
+ prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_1/a_52_123# prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_39/B
+ prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_21/a_132_392# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_13/a_206_368#
+ prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_43/a_52_123# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_51/a_206_368#
+ prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_47/X prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_23/a_437_503#
+ prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_11/a_52_123# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_61/a_437_503#
+ prbs_generator_syn_15/sky130_fd_sc_hs__nor2b_1_7/Y prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_51/A
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_15/a_696_458# prbs_generator_syn_15/sky130_fd_sc_hs__nor2b_1_5/Y
+ prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_9/a_230_79# prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_25/X
+ prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_19/a_112_119# prbs_generator_syn_15/sky130_fd_sc_hs__nand2_1_45/B
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_5/a_1178_124# prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_19/a_230_79#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_41/a_1226_296# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_59/a_1226_296#
+ prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_63/a_230_79# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_51/Q
+ prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_7/a_132_392# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_9/a_437_503#
+ prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_46/a_376_368# prbs_generator_syn_15/sky130_fd_sc_hs__nand2_1_33/a_117_74#
+ prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_11/a_293_74# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_27/a_1178_124#
+ prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_11/a_132_392# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_13/a_437_503#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_51/a_437_503# prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_5/a_52_123#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_35/a_544_485# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_73/a_651_503#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_45/a_696_458# prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_15/a_52_123#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_47/a_1141_508# prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_47/a_112_119#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_4/a_1178_124# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_17/a_1034_424#
+ prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_23/B prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_37/a_376_368#
+ prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_15/B prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_7/Y
+ prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_29/a_138_385# prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_33/a_230_79#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_25/a_1178_124# prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_47/a_293_74#
+ prbs_generator_syn_15/sky130_fd_sc_hs__nand2_1_37/a_117_74# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_33/a_206_368#
+ prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_15/a_293_74# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_71/a_206_368#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_25/a_544_485# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_67/a_1034_424#
+ prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_13/a_222_392# prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_9/a_52_123#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_15/a_1034_424# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_57/a_1226_296#
+ prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_19/a_52_123# prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_23/X
+ prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_63/a_52_123# prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_19/a_138_385#
+ prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_9/a_376_368# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_21/a_206_368#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_33/a_437_503# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_71/a_437_503#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_53/a_651_503# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_15/a_544_485#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_63/a_696_458# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_65/a_1034_424#
+ prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_19/a_293_74# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_45/a_1141_508#
+ prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_27/a_112_119# prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_67/a_112_119#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_1/a_1178_124# prbs_generator_syn_15/sky130_fd_sc_hs__conb_1_1/a_21_290#
+ prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_63/a_293_74# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_8/a_206_368#
+ prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_17/a_376_368# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_63/a_27_74#
+ prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_21/A prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_55/a_376_368#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_1/a_696_458# prbs_generator_syn_15/sky130_fd_sc_hs__nor2b_1_1/a_278_368#
+ prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_47/a_138_385# prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_33/a_52_123#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_9/a_1034_424# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_21/a_437_503#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_1/a_27_74# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_43/a_651_503#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_1/Q prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_45/a_544_485#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_69/a_735_102# prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_57/a_112_119#
+ prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_31/a_222_392# prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_13/A
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_55/a_1226_296# prbs_generator_syn_15/sky130_fd_sc_hs__nand2_2_5/a_27_74#
+ prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_53/a_230_79# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_8/a_437_503#
+ prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_67/a_293_74# prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_33/a_293_74#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_7/a_735_102# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_23/a_1178_124#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_41/a_206_368# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_8/a_1034_424#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_63/a_1034_424# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_59/a_735_102#
+ prbs_generator_syn_15/sky130_fd_sc_hs__nand2_1_5/B prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_43/a_1141_508#
+ prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_46/a_112_119# prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_61/a_222_392#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_13/a_1034_424# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_73/a_1178_124#
+ prbs_generator_syn_15/sky130_fd_sc_hs__nand2_1_27/B prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_13/B
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_57/a_27_74# prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_57/a_230_79#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_21/a_1178_124# prbs_generator_syn_15/sky130_fd_sc_hs__nor2b_1_1/a_27_112#
+ prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_27/a_138_385# prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_23/a_230_79#
+ prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_67/a_138_385# prbs_generator_syn_15/sky130_fd_sc_hs__nand2_1_41/B
+ prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_9/a_222_392# prbs_generator_syn_15/sky130_fd_sc_hs__nand2_1_27/a_117_74#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_32/a_206_368# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_23/a_651_503#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_41/a_437_503# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_73/a_27_74#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_61/a_651_503# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_63/a_544_485#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_49/a_735_102# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_73/a_696_458#
+ prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_37/a_112_119# prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_51/a_222_392#
+ prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_43/X prbs_generator_syn_15/sky130_fd_sc_hs__nand2_2_1/B
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_9/a_651_503# prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_53/a_52_123#
+ prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_49/X prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_25/a_376_368#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_1/a_544_485# prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_65/a_376_368#
+ prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_57/a_138_385# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_27/a_27_74#
+ prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_39/a_132_392# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_7/a_1034_424#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_13/a_651_503# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_32/a_437_503#
+ prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_27/a_230_79# prbs_generator_syn_15/m3_13600_12265#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_51/a_651_503# prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_59/B
+ prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_47/A prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_61/a_1034_424#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_41/a_1141_508# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_59/a_1141_508#
+ prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_41/a_222_392# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_53/a_1226_296#
+ prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_3/A prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_71/a_1178_124#
+ prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_9/a_112_119# prbs_generator_syn_15/sky130_fd_sc_hs__nand2_1_3/a_117_74#
+ prbs_generator_syn_15/m3_13600_8483# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_39/a_1178_124#
+ prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_57/a_52_123# prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_46/a_138_385#
+ prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_23/a_52_123# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_67/a_27_74#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_53/a_696_458# prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_17/a_112_119#
+ prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_11/A prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_55/a_112_119#
+ prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_1/A prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_51/a_1226_296#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_29/a_1034_424# prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_59/A
+ prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_23/A prbs_generator_syn_15/sky130_fd_sc_hs__nand2_1_39/B
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_5/a_27_74# prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_57/a_293_74#
+ prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_37/a_138_385# prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_59/a_132_392#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_33/a_651_503# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_71/a_651_503#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_43/a_696_458# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_73/a_544_485#
+ prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_27/a_52_123# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_57/a_1141_508#
+ prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_21/a_222_392# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_35/a_27_74#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_69/a_1226_296# prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_37/B
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_19/a_1226_296# prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_35/a_376_368#
+ prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_47/a_230_79# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_37/a_1178_124#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_5/a_1034_424# prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_49/a_132_392#
+ prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_7/a_222_392# prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_27/a_293_74#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_21/a_651_503# prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_9/a_138_385#
+ prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_11/a_222_392# prbs_generator_syn_15/m3_13600_14095#
+ prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_50/A prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_27/a_1034_424#
+ prbs_generator_syn_15/sky130_fd_sc_hs__nand2_1_13/B prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_8/a_651_503#
+ prbs_generator_syn_15/m3_13600_9703# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_35/a_1178_124#
+ prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_17/a_138_385# prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_55/a_138_385#
+ prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_7/a_230_79# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_4/a_1034_424#
+ prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_7/a_376_368# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_69/a_206_368#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_23/a_696_458# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_53/a_544_485#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_39/a_735_102# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_61/a_696_458#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_55/a_1141_508# prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_25/a_112_119#
+ prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_65/a_112_119# prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_43/a_293_74#
+ prbs_generator_syn_15/sky130_fd_sc_hs__nand2_1_57/B prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_25/a_1034_424#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_7/a_206_368# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_17/a_1226_296#
+ prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_15/a_376_368# prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_53/a_376_368#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_9/a_696_458# prbs_generator_syn_15/m3_13600_431#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_45/a_27_74# prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_47/a_52_123#
+ prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_29/a_132_392# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_59/a_206_368#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_69/a_437_503# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_41/a_651_503#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_43/a_544_485# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_13/a_696_458#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_29/a_735_102# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_51/a_696_458#
+ prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_61/Y prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_67/a_1226_296#
+ prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_5/a_132_392# prbs_generator_syn_15/sky130_fd_sc_hs__and2b_2_1/a_198_48#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_7/a_437_503# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_15/a_1226_296#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_69/a_27_74# prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_46/a_293_74#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_1/a_1034_424# prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_19/a_132_392#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_49/a_206_368# prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_7/a_52_123#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_59/a_437_503# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_32/a_651_503#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_7/a_27_74# prbs_generator_syn_15/sky130_fd_sc_hs__nand2_2_1/a_27_74#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_19/a_735_102# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_57/a_735_102#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_65/a_1226_296# prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_37/A
+ prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_33/a_376_368# prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_37/a_230_79#
+ prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_25/a_138_385# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_39/a_27_74#
+ prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_65/a_138_385# prbs_generator_syn_15/sky130_fd_sc_hs__nor2b_1_9/a_278_368#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_49/a_437_503# prbs_generator_syn_15/sky130_fd_sc_hs__and2b_2_1/a_505_74#
+ prbs_generator_syn_15/sky130_fd_sc_hs__nand2_1_51/a_117_74# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_23/a_544_485#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_33/a_696_458# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_61/a_544_485#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_9/a_1226_296# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_53/a_1141_508#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_71/a_696_458# prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_35/a_112_119#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_23/a_1034_424# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_9/a_544_485#
+ prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_63/a_376_368# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_33/a_1178_124#
+ prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_5/a_376_368# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_13/a_544_485#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_73/a_1034_424# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_21/a_696_458#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_51/a_544_485# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_8/a_1226_296#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_51/a_1141_508# prbs_generator_syn_15/sky130_fd_sc_hs__nand2_1_55/a_117_74#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_21/a_1034_424# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_63/a_1226_296#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_23/a_27_74# prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_7/a_112_119#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_13/a_1226_296# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_8/a_696_458#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_32/a_1178_124# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_49/a_1178_124#
+ prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_37/a_52_123# prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_27/a_132_392#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_71/Q prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_67/a_735_102#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_69/a_1141_508# prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_15/a_112_119#
+ prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_53/a_112_119# prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_39/a_222_392#
+ prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_55/a_230_79# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_19/a_1141_508#
+ prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_37/a_293_74# prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_43/a_376_368#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_5/a_735_102# prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_35/a_138_385#
+ prbs_generator_syn_15/sky130_fd_sc_hs__sdlclkp_2_1/a_114_424# prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_57/a_132_392#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_71/a_1034_424# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_7/a_1226_296#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_33/a_544_485# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_41/a_696_458#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_71/a_544_485# prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_21/B
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_61/a_1226_296# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_39/a_1034_424#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_17/a_27_74# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_9/a_27_74#
+ prbs_generator_syn_15/sky130_fd_sc_hs__nor2b_1_5/a_27_112# prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_47/a_132_392#
+ prbs_generator_syn_15/sky130_fd_sc_hs__nor2b_1_8/a_278_368# prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_9/B
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_39/a_206_368# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_33/a_27_74#
+ prbs_generator_syn_15/sky130_fd_sc_hs__nand2_1_41/a_117_74# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_69/a_651_503#
+ prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_51/a_293_74# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_21/a_544_485#
+ prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_7/a_138_385# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_32/a_696_458#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_47/a_735_102# prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_33/a_112_119#
+ prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_59/a_222_392# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_17/a_1141_508#
+ prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_55/a_52_123# prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_3/a_293_74#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_7/a_651_503# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_29/a_1226_296#
+ prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_23/a_376_368# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_8/a_544_485#
+ prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_47/B prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_47/a_1178_124#
+ prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_15/a_138_385# prbs_generator_syn_15/sky130_fd_sc_hs__sdlclkp_2_1/a_1195_374#
+ prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_53/a_138_385# prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_37/a_132_392#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_29/a_206_368# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_39/a_437_503#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_59/a_651_503# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_37/a_735_102#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_67/a_1141_508# prbs_generator_syn_15/sky130_fd_sc_hs__and2b_2_1/a_27_74#
+ prbs_generator_syn_15/sky130_fd_sc_hs__conb_1_1/a_165_290# prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_55/a_293_74#
+ prbs_generator_syn_15/sky130_fd_sc_hs__nand2_1_45/a_117_74# prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_63/a_112_119#
+ prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_49/a_222_392# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_37/a_1034_424#
+ prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_23/a_293_74# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_15/a_1141_508#
+ prbs_generator_syn_15/sky130_fd_sc_hs__nand2_1_5/a_117_74# prbs_generator_syn_15/m3_13600_13485#
+ prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_5/a_112_119# prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_13/a_376_368#
+ prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_51/a_376_368# prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_7/a_293_74#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_19/a_206_368# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_57/a_206_368#
+ prbs_generator_syn_15/sky130_fd_sc_hs__sdlclkp_2_1/a_318_74# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_29/a_437_503#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_49/a_651_503# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_25/a_27_74#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_5/a_1226_296# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_41/a_544_485#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_27/a_735_102# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_65/a_1141_508#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_65/a_735_102# prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_3/a_230_79#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_35/a_1034_424# prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_13/a_230_79#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_41/a_27_74# prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_3/a_132_392#
+ prbs_generator_syn_15/sky130_fd_sc_hs__nand2_1_49/a_117_74# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_27/a_1226_296#
+ prbs_generator_syn_15/sky130_fd_sc_hs__nand2_1_15/a_117_74# prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_41/a_376_368#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_45/a_1178_124# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_4/a_735_102#
+ prbs_generator_syn_15/sky130_fd_sc_hs__nand2_1_9/a_117_74# prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_33/a_138_385#
+ prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_17/a_132_392# prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_55/a_132_392#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_9/a_1141_508# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_19/a_437_503#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_57/a_437_503# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_4/a_1226_296#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_32/a_544_485# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_17/a_735_102#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_55/a_735_102# prbs_generator_syn_15/m3_13600_2261#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_65/a_27_74# prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_29/a_222_392#
+ prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_43/a_112_119# prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_19/X
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_25/a_1226_296# prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_31/a_376_368#
+ prbs_generator_syn_15/sky130_fd_sc_hs__or2_1_1/a_63_368# prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_17/a_230_79#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_4/a_27_74# prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_61/a_230_79#
+ prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_63/a_138_385# prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_5/a_222_392#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_8/a_1141_508# prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_41/a_293_74#
+ prbs_generator_syn_15/sky130_fd_sc_hs__nand2_1_31/a_117_74# prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_5/a_138_385#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_63/a_1141_508# prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_19/a_222_392#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_13/a_1141_508# prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_3/a_52_123#
+ prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_13/a_52_123# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_43/a_1178_124#
+ prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_61/a_376_368# prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_35/a_132_392#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_67/a_206_368# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_1/a_1226_296#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_69/a_696_458# prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_31/a_230_79#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_35/a_735_102# prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_23/a_112_119#
+ prbs_generator_syn_15/sky130_fd_sc_hs__nand2_1_35/a_117_74# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_59/a_27_74#
+ prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_13/a_293_74# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_5/a_206_368#
+ prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_50/a_376_368# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_7/a_696_458#
+ prbs_generator_syn_15/sky130_fd_sc_hs__nor2b_1_7/a_278_368# prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_17/a_52_123#
+ prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_43/a_138_385# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_7/a_1141_508#
+ prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_61/a_52_123# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_67/a_437_503#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_61/a_1141_508# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_25/a_735_102#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_59/a_696_458# prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_13/a_112_119#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_33/a_1034_424# prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_51/a_112_119#
+ prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_35/a_230_79# prbs_generator_syn_15/m3_13600_4091#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_23/a_1226_296# prbs_generator_syn_15/sky130_fd_sc_hs__nand2_1_39/a_117_74#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_29/a_27_74# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_5/a_437_503#
+ prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_17/a_293_74# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_41/a_1178_124#
+ prbs_generator_syn_15/sky130_fd_sc_hs__or2_1_1/a_152_368# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_59/a_1178_124#
+ prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_61/a_293_74# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_47/a_206_368#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_39/a_651_503# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_49/a_696_458#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_15/a_735_102# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_32/a_1034_424#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_73/a_1226_296# prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_27/a_222_392#
+ prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_41/a_112_119# prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_31/a_52_123#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_49/a_1034_424# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_29/a_1141_508#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_21/a_1226_296# prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_39/a_230_79#
+ prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_23/a_138_385# prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_51/a_230_79#
+ prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_45/a_132_392# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_37/a_206_368#
+ prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_65/a_293_74# prbs_generator_syn_15/sky130_fd_sc_hs__nand2_1_53/a_117_74#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_47/a_437_503# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_29/a_651_503#
+ prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_31/a_293_74# prbs_generator_syn_15/sky130_fd_sc_hs__nand2_1_21/a_117_74#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_69/a_544_485# prbs_generator_syn_15/sky130_fd_sc_hs__clkbuf_16_1/a_114_74#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_45/a_735_102# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_13/a_27_74#
+ prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_31/a_112_119# prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_57/a_222_392#
+ prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_35/a_52_123# prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_21/a_376_368#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_7/a_544_485# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_57/a_1178_124#
+ prbs_generator_syn_15/m3_13600_6043# prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_13/a_138_385#
+ prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_51/a_138_385# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_5/a_1141_508#
+ prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_3/a_376_368# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_27/a_206_368#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_65/a_206_368# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_37/a_437_503#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_19/a_651_503# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_57/a_651_503#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_59/a_544_485# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_71/a_1226_296#
+ prbs_generator_syn_15/sky130_fd_sc_hs__nand2_1_25/a_117_74# prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_61/a_112_119#
+ prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_47/a_222_392# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_27/a_1141_508#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_53/a_27_74# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_4/a_206_368#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_39/a_1226_296# prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_11/a_376_368#
+ prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_39/a_52_123# prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_41/a_138_385#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_4/a_1141_508# prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_25/a_132_392#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_17/a_206_368# prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_41/A
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_55/a_206_368# prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_51/a_52_123#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_27/a_437_503# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_65/a_437_503#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_49/a_544_485# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_63/a_735_102#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_47/a_1034_424# prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_50/a_112_119#
+ prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_37/a_222_392# prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_59/a_230_79#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_25/a_1141_508# prbs_generator_syn_15/sky130_fd_sc_hs__nor2b_1_4/a_27_112#
+ prbs_generator_syn_15/sky130_fd_sc_hs__sdlclkp_2_1/a_685_81# prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_1/a_132_392#
+ prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_39/a_293_74# prbs_generator_syn_15/sky130_fd_sc_hs__nand2_1_29/a_117_74#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_4/a_437_503# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_55/a_1178_124#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_21/a_27_74# prbs_generator_syn_15/m3_13600_12875#
+ prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_50/a_293_74# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_1/a_735_102#
+ prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_31/a_138_385# prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_15/a_132_392#
+ prbs_generator_syn_15/sky130_fd_sc_hs__nand2_1_1/a_117_74# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_17/a_437_503#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_55/a_437_503# prbs_generator_syn
Xprbs_generator_syn_25 prbs_generator_syn_31/clk prbs_generator_syn_27/rst prbs_generator_syn_25/cke
+ sky130_fd_sc_hs__conb_1_249/LO sky130_fd_sc_hs__conb_1_249/HI sky130_fd_sc_hs__conb_1_249/HI
+ sky130_fd_sc_hs__conb_1_249/HI sky130_fd_sc_hs__conb_1_249/HI sky130_fd_sc_hs__conb_1_249/HI
+ sky130_fd_sc_hs__conb_1_249/HI sky130_fd_sc_hs__conb_1_249/HI sky130_fd_sc_hs__conb_1_249/HI
+ sky130_fd_sc_hs__conb_1_249/LO sky130_fd_sc_hs__conb_1_249/LO prbs_generator_syn_25/eqn[31]
+ prbs_generator_syn_25/cke prbs_generator_syn_25/eqn[31] prbs_generator_syn_25/cke
+ prbs_generator_syn_25/eqn[31] prbs_generator_syn_25/cke prbs_generator_syn_25/cke
+ sky130_fd_sc_hs__conb_1_233/HI prbs_generator_syn_27/eqn[20] prbs_generator_syn_27/eqn[20]
+ prbs_generator_syn_27/eqn[20] prbs_generator_syn_27/eqn[22] prbs_generator_syn_27/eqn[28]
+ sky130_fd_sc_hs__conb_1_251/HI sky130_fd_sc_hs__conb_1_251/HI prbs_generator_syn_27/eqn[28]
+ prbs_generator_syn_27/eqn[30] sky130_fd_sc_hs__conb_1_253/HI sky130_fd_sc_hs__conb_1_253/HI
+ sky130_fd_sc_hs__conb_1_253/HI sky130_fd_sc_hs__conb_1_253/HI prbs_generator_syn_25/eqn[31]
+ prbs_generator_syn_25/eqn[30] prbs_generator_syn_25/eqn[30] prbs_generator_syn_25/eqn[30]
+ prbs_generator_syn_25/eqn[30] prbs_generator_syn_25/eqn[30] prbs_generator_syn_25/eqn[30]
+ prbs_generator_syn_25/eqn[30] prbs_generator_syn_25/eqn[30] prbs_generator_syn_25/eqn[22]
+ prbs_generator_syn_25/eqn[22] prbs_generator_syn_25/eqn[20] prbs_generator_syn_25/eqn[22]
+ prbs_generator_syn_25/eqn[22] prbs_generator_syn_25/eqn[22] prbs_generator_syn_25/eqn[22]
+ prbs_generator_syn_25/eqn[22] prbs_generator_syn_25/eqn[22] prbs_generator_syn_25/eqn[9]
+ prbs_generator_syn_25/eqn[9] prbs_generator_syn_25/eqn[9] prbs_generator_syn_25/eqn[9]
+ prbs_generator_syn_25/eqn[9] prbs_generator_syn_25/eqn[8] prbs_generator_syn_25/eqn[8]
+ prbs_generator_syn_25/eqn[8] prbs_generator_syn_25/eqn[8] prbs_generator_syn_25/eqn[8]
+ prbs_generator_syn_25/eqn[8] prbs_generator_syn_25/eqn[8] prbs_generator_syn_25/eqn[1]
+ prbs_generator_syn_27/eqn[9] prbs_generator_syn_27/inj_err prbs_generator_syn_25/eqn[31]
+ prbs_generator_syn_25/eqn[31] hr_16t4_mux_top_1/din[0] DVSS: DVDD: prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_1/a_293_74#
+ prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_15/X prbs_generator_syn_25/sky130_fd_sc_hs__nand2_1_35/B
+ prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_51/Y prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_9/A
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_9/CLK prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_47/a_27_74#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_37/a_1226_296# prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_3/B
+ prbs_generator_syn_25/sky130_fd_sc_hs__nor2b_1_7/a_27_112# prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_29/B
+ prbs_generator_syn_25/sky130_fd_sc_hs__sdlclkp_2_1/a_580_74# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_1/a_1141_508#
+ prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_5/Y prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_41/a_230_79#
+ prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_61/a_138_385# prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_43/a_132_392#
+ prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_3/a_222_392# prbs_generator_syn_25/sky130_fd_sc_hs__nor2b_1_9/a_27_112#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_61/a_27_74# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_35/a_206_368#
+ prbs_generator_syn_25/sky130_fd_sc_hs__nand2_2_3/Y prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_25/B
+ prbs_generator_syn_25/sky130_fd_sc_hs__nand2_1_11/a_117_74# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_67/a_651_503#
+ prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_45/X prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_39/a_696_458#
+ prbs_generator_syn_25/sky130_fd_sc_hs__sdlclkp_2_1/a_1198_74# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_45/a_1034_424#
+ prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_17/a_222_392# prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_55/a_222_392#
+ prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_53/Y prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_35/A
+ prbs_generator_syn_25/m3_13600_1651# prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_59/a_52_123#
+ prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_5/a_293_74# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_35/a_1226_296#
+ prbs_generator_syn_25/sky130_fd_sc_hs__nand2_1_51/B prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_5/a_651_503#
+ prbs_generator_syn_25/sky130_fd_sc_hs__nand2_1_21/B prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_8/a_27_74#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_15/a_27_74# prbs_generator_syn_25/sky130_fd_sc_hs__and2b_2_1/X
+ prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_13/X prbs_generator_syn_25/sky130_fd_sc_hs__nand2_2_3/a_27_74#
+ prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_50/a_138_385# prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_33/a_132_392#
+ prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_1/a_376_368# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_25/a_206_368#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_35/a_437_503# prbs_generator_syn_25/sky130_fd_sc_hs__sdlclkp_2_1/a_708_451#
+ prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_45/a_230_79# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_29/a_696_458#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_32/a_27_74# prbs_generator_syn_25/sky130_fd_sc_hs__nor2b_1_4/Y
+ prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_59/a_293_74# prbs_generator_syn_25/sky130_fd_sc_hs__nand2_1_47/a_117_74#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_73/a_735_102# prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_21/a_112_119#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_23/a_1141_508# prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_25/a_293_74#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_7/Q prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_3/a_112_119#
+ prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_35/B prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_51/X
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_53/a_1178_124# prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_23/a_132_392#
+ prbs_generator_syn_25/sky130_fd_sc_hs__nand2_1_3/B prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_15/a_206_368#
+ prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_63/a_132_392# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_55/a_27_74#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_25/a_437_503# prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_41/a_52_123#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_47/a_651_503# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_73/a_1141_508#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_19/a_696_458# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_57/a_696_458#
+ prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_7/X prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_43/a_1034_424#
+ prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_55/A prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_11/a_112_119#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_21/a_1141_508# prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_35/a_222_392#
+ prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_49/a_230_79# prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_67/Y
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_71/a_27_74# prbs_generator_syn_25/sky130_fd_sc_hs__nand2_1_33/B
+ prbs_generator_syn_25/sky130_fd_sc_hs__conb_1_1/LO prbs_generator_syn_25/sky130_fd_sc_hs__nand2_1_19/a_117_74#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_51/a_1178_124# prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_33/X
+ prbs_generator_syn_25/sky130_fd_sc_hs__nand2_1_29/B prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_41/Y
+ prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_53/a_132_392# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_45/a_206_368#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_15/a_437_503# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_37/a_651_503#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_39/a_544_485# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_53/a_735_102#
+ prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_45/a_52_123# prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_1/B
+ prbs_generator_syn_25/sky130_fd_sc_hs__nand2_2_3/B prbs_generator_syn_25/sky130_fd_sc_hs__clkbuf_16_1/A
+ prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_21/X prbs_generator_syn_25/sky130_fd_sc_hs__nand2_1_25/B
+ prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_39/a_376_368# prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_63/X
+ prbs_generator_syn_25/m3_13600_3481# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_69/a_1178_124#
+ prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_21/a_138_385# prbs_generator_syn_25/sky130_fd_sc_hs__nor2b_1_8/Y
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_19/a_1178_124# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_49/a_27_74#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_45/a_437_503# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_27/a_651_503#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_71/a_1141_508# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_65/a_651_503#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_29/a_544_485# prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_3/a_138_385#
+ prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_55/X prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_43/a_735_102#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_41/a_1034_424# prbs_generator_syn_25/sky130_fd_sc_hs__nand2_1_9/B
+ prbs_generator_syn_25/sky130_fd_sc_hs__nor2b_1_9/Y prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_59/a_1034_424#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_39/a_1141_508# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_33/a_1226_296#
+ prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_49/a_52_123# prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_47/Y
+ prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_43/Y prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_4/a_651_503#
+ prbs_generator_syn_25/sky130_fd_sc_hs__nand2_1_49/B prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_19/A
+ prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_11/a_138_385# prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_5/X
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_63/a_206_368# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_17/a_651_503#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_19/a_544_485# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_55/a_651_503#
+ prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_9/Y prbs_generator_syn_25/sky130_fd_sc_hs__nand2_1_17/B
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_57/a_544_485# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_67/a_696_458#
+ prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_35/X prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_19/a_27_74#
+ prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_45/a_222_392# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_32/a_1226_296#
+ prbs_generator_syn_25/sky130_fd_sc_hs__nand2_1_43/B prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_25/A
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_1/a_206_368# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_49/a_1226_296#
+ prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_1/a_112_119# prbs_generator_syn_25/sky130_fd_sc_hs__or2_1_1/X
+ prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_59/a_376_368# prbs_generator_syn_25/sky130_fd_sc_hs__nand2_1_19/B
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_5/a_696_458# prbs_generator_syn_25/sky130_fd_sc_hs__nor2b_1_1/Y
+ prbs_generator_syn_25/sky130_fd_sc_hs__nor2b_1_5/a_278_368# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_17/a_1178_124#
+ prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_39/X prbs_generator_syn_25/m3_13600_5433#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_63/a_437_503# prbs_generator_syn_25/sky130_fd_sc_hs__nand2_2_5/B
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_23/a_735_102# prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_53/A
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_61/a_735_102# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_57/a_1034_424#
+ prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_63/B prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_37/a_1141_508#
+ prbs_generator_syn_25/sky130_fd_sc_hs__nand2_1_47/B prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_29/X
+ prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_65/Y prbs_generator_syn_25/m3_13600_4701#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_1/a_437_503# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_67/a_1178_124#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_9/a_735_102# prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_13/a_132_392#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_15/a_1178_124# prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_15/A
+ prbs_generator_syn_25/sky130_fd_sc_hs__nand2_1_1/B prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_43/B
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_35/a_651_503# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_8/D
+ prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_29/A prbs_generator_syn_25/sky130_fd_sc_hs__nand2_1_7/B
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_13/a_735_102# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_47/a_696_458#
+ prbs_generator_syn_25/sky130_fd_sc_hs__nand2_1_31/B prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_51/a_735_102#
+ prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_59/X prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_35/a_1141_508#
+ prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_25/a_222_392# prbs_generator_syn_25/sky130_fd_sc_hs__sdlclkp_2_1/a_288_48#
+ prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_55/B prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_17/B
+ prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_43/A prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_7/A
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_65/a_1178_124# prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_59/Y
+ prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_41/X prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_21/a_230_79#
+ prbs_generator_syn_25/sky130_fd_sc_hs__nand2_1_57/a_117_74# prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_1/a_222_392#
+ prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_19/B prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_35/a_293_74#
+ prbs_generator_syn_25/sky130_fd_sc_hs__nand2_1_23/a_117_74# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_73/a_206_368#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_25/a_651_503# prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_1/a_138_385#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_37/a_696_458# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_67/a_544_485#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_43/a_27_74# prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_9/X
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_55/a_1034_424# prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_39/a_112_119#
+ prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_15/a_222_392# prbs_generator_syn_25/sky130_fd_sc_hs__conb_1_1/HI
+ prbs_generator_syn_25/sky130_fd_sc_hs__nand2_1_23/B prbs_generator_syn_25/sky130_fd_sc_hs__nand2_1_53/B
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_9/a_1178_124# prbs_generator_syn_25/sky130_fd_sc_hs__nor2b_1_4/A
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_47/a_1226_296# prbs_generator_syn_25/m3_13600_11045#
+ prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_17/X prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_29/a_376_368#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_5/a_544_485# prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_3/X
+ prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_31/a_132_392# prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_61/A
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_15/a_651_503# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_73/a_437_503#
+ prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_25/a_230_79# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_27/a_696_458#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_65/a_696_458# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_33/a_735_102#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_71/a_735_102# prbs_generator_syn_25/m3_13600_7263#
+ prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_43/a_222_392# prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_50/Y
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_8/a_1178_124# prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_53/B
+ prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_19/a_376_368# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_63/a_1178_124#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_4/a_696_458# prbs_generator_syn_25/sky130_fd_sc_hs__nor2b_1_4/a_278_368#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_13/a_1178_124# prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_61/a_132_392#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_53/a_206_368# prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_21/a_52_123#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_45/a_651_503# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_17/a_696_458#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_47/a_544_485# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_55/a_696_458#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_21/a_735_102# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_37/a_27_74#
+ prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_61/B prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_61/X
+ prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_59/a_112_119# prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_31/A
+ prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_33/a_222_392# prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_29/a_230_79#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_45/a_1226_296# prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_9/a_132_392#
+ prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_5/A prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_57/Y
+ prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_31/X prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_51/a_27_74#
+ prbs_generator_syn_25/sky130_fd_sc_hs__nor2b_1_8/a_27_112# prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_47/a_376_368#
+ prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_53/a_293_74# prbs_generator_syn_25/sky130_fd_sc_hs__nand2_1_43/a_117_74#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_8/a_735_102# prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_21/a_293_74#
+ prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_39/a_138_385# prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_63/Y
+ prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_51/a_132_392# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_43/a_206_368#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_53/a_437_503# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_37/a_544_485#
+ prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_57/X prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_53/a_1034_424#
+ prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_25/a_52_123# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_33/a_1141_508#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_63/Q prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_23/a_222_392#
+ prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_63/a_222_392# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_7/a_1178_124#
+ prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_53/X prbs_generator_syn_25/sky130_fd_sc_hs__nand2_2_5/Y
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_61/a_1178_124# prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_1/a_230_79#
+ prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_43/a_230_79# prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_11/a_230_79#
+ prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_41/a_132_392# prbs_generator_syn_25/sky130_fd_sc_hs__nand2_1_13/a_117_74#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_43/a_437_503# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_27/a_544_485#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_63/a_651_503# prbs_generator_syn_25/sky130_fd_sc_hs__nand2_1_7/a_117_74#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_35/a_696_458# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_65/a_544_485#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_51/a_1034_424# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_41/a_735_102#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_32/a_1141_508# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_49/a_1141_508#
+ prbs_generator_syn_25/sky130_fd_sc_hs__nand2_1_55/B prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_53/a_222_392#
+ prbs_generator_syn_25/sky130_fd_sc_hs__sdlclkp_2_1/a_114_112# prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_9/a_293_74#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_43/a_1226_296# prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_29/a_52_123#
+ prbs_generator_syn_25/sky130_fd_sc_hs__nand2_1_37/B prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_1/a_651_503#
+ prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_27/a_376_368# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_4/a_544_485#
+ prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_67/a_376_368# prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_27/X
+ prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_1/X prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_59/a_138_385#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_29/a_1178_124# prbs_generator_syn_25/m3_13600_2871#
+ prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_5/a_230_79# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_23/a_206_368#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_61/a_206_368# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_17/a_544_485#
+ prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_15/a_230_79# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_25/a_696_458#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_55/a_544_485# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_32/a_735_102#
+ prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_29/a_293_74# prbs_generator_syn_25/sky130_fd_sc_hs__nand2_1_17/a_117_74#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_69/a_1034_424# prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_29/a_112_119#
+ prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_37/X prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_31/B
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_19/a_1034_424# prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_33/A
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_9/a_206_368# prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_57/a_376_368#
+ prbs_generator_syn_25/sky130_fd_sc_hs__sdlclkp_2_1/a_706_317# prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_11/B
+ prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_1/a_52_123# prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_39/B
+ prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_21/a_132_392# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_13/a_206_368#
+ prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_43/a_52_123# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_51/a_206_368#
+ prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_47/X prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_23/a_437_503#
+ prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_11/a_52_123# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_61/a_437_503#
+ prbs_generator_syn_25/sky130_fd_sc_hs__nor2b_1_7/Y prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_51/A
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_15/a_696_458# prbs_generator_syn_25/sky130_fd_sc_hs__nor2b_1_5/Y
+ prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_9/a_230_79# prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_25/X
+ prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_19/a_112_119# prbs_generator_syn_25/sky130_fd_sc_hs__nand2_1_45/B
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_5/a_1178_124# prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_19/a_230_79#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_41/a_1226_296# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_59/a_1226_296#
+ prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_63/a_230_79# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_51/Q
+ prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_7/a_132_392# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_9/a_437_503#
+ prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_46/a_376_368# prbs_generator_syn_25/sky130_fd_sc_hs__nand2_1_33/a_117_74#
+ prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_11/a_293_74# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_27/a_1178_124#
+ prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_11/a_132_392# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_13/a_437_503#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_51/a_437_503# prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_5/a_52_123#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_35/a_544_485# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_73/a_651_503#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_45/a_696_458# prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_15/a_52_123#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_47/a_1141_508# prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_47/a_112_119#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_4/a_1178_124# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_17/a_1034_424#
+ prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_23/B prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_37/a_376_368#
+ prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_15/B prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_7/Y
+ prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_29/a_138_385# prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_33/a_230_79#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_25/a_1178_124# prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_47/a_293_74#
+ prbs_generator_syn_25/sky130_fd_sc_hs__nand2_1_37/a_117_74# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_33/a_206_368#
+ prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_15/a_293_74# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_71/a_206_368#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_25/a_544_485# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_67/a_1034_424#
+ prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_13/a_222_392# prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_9/a_52_123#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_15/a_1034_424# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_57/a_1226_296#
+ prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_19/a_52_123# prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_23/X
+ prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_63/a_52_123# prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_19/a_138_385#
+ prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_9/a_376_368# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_21/a_206_368#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_33/a_437_503# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_71/a_437_503#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_53/a_651_503# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_15/a_544_485#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_63/a_696_458# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_65/a_1034_424#
+ prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_19/a_293_74# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_45/a_1141_508#
+ prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_27/a_112_119# prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_67/a_112_119#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_1/a_1178_124# prbs_generator_syn_25/sky130_fd_sc_hs__conb_1_1/a_21_290#
+ prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_63/a_293_74# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_8/a_206_368#
+ prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_17/a_376_368# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_63/a_27_74#
+ prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_21/A prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_55/a_376_368#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_1/a_696_458# prbs_generator_syn_25/sky130_fd_sc_hs__nor2b_1_1/a_278_368#
+ prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_47/a_138_385# prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_33/a_52_123#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_9/a_1034_424# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_21/a_437_503#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_1/a_27_74# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_43/a_651_503#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_1/Q prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_45/a_544_485#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_69/a_735_102# prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_57/a_112_119#
+ prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_31/a_222_392# prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_13/A
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_55/a_1226_296# prbs_generator_syn_25/sky130_fd_sc_hs__nand2_2_5/a_27_74#
+ prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_53/a_230_79# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_8/a_437_503#
+ prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_67/a_293_74# prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_33/a_293_74#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_7/a_735_102# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_23/a_1178_124#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_41/a_206_368# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_8/a_1034_424#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_63/a_1034_424# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_59/a_735_102#
+ prbs_generator_syn_25/sky130_fd_sc_hs__nand2_1_5/B prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_43/a_1141_508#
+ prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_46/a_112_119# prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_61/a_222_392#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_13/a_1034_424# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_73/a_1178_124#
+ prbs_generator_syn_25/sky130_fd_sc_hs__nand2_1_27/B prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_13/B
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_57/a_27_74# prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_57/a_230_79#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_21/a_1178_124# prbs_generator_syn_25/sky130_fd_sc_hs__nor2b_1_1/a_27_112#
+ prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_27/a_138_385# prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_23/a_230_79#
+ prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_67/a_138_385# prbs_generator_syn_25/sky130_fd_sc_hs__nand2_1_41/B
+ prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_9/a_222_392# prbs_generator_syn_25/sky130_fd_sc_hs__nand2_1_27/a_117_74#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_32/a_206_368# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_23/a_651_503#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_41/a_437_503# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_73/a_27_74#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_61/a_651_503# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_63/a_544_485#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_49/a_735_102# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_73/a_696_458#
+ prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_37/a_112_119# prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_51/a_222_392#
+ prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_43/X prbs_generator_syn_25/sky130_fd_sc_hs__nand2_2_1/B
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_9/a_651_503# prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_53/a_52_123#
+ prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_49/X prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_25/a_376_368#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_1/a_544_485# prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_65/a_376_368#
+ prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_57/a_138_385# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_27/a_27_74#
+ prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_39/a_132_392# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_7/a_1034_424#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_13/a_651_503# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_32/a_437_503#
+ prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_27/a_230_79# prbs_generator_syn_25/m3_13600_12265#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_51/a_651_503# prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_59/B
+ prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_47/A prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_61/a_1034_424#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_41/a_1141_508# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_59/a_1141_508#
+ prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_41/a_222_392# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_53/a_1226_296#
+ prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_3/A prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_71/a_1178_124#
+ prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_9/a_112_119# prbs_generator_syn_25/sky130_fd_sc_hs__nand2_1_3/a_117_74#
+ prbs_generator_syn_25/m3_13600_8483# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_39/a_1178_124#
+ prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_57/a_52_123# prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_46/a_138_385#
+ prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_23/a_52_123# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_67/a_27_74#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_53/a_696_458# prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_17/a_112_119#
+ prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_11/A prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_55/a_112_119#
+ prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_1/A prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_51/a_1226_296#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_29/a_1034_424# prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_59/A
+ prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_23/A prbs_generator_syn_25/sky130_fd_sc_hs__nand2_1_39/B
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_5/a_27_74# prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_57/a_293_74#
+ prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_37/a_138_385# prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_59/a_132_392#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_33/a_651_503# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_71/a_651_503#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_43/a_696_458# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_73/a_544_485#
+ prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_27/a_52_123# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_57/a_1141_508#
+ prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_21/a_222_392# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_35/a_27_74#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_69/a_1226_296# prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_37/B
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_19/a_1226_296# prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_35/a_376_368#
+ prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_47/a_230_79# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_37/a_1178_124#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_5/a_1034_424# prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_49/a_132_392#
+ prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_7/a_222_392# prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_27/a_293_74#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_21/a_651_503# prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_9/a_138_385#
+ prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_11/a_222_392# prbs_generator_syn_25/m3_13600_14095#
+ prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_50/A prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_27/a_1034_424#
+ prbs_generator_syn_25/sky130_fd_sc_hs__nand2_1_13/B prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_8/a_651_503#
+ prbs_generator_syn_25/m3_13600_9703# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_35/a_1178_124#
+ prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_17/a_138_385# prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_55/a_138_385#
+ prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_7/a_230_79# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_4/a_1034_424#
+ prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_7/a_376_368# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_69/a_206_368#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_23/a_696_458# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_53/a_544_485#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_39/a_735_102# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_61/a_696_458#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_55/a_1141_508# prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_25/a_112_119#
+ prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_65/a_112_119# prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_43/a_293_74#
+ prbs_generator_syn_25/sky130_fd_sc_hs__nand2_1_57/B prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_25/a_1034_424#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_7/a_206_368# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_17/a_1226_296#
+ prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_15/a_376_368# prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_53/a_376_368#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_9/a_696_458# prbs_generator_syn_25/m3_13600_431#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_45/a_27_74# prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_47/a_52_123#
+ prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_29/a_132_392# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_59/a_206_368#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_69/a_437_503# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_41/a_651_503#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_43/a_544_485# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_13/a_696_458#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_29/a_735_102# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_51/a_696_458#
+ prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_61/Y prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_67/a_1226_296#
+ prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_5/a_132_392# prbs_generator_syn_25/sky130_fd_sc_hs__and2b_2_1/a_198_48#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_7/a_437_503# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_15/a_1226_296#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_69/a_27_74# prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_46/a_293_74#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_1/a_1034_424# prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_19/a_132_392#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_49/a_206_368# prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_7/a_52_123#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_59/a_437_503# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_32/a_651_503#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_7/a_27_74# prbs_generator_syn_25/sky130_fd_sc_hs__nand2_2_1/a_27_74#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_19/a_735_102# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_57/a_735_102#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_65/a_1226_296# prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_37/A
+ prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_33/a_376_368# prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_37/a_230_79#
+ prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_25/a_138_385# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_39/a_27_74#
+ prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_65/a_138_385# prbs_generator_syn_25/sky130_fd_sc_hs__nor2b_1_9/a_278_368#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_49/a_437_503# prbs_generator_syn_25/sky130_fd_sc_hs__and2b_2_1/a_505_74#
+ prbs_generator_syn_25/sky130_fd_sc_hs__nand2_1_51/a_117_74# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_23/a_544_485#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_33/a_696_458# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_61/a_544_485#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_9/a_1226_296# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_53/a_1141_508#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_71/a_696_458# prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_35/a_112_119#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_23/a_1034_424# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_9/a_544_485#
+ prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_63/a_376_368# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_33/a_1178_124#
+ prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_5/a_376_368# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_13/a_544_485#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_73/a_1034_424# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_21/a_696_458#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_51/a_544_485# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_8/a_1226_296#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_51/a_1141_508# prbs_generator_syn_25/sky130_fd_sc_hs__nand2_1_55/a_117_74#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_21/a_1034_424# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_63/a_1226_296#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_23/a_27_74# prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_7/a_112_119#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_13/a_1226_296# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_8/a_696_458#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_32/a_1178_124# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_49/a_1178_124#
+ prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_37/a_52_123# prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_27/a_132_392#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_71/Q prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_67/a_735_102#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_69/a_1141_508# prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_15/a_112_119#
+ prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_53/a_112_119# prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_39/a_222_392#
+ prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_55/a_230_79# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_19/a_1141_508#
+ prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_37/a_293_74# prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_43/a_376_368#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_5/a_735_102# prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_35/a_138_385#
+ prbs_generator_syn_25/sky130_fd_sc_hs__sdlclkp_2_1/a_114_424# prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_57/a_132_392#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_71/a_1034_424# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_7/a_1226_296#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_33/a_544_485# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_41/a_696_458#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_71/a_544_485# prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_21/B
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_61/a_1226_296# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_39/a_1034_424#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_17/a_27_74# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_9/a_27_74#
+ prbs_generator_syn_25/sky130_fd_sc_hs__nor2b_1_5/a_27_112# prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_47/a_132_392#
+ prbs_generator_syn_25/sky130_fd_sc_hs__nor2b_1_8/a_278_368# prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_9/B
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_39/a_206_368# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_33/a_27_74#
+ prbs_generator_syn_25/sky130_fd_sc_hs__nand2_1_41/a_117_74# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_69/a_651_503#
+ prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_51/a_293_74# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_21/a_544_485#
+ prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_7/a_138_385# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_32/a_696_458#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_47/a_735_102# prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_33/a_112_119#
+ prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_59/a_222_392# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_17/a_1141_508#
+ prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_55/a_52_123# prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_3/a_293_74#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_7/a_651_503# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_29/a_1226_296#
+ prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_23/a_376_368# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_8/a_544_485#
+ prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_47/B prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_47/a_1178_124#
+ prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_15/a_138_385# prbs_generator_syn_25/sky130_fd_sc_hs__sdlclkp_2_1/a_1195_374#
+ prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_53/a_138_385# prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_37/a_132_392#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_29/a_206_368# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_39/a_437_503#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_59/a_651_503# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_37/a_735_102#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_67/a_1141_508# prbs_generator_syn_25/sky130_fd_sc_hs__and2b_2_1/a_27_74#
+ prbs_generator_syn_25/sky130_fd_sc_hs__conb_1_1/a_165_290# prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_55/a_293_74#
+ prbs_generator_syn_25/sky130_fd_sc_hs__nand2_1_45/a_117_74# prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_63/a_112_119#
+ prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_49/a_222_392# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_37/a_1034_424#
+ prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_23/a_293_74# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_15/a_1141_508#
+ prbs_generator_syn_25/sky130_fd_sc_hs__nand2_1_5/a_117_74# prbs_generator_syn_25/m3_13600_13485#
+ prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_5/a_112_119# prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_13/a_376_368#
+ prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_51/a_376_368# prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_7/a_293_74#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_19/a_206_368# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_57/a_206_368#
+ prbs_generator_syn_25/sky130_fd_sc_hs__sdlclkp_2_1/a_318_74# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_29/a_437_503#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_49/a_651_503# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_25/a_27_74#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_5/a_1226_296# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_41/a_544_485#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_27/a_735_102# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_65/a_1141_508#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_65/a_735_102# prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_3/a_230_79#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_35/a_1034_424# prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_13/a_230_79#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_41/a_27_74# prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_3/a_132_392#
+ prbs_generator_syn_25/sky130_fd_sc_hs__nand2_1_49/a_117_74# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_27/a_1226_296#
+ prbs_generator_syn_25/sky130_fd_sc_hs__nand2_1_15/a_117_74# prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_41/a_376_368#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_45/a_1178_124# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_4/a_735_102#
+ prbs_generator_syn_25/sky130_fd_sc_hs__nand2_1_9/a_117_74# prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_33/a_138_385#
+ prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_17/a_132_392# prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_55/a_132_392#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_9/a_1141_508# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_19/a_437_503#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_57/a_437_503# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_4/a_1226_296#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_32/a_544_485# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_17/a_735_102#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_55/a_735_102# prbs_generator_syn_25/m3_13600_2261#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_65/a_27_74# prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_29/a_222_392#
+ prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_43/a_112_119# prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_19/X
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_25/a_1226_296# prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_31/a_376_368#
+ prbs_generator_syn_25/sky130_fd_sc_hs__or2_1_1/a_63_368# prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_17/a_230_79#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_4/a_27_74# prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_61/a_230_79#
+ prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_63/a_138_385# prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_5/a_222_392#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_8/a_1141_508# prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_41/a_293_74#
+ prbs_generator_syn_25/sky130_fd_sc_hs__nand2_1_31/a_117_74# prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_5/a_138_385#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_63/a_1141_508# prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_19/a_222_392#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_13/a_1141_508# prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_3/a_52_123#
+ prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_13/a_52_123# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_43/a_1178_124#
+ prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_61/a_376_368# prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_35/a_132_392#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_67/a_206_368# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_1/a_1226_296#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_69/a_696_458# prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_31/a_230_79#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_35/a_735_102# prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_23/a_112_119#
+ prbs_generator_syn_25/sky130_fd_sc_hs__nand2_1_35/a_117_74# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_59/a_27_74#
+ prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_13/a_293_74# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_5/a_206_368#
+ prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_50/a_376_368# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_7/a_696_458#
+ prbs_generator_syn_25/sky130_fd_sc_hs__nor2b_1_7/a_278_368# prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_17/a_52_123#
+ prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_43/a_138_385# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_7/a_1141_508#
+ prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_61/a_52_123# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_67/a_437_503#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_61/a_1141_508# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_25/a_735_102#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_59/a_696_458# prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_13/a_112_119#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_33/a_1034_424# prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_51/a_112_119#
+ prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_35/a_230_79# prbs_generator_syn_25/m3_13600_4091#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_23/a_1226_296# prbs_generator_syn_25/sky130_fd_sc_hs__nand2_1_39/a_117_74#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_29/a_27_74# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_5/a_437_503#
+ prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_17/a_293_74# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_41/a_1178_124#
+ prbs_generator_syn_25/sky130_fd_sc_hs__or2_1_1/a_152_368# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_59/a_1178_124#
+ prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_61/a_293_74# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_47/a_206_368#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_39/a_651_503# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_49/a_696_458#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_15/a_735_102# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_32/a_1034_424#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_73/a_1226_296# prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_27/a_222_392#
+ prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_41/a_112_119# prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_31/a_52_123#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_49/a_1034_424# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_29/a_1141_508#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_21/a_1226_296# prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_39/a_230_79#
+ prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_23/a_138_385# prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_51/a_230_79#
+ prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_45/a_132_392# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_37/a_206_368#
+ prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_65/a_293_74# prbs_generator_syn_25/sky130_fd_sc_hs__nand2_1_53/a_117_74#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_47/a_437_503# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_29/a_651_503#
+ prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_31/a_293_74# prbs_generator_syn_25/sky130_fd_sc_hs__nand2_1_21/a_117_74#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_69/a_544_485# prbs_generator_syn_25/sky130_fd_sc_hs__clkbuf_16_1/a_114_74#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_45/a_735_102# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_13/a_27_74#
+ prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_31/a_112_119# prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_57/a_222_392#
+ prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_35/a_52_123# prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_21/a_376_368#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_7/a_544_485# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_57/a_1178_124#
+ prbs_generator_syn_25/m3_13600_6043# prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_13/a_138_385#
+ prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_51/a_138_385# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_5/a_1141_508#
+ prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_3/a_376_368# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_27/a_206_368#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_65/a_206_368# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_37/a_437_503#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_19/a_651_503# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_57/a_651_503#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_59/a_544_485# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_71/a_1226_296#
+ prbs_generator_syn_25/sky130_fd_sc_hs__nand2_1_25/a_117_74# prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_61/a_112_119#
+ prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_47/a_222_392# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_27/a_1141_508#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_53/a_27_74# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_4/a_206_368#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_39/a_1226_296# prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_11/a_376_368#
+ prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_39/a_52_123# prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_41/a_138_385#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_4/a_1141_508# prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_25/a_132_392#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_17/a_206_368# prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_41/A
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_55/a_206_368# prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_51/a_52_123#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_27/a_437_503# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_65/a_437_503#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_49/a_544_485# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_63/a_735_102#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_47/a_1034_424# prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_50/a_112_119#
+ prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_37/a_222_392# prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_59/a_230_79#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_25/a_1141_508# prbs_generator_syn_25/sky130_fd_sc_hs__nor2b_1_4/a_27_112#
+ prbs_generator_syn_25/sky130_fd_sc_hs__sdlclkp_2_1/a_685_81# prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_1/a_132_392#
+ prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_39/a_293_74# prbs_generator_syn_25/sky130_fd_sc_hs__nand2_1_29/a_117_74#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_4/a_437_503# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_55/a_1178_124#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_21/a_27_74# prbs_generator_syn_25/m3_13600_12875#
+ prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_50/a_293_74# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_1/a_735_102#
+ prbs_generator_syn_25/sky130_fd_sc_hs__xnor2_1_31/a_138_385# prbs_generator_syn_25/sky130_fd_sc_hs__a22o_1_15/a_132_392#
+ prbs_generator_syn_25/sky130_fd_sc_hs__nand2_1_1/a_117_74# prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_17/a_437_503#
+ prbs_generator_syn_25/sky130_fd_sc_hs__dfxtp_4_55/a_437_503# prbs_generator_syn
Xsky130_fd_sc_hs__conb_1_5 DVSS: DVDD: DVDD: DVSS: prbs_generator_syn_1/eqn[8] prbs_generator_syn_1/eqn[1]
+ sky130_fd_sc_hs__conb_1_5/a_165_290# sky130_fd_sc_hs__conb_1_5/a_21_290# sky130_fd_sc_hs__conb_1
Xsky130_fd_sc_hs__buf_2_101 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__buf_2_91/X sky130_fd_sc_hs__buf_2_101/X
+ sky130_fd_sc_hs__buf_2_101/a_21_260# sky130_fd_sc_hs__buf_2
Xsky130_fd_sc_hs__buf_2_112 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__buf_2_113/A sky130_fd_sc_hs__buf_2_113/X
+ sky130_fd_sc_hs__buf_2_113/a_21_260# sky130_fd_sc_hs__buf_2
Xsky130_fd_sc_hs__buf_2_123 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__buf_2_123/A sky130_fd_sc_hs__buf_2_123/X
+ sky130_fd_sc_hs__buf_2_123/a_21_260# sky130_fd_sc_hs__buf_2
Xsky130_fd_sc_hs__buf_2_134 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__buf_2_135/A sky130_fd_sc_hs__buf_2_135/X
+ sky130_fd_sc_hs__buf_2_135/a_21_260# sky130_fd_sc_hs__buf_2
Xsky130_fd_sc_hs__buf_2_145 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__buf_2_151/X sky130_fd_sc_hs__buf_2_145/X
+ sky130_fd_sc_hs__buf_2_145/a_21_260# sky130_fd_sc_hs__buf_2
Xsky130_fd_sc_hs__buf_2_156 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__buf_2_157/A sky130_fd_sc_hs__buf_2_157/X
+ sky130_fd_sc_hs__buf_2_157/a_21_260# sky130_fd_sc_hs__buf_2
Xsky130_fd_sc_hs__einvp_2_13 DVSS: DVDD: DVDD: DVSS: dout_n sky130_fd_sc_hs__buf_8_1/A
+ sky130_fd_sc_hs__dlrtp_1_15/Q sky130_fd_sc_hs__einvp_2_13/a_263_323# sky130_fd_sc_hs__einvp_2_13/a_36_74#
+ sky130_fd_sc_hs__einvp_2_13/a_27_368# sky130_fd_sc_hs__einvp_2
Xsky130_fd_sc_hs__einvp_2_24 DVSS: DVDD: DVDD: DVSS: dout_n sky130_fd_sc_hs__einvp_2_9/A
+ sky130_fd_sc_hs__dlrtp_1_19/Q sky130_fd_sc_hs__einvp_2_25/a_263_323# sky130_fd_sc_hs__einvp_2_25/a_36_74#
+ sky130_fd_sc_hs__einvp_2_25/a_27_368# sky130_fd_sc_hs__einvp_2
Xsky130_fd_sc_hs__einvp_2_35 DVSS: DVDD: DVDD: DVSS: dout_n sky130_fd_sc_hs__buf_8_1/X
+ sky130_fd_sc_hs__buf_2_123/X sky130_fd_sc_hs__einvp_2_35/a_263_323# sky130_fd_sc_hs__einvp_2_35/a_36_74#
+ sky130_fd_sc_hs__einvp_2_35/a_27_368# sky130_fd_sc_hs__einvp_2
Xsky130_fd_sc_hs__einvp_2_46 DVSS: DVDD: DVDD: DVSS: dout_n sky130_fd_sc_hs__buf_8_1/A
+ sky130_fd_sc_hs__dlrtp_1_33/Q sky130_fd_sc_hs__einvp_2_47/a_263_323# sky130_fd_sc_hs__einvp_2_47/a_36_74#
+ sky130_fd_sc_hs__einvp_2_47/a_27_368# sky130_fd_sc_hs__einvp_2
Xsky130_fd_sc_hs__einvp_2_57 DVSS: DVDD: DVDD: DVSS: dout_p sky130_fd_sc_hs__einvp_2_65/A
+ sky130_fd_sc_hs__dlrtp_1_41/Q sky130_fd_sc_hs__einvp_2_57/a_263_323# sky130_fd_sc_hs__einvp_2_57/a_36_74#
+ sky130_fd_sc_hs__einvp_2_57/a_27_368# sky130_fd_sc_hs__einvp_2
Xsky130_fd_sc_hs__einvp_2_68 DVSS: DVDD: DVDD: DVSS: dout_p sky130_fd_sc_hs__einvp_2_97/A
+ sky130_fd_sc_hs__dlrtp_1_59/Q sky130_fd_sc_hs__einvp_2_69/a_263_323# sky130_fd_sc_hs__einvp_2_69/a_36_74#
+ sky130_fd_sc_hs__einvp_2_69/a_27_368# sky130_fd_sc_hs__einvp_2
Xsky130_fd_sc_hs__einvp_2_79 DVSS: DVDD: DVDD: DVSS: dout_p sky130_fd_sc_hs__einvp_2_97/A
+ sky130_fd_sc_hs__dlrtp_1_67/Q sky130_fd_sc_hs__einvp_2_79/a_263_323# sky130_fd_sc_hs__einvp_2_79/a_36_74#
+ sky130_fd_sc_hs__einvp_2_79/a_27_368# sky130_fd_sc_hs__einvp_2
Xsky130_fd_sc_hs__or2b_2_5 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__or2b_2_5/X sky130_fd_sc_hs__or2b_4_3/A
+ sky130_fd_sc_hs__or2b_2_5/A sky130_fd_sc_hs__or2b_2_5/a_470_368# sky130_fd_sc_hs__or2b_2_5/a_27_368#
+ sky130_fd_sc_hs__or2b_2_5/a_187_48# sky130_fd_sc_hs__or2b_2
Xsky130_fd_sc_hs__conb_1_12 DVSS: DVDD: DVDD: DVSS: prbs_generator_syn_9/eqn[9] sky130_fd_sc_hs__conb_1_13/HI
+ sky130_fd_sc_hs__conb_1_13/a_165_290# sky130_fd_sc_hs__conb_1_13/a_21_290# sky130_fd_sc_hs__conb_1
Xsky130_fd_sc_hs__conb_1_23 DVSS: DVDD: DVDD: DVSS: prbs_generator_syn_1/eqn[30] sky130_fd_sc_hs__conb_1_23/HI
+ sky130_fd_sc_hs__conb_1_23/a_165_290# sky130_fd_sc_hs__conb_1_23/a_21_290# sky130_fd_sc_hs__conb_1
Xsky130_fd_sc_hs__conb_1_34 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__conb_1_35/LO
+ sky130_fd_sc_hs__conb_1_35/HI sky130_fd_sc_hs__conb_1_35/a_165_290# sky130_fd_sc_hs__conb_1_35/a_21_290#
+ sky130_fd_sc_hs__conb_1
Xsky130_fd_sc_hs__conb_1_45 DVSS: DVDD: DVDD: DVSS: prbs_generator_syn_3/eqn[30] sky130_fd_sc_hs__conb_1_45/HI
+ sky130_fd_sc_hs__conb_1_45/a_165_290# sky130_fd_sc_hs__conb_1_45/a_21_290# sky130_fd_sc_hs__conb_1
Xsky130_fd_sc_hs__conb_1_56 DVSS: DVDD: DVDD: DVSS: prbs_generator_syn_9/eqn[31] prbs_generator_syn_9/cke
+ sky130_fd_sc_hs__conb_1_57/a_165_290# sky130_fd_sc_hs__conb_1_57/a_21_290# sky130_fd_sc_hs__conb_1
Xsky130_fd_sc_hs__conb_1_67 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__conb_1_67/LO
+ sky130_fd_sc_hs__conb_1_67/HI sky130_fd_sc_hs__conb_1_67/a_165_290# sky130_fd_sc_hs__conb_1_67/a_21_290#
+ sky130_fd_sc_hs__conb_1
Xsky130_fd_sc_hs__conb_1_78 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__conb_1_79/LO
+ sky130_fd_sc_hs__conb_1_79/HI sky130_fd_sc_hs__conb_1_79/a_165_290# sky130_fd_sc_hs__conb_1_79/a_21_290#
+ sky130_fd_sc_hs__conb_1
Xsky130_fd_sc_hs__inv_4_30 DVSS: DVDD: DVDD: DVSS: osc_core_1/pi1_r[3] osc_core_1/pi1_l[3]
+ sky130_fd_sc_hs__inv_4
Xsky130_fd_sc_hs__conb_1_89 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__conb_1_89/LO
+ sky130_fd_sc_hs__conb_1_89/HI sky130_fd_sc_hs__conb_1_89/a_165_290# sky130_fd_sc_hs__conb_1_89/a_21_290#
+ sky130_fd_sc_hs__conb_1
Xsky130_fd_sc_hs__inv_4_41 DVSS: DVDD: DVDD: DVSS: osc_core_1/pi2_r[2] osc_core_1/pi2_l[2]
+ sky130_fd_sc_hs__inv_4
Xsky130_fd_sc_hs__inv_4_52 DVSS: DVDD: DVDD: DVSS: osc_core_1/pi4_r[3] osc_core_1/pi4_l[3]
+ sky130_fd_sc_hs__inv_4
Xsky130_fd_sc_hs__inv_4_63 DVSS: DVDD: DVDD: DVSS: osc_core_1/pi4_r[1] osc_core_1/pi4_l[1]
+ sky130_fd_sc_hs__inv_4
Xsky130_fd_sc_hs__inv_4_74 DVSS: DVDD: DVDD: DVSS: osc_core_1/pi5_r[1] osc_core_1/pi5_l[1]
+ sky130_fd_sc_hs__inv_4
Xsky130_fd_sc_hs__inv_4_85 DVSS: DVDD: DVDD: DVSS: hr_16t4_mux_top_3/din[4] hr_16t4_mux_top_1/din[4]
+ sky130_fd_sc_hs__inv_4
Xsky130_fd_sc_hs__dlrtp_1_14 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__dlrtp_1_15/Q
+ sky130_fd_sc_hs__clkbuf_2_3/X sky130_fd_sc_hs__conb_1_119/HI sky130_fd_sc_hs__buf_2_103/X
+ sky130_fd_sc_hs__dlrtp_1_15/a_216_424# sky130_fd_sc_hs__dlrtp_1_15/a_759_508# sky130_fd_sc_hs__dlrtp_1_15/a_565_74#
+ sky130_fd_sc_hs__dlrtp_1_15/a_27_424# sky130_fd_sc_hs__dlrtp_1_15/a_1045_74# sky130_fd_sc_hs__dlrtp_1_15/a_643_74#
+ sky130_fd_sc_hs__dlrtp_1_15/a_817_48# sky130_fd_sc_hs__dlrtp_1_15/a_568_392# sky130_fd_sc_hs__dlrtp_1_15/a_363_74#
+ sky130_fd_sc_hs__dlrtp_1_15/a_769_74# sky130_fd_sc_hs__dlrtp_1
Xsky130_fd_sc_hs__dlrtp_1_25 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__dlrtp_1_25/Q
+ sky130_fd_sc_hs__clkbuf_2_3/X sky130_fd_sc_hs__conb_1_119/HI sky130_fd_sc_hs__dlrtp_1_25/D
+ sky130_fd_sc_hs__dlrtp_1_25/a_216_424# sky130_fd_sc_hs__dlrtp_1_25/a_759_508# sky130_fd_sc_hs__dlrtp_1_25/a_565_74#
+ sky130_fd_sc_hs__dlrtp_1_25/a_27_424# sky130_fd_sc_hs__dlrtp_1_25/a_1045_74# sky130_fd_sc_hs__dlrtp_1_25/a_643_74#
+ sky130_fd_sc_hs__dlrtp_1_25/a_817_48# sky130_fd_sc_hs__dlrtp_1_25/a_568_392# sky130_fd_sc_hs__dlrtp_1_25/a_363_74#
+ sky130_fd_sc_hs__dlrtp_1_25/a_769_74# sky130_fd_sc_hs__dlrtp_1
Xsky130_fd_sc_hs__dlrtp_1_36 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__dlrtp_1_37/Q
+ sky130_fd_sc_hs__clkbuf_2_3/A sky130_fd_sc_hs__conb_1_121/HI sky130_fd_sc_hs__buf_2_135/X
+ sky130_fd_sc_hs__dlrtp_1_37/a_216_424# sky130_fd_sc_hs__dlrtp_1_37/a_759_508# sky130_fd_sc_hs__dlrtp_1_37/a_565_74#
+ sky130_fd_sc_hs__dlrtp_1_37/a_27_424# sky130_fd_sc_hs__dlrtp_1_37/a_1045_74# sky130_fd_sc_hs__dlrtp_1_37/a_643_74#
+ sky130_fd_sc_hs__dlrtp_1_37/a_817_48# sky130_fd_sc_hs__dlrtp_1_37/a_568_392# sky130_fd_sc_hs__dlrtp_1_37/a_363_74#
+ sky130_fd_sc_hs__dlrtp_1_37/a_769_74# sky130_fd_sc_hs__dlrtp_1
Xsky130_fd_sc_hs__dlrtp_1_47 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__dlrtp_1_47/Q
+ sky130_fd_sc_hs__clkbuf_16_53/A sky130_fd_sc_hs__conb_1_121/HI sky130_fd_sc_hs__buf_2_21/X
+ sky130_fd_sc_hs__dlrtp_1_47/a_216_424# sky130_fd_sc_hs__dlrtp_1_47/a_759_508# sky130_fd_sc_hs__dlrtp_1_47/a_565_74#
+ sky130_fd_sc_hs__dlrtp_1_47/a_27_424# sky130_fd_sc_hs__dlrtp_1_47/a_1045_74# sky130_fd_sc_hs__dlrtp_1_47/a_643_74#
+ sky130_fd_sc_hs__dlrtp_1_47/a_817_48# sky130_fd_sc_hs__dlrtp_1_47/a_568_392# sky130_fd_sc_hs__dlrtp_1_47/a_363_74#
+ sky130_fd_sc_hs__dlrtp_1_47/a_769_74# sky130_fd_sc_hs__dlrtp_1
Xsky130_fd_sc_hs__dlrtp_1_58 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__dlrtp_1_58/Q
+ sky130_fd_sc_hs__clkbuf_16_53/A sky130_fd_sc_hs__conb_1_125/HI sky130_fd_sc_hs__dlrtp_1_58/D
+ sky130_fd_sc_hs__dlrtp_1_58/a_216_424# sky130_fd_sc_hs__dlrtp_1_58/a_759_508# sky130_fd_sc_hs__dlrtp_1_58/a_565_74#
+ sky130_fd_sc_hs__dlrtp_1_58/a_27_424# sky130_fd_sc_hs__dlrtp_1_58/a_1045_74# sky130_fd_sc_hs__dlrtp_1_58/a_643_74#
+ sky130_fd_sc_hs__dlrtp_1_58/a_817_48# sky130_fd_sc_hs__dlrtp_1_58/a_568_392# sky130_fd_sc_hs__dlrtp_1_58/a_363_74#
+ sky130_fd_sc_hs__dlrtp_1_58/a_769_74# sky130_fd_sc_hs__dlrtp_1
Xsky130_fd_sc_hs__dlrtp_1_69 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__dlrtp_1_69/Q
+ sky130_fd_sc_hs__clkbuf_16_53/A sky130_fd_sc_hs__conb_1_129/HI sky130_fd_sc_hs__dlrtp_1_69/D
+ sky130_fd_sc_hs__dlrtp_1_69/a_216_424# sky130_fd_sc_hs__dlrtp_1_69/a_759_508# sky130_fd_sc_hs__dlrtp_1_69/a_565_74#
+ sky130_fd_sc_hs__dlrtp_1_69/a_27_424# sky130_fd_sc_hs__dlrtp_1_69/a_1045_74# sky130_fd_sc_hs__dlrtp_1_69/a_643_74#
+ sky130_fd_sc_hs__dlrtp_1_69/a_817_48# sky130_fd_sc_hs__dlrtp_1_69/a_568_392# sky130_fd_sc_hs__dlrtp_1_69/a_363_74#
+ sky130_fd_sc_hs__dlrtp_1_69/a_769_74# sky130_fd_sc_hs__dlrtp_1
Xsky130_fd_sc_hs__einvp_2_7 DVSS: DVDD: DVDD: DVSS: dout_n sky130_fd_sc_hs__buf_8_1/A
+ sky130_fd_sc_hs__dlrtp_1_3/Q sky130_fd_sc_hs__einvp_2_7/a_263_323# sky130_fd_sc_hs__einvp_2_7/a_36_74#
+ sky130_fd_sc_hs__einvp_2_7/a_27_368# sky130_fd_sc_hs__einvp_2
Xfine_freq_track_1 osc_core_1/p3 sky130_fd_sc_hs__clkbuf_4_89/X sky130_fd_sc_hs__clkbuf_4_91/X
+ sky130_fd_sc_hs__clkbuf_4_93/X sky130_fd_sc_hs__clkbuf_4_95/X sky130_fd_sc_hs__clkbuf_4_97/X
+ sky130_fd_sc_hs__clkbuf_4_99/X osc_core_1/ref_clk qr_4t1_mux_top_1/rst fine_freq_track_1/aux_osc_en
+ fine_freq_track_1/fftl_en sky130_fd_sc_hs__clkbuf_4_65/X sky130_fd_sc_hs__clkbuf_4_61/X
+ sky130_fd_sc_hs__clkbuf_4_63/X sky130_fd_sc_hs__clkinv_2_3/Y sky130_fd_sc_hs__clkbuf_4_67/X
+ sky130_fd_sc_hs__clkbuf_4_53/X sky130_fd_sc_hs__clkbuf_4_57/X sky130_fd_sc_hs__clkbuf_4_59/X
+ sky130_fd_sc_hs__clkbuf_4_55/X sky130_fd_sc_hs__clkbuf_8_15/X sky130_fd_sc_hs__clkbuf_8_17/X
+ sky130_fd_sc_hs__clkbuf_8_19/X sky130_fd_sc_hs__clkbuf_8_13/X sky130_fd_sc_hs__clkbuf_8_21/X
+ sky130_fd_sc_hs__clkbuf_16_19/X sky130_fd_sc_hs__clkbuf_16_17/X sky130_fd_sc_hs__clkbuf_8_23/X
+ sky130_fd_sc_hs__clkbuf_8_25/X sky130_fd_sc_hs__clkbuf_8_27/X sky130_fd_sc_hs__clkbuf_8_29/X
+ sky130_fd_sc_hs__clkbuf_8_31/X sky130_fd_sc_hs__clkbuf_4_41/X sky130_fd_sc_hs__einvp_8_5/A
+ fine_freq_track_1/out_star osc_core_1/delay_con_msb[7] osc_core_1/delay_con_msb[6]
+ osc_core_1/delay_con_msb[5] osc_core_1/delay_con_msb[4] osc_core_1/delay_con_msb[3]
+ osc_core_1/delay_con_msb[2] osc_core_1/delay_con_msb[1] osc_core_1/delay_con_msb[0]
+ osc_core_1/delay_con_lsb[4] osc_core_1/delay_con_lsb[3] osc_core_1/delay_con_lsb[2]
+ osc_core_1/delay_con_lsb[1] osc_core_1/delay_con_lsb[0] DVSS: DVDD: fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_9/a_1827_81#
+ fine_freq_track_1/sky130_fd_sc_hs__nor2b_1_23/Y fine_freq_track_1/sky130_fd_sc_hs__o21a_1_51/B1
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_19/a_498_360# fine_freq_track_1/sky130_fd_sc_hs__inv_4_65/Y
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_79/a_1350_392# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_63/a_789_463#
+ fine_freq_track_1/sky130_fd_sc_hs__dfstp_2_4/a_2022_94# fine_freq_track_1/sky130_fd_sc_hs__nor2_1_35/B
+ fine_freq_track_1/sky130_fd_sc_hs__dfstp_2_7/a_1278_74# fine_freq_track_1/sky130_fd_sc_hs__nor2_1_3/a_116_368#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_15/a_706_463# fine_freq_track_1/sky130_fd_sc_hs__inv_2_7/Y
+ fine_freq_track_1/sky130_fd_sc_hs__a22o_1_27/a_222_392# fine_freq_track_1/sky130_fd_sc_hs__a32oi_1_3/Y
+ fine_freq_track_1/sky130_fd_sc_hs__a22o_1_21/a_52_123# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_3/a_37_78#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_75/a_1678_395# fine_freq_track_1/sky130_fd_sc_hs__inv_4_45/A
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_45/a_834_355# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_37/a_1627_493#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_45/a_319_360# fine_freq_track_1/sky130_fd_sc_hs__fa_2_11/a_1205_79#
+ fine_freq_track_1/sky130_fd_sc_hs__fa_2_1/CIN fine_freq_track_1/sky130_fd_sc_hs__nor2_1_31/Y
+ fine_freq_track_1/sky130_fd_sc_hs__a32oi_1_3/B1 fine_freq_track_1/sky130_fd_sc_hs__nand2_4_13/Y
+ fine_freq_track_1/sky130_fd_sc_hs__nand3_1_1/a_155_74# fine_freq_track_1/sky130_fd_sc_hs__nor2_1_37/B
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_59/a_313_74# fine_freq_track_1/sky130_fd_sc_hs__sdlclkp_1_1/a_114_112#
+ fine_freq_track_1/sky130_fd_sc_hs__nor2b_1_25/Y fine_freq_track_1/sky130_fd_sc_hs__o21a_1_7/A1
+ fine_freq_track_1/sky130_fd_sc_hs__sdlclkp_4_1/a_634_74# fine_freq_track_1/sky130_fd_sc_hs__nor4_1_1/D
+ fine_freq_track_1/sky130_fd_sc_hs__inv_4_63/Y fine_freq_track_1/sky130_fd_sc_hs__inv_4_125/A
+ fine_freq_track_1/sky130_fd_sc_hs__inv_4_59/A fine_freq_track_1/sky130_fd_sc_hs__dfxtp_2_3/a_1217_314#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_25/a_313_74# fine_freq_track_1/sky130_fd_sc_hs__clkbuf_8_1/X
+ fine_freq_track_1/sky130_fd_sc_hs__inv_4_47/A fine_freq_track_1/sky130_fd_sc_hs__o21a_1_5/X
+ fine_freq_track_1/sky130_fd_sc_hs__o21a_1_37/a_376_387# fine_freq_track_1/sky130_fd_sc_hs__inv_4_55/Y
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_39/a_890_138# fine_freq_track_1/sky130_fd_sc_hs__clkbuf_2_1/X
+ fine_freq_track_1/sky130_fd_sc_hs__dfxtp_2_9/a_206_368# fine_freq_track_1/sky130_fd_sc_hs__xnor2_1_3/B
+ fine_freq_track_1/sky130_fd_sc_hs__nor2_1_61/B fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_25/a_125_78#
+ fine_freq_track_1/sky130_fd_sc_hs__o21a_1_77/a_376_387# fine_freq_track_1/sky130_fd_sc_hs__dfsbp_2_1/a_225_74#
+ fine_freq_track_1/sky130_fd_sc_hs__nor2b_1_7/a_27_112# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_7/a_714_127#
+ fine_freq_track_1/sky130_fd_sc_hs__o21a_1_77/a_83_244# fine_freq_track_1/sky130_fd_sc_hs__nand2_1_9/A
+ fine_freq_track_1/sky130_fd_sc_hs__nand2_1_113/a_117_74# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_15/a_38_78#
+ fine_freq_track_1/sky130_fd_sc_hs__inv_4_135/Y fine_freq_track_1/sky130_fd_sc_hs__nand4_2_1/B
+ fine_freq_track_1/sky130_fd_sc_hs__inv_4_73/A fine_freq_track_1/sky130_fd_sc_hs__nand2_1_47/B
+ fine_freq_track_1/sky130_fd_sc_hs__nor2_1_43/a_116_368# fine_freq_track_1/sky130_fd_sc_hs__a22oi_1_19/a_339_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_5/a_1224_74# fine_freq_track_1/sky130_fd_sc_hs__xnor2_1_15/Y
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_43/D fine_freq_track_1/sky130_fd_sc_hs__inv_4_137/A
+ fine_freq_track_1/sky130_fd_sc_hs__dfstp_2_1/CLK fine_freq_track_1/sky130_fd_sc_hs__nor2_1_41/Y
+ fine_freq_track_1/sky130_fd_sc_hs__dfxtp_4_2/a_1141_508# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_5/a_124_78#
+ fine_freq_track_1/sky130_fd_sc_hs__inv_4_103/A fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_23/D
+ fine_freq_track_1/sky130_fd_sc_hs__nor2_1_45/B fine_freq_track_1/sky130_fd_sc_hs__nor2b_1_45/a_27_112#
+ fine_freq_track_1/sky130_fd_sc_hs__dfstp_2_7/Q fine_freq_track_1/sky130_fd_sc_hs__a31oi_2_1/Y
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_81/a_699_463# fine_freq_track_1/sky130_fd_sc_hs__o22ai_1_9/B1
+ fine_freq_track_1/sky130_fd_sc_hs__xnor2_1_1/B fine_freq_track_1/sky130_fd_sc_hs__nor2b_1_19/a_278_368#
+ fine_freq_track_1/sky130_fd_sc_hs__nor3_1_5/Y fine_freq_track_1/sky130_fd_sc_hs__inv_4_87/Y
+ fine_freq_track_1/sky130_fd_sc_hs__nand2_1_77/a_117_74# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_43/a_841_401#
+ fine_freq_track_1/sky130_fd_sc_hs__o22ai_1_9/a_27_74# fine_freq_track_1/sky130_fd_sc_hs__inv_4_133/Y
+ fine_freq_track_1/sky130_fd_sc_hs__nor3_1_1/a_198_368# fine_freq_track_1/sky130_fd_sc_hs__o21a_1_71/A1
+ fine_freq_track_1/sky130_fd_sc_hs__a22o_1_3/a_222_392# fine_freq_track_1/sky130_fd_sc_hs__a21oi_1_97/Y
+ fine_freq_track_1/sky130_fd_sc_hs__nor3_1_13/A fine_freq_track_1/sky130_fd_sc_hs__inv_4_17/Y
+ fine_freq_track_1/sky130_fd_sc_hs__nand2_1_43/a_117_74# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_45/a_812_138#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_23/a_856_304# fine_freq_track_1/sky130_fd_sc_hs__o31ai_1_1/a_119_368#
+ fine_freq_track_1/sky130_fd_sc_hs__fa_2_21/a_27_79# fine_freq_track_1/sky130_fd_sc_hs__o211ai_1_7/a_311_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_23/a_850_127# fine_freq_track_1/sky130_fd_sc_hs__nor3_1_13/C
+ fine_freq_track_1/sky130_fd_sc_hs__nand2_1_11/a_117_74# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_17/a_33_74#
+ fine_freq_track_1/sky130_fd_sc_hs__nand4_1_5/C fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_29/a_1647_81#
+ fine_freq_track_1/sky130_fd_sc_hs__fa_2_21/a_484_347# fine_freq_track_1/sky130_fd_sc_hs__dfxtp_2_3/a_695_459#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_81/a_124_78# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_31/a_38_78#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_67/a_1647_81# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_29/a_1224_74#
+ fine_freq_track_1/sky130_fd_sc_hs__inv_4_75/A fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_5/a_38_78#
+ fine_freq_track_1/sky130_fd_sc_hs__nand2_1_5/a_117_74# fine_freq_track_1/sky130_fd_sc_hs__nor2_1_51/Y
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_41/a_507_368# fine_freq_track_1/sky130_fd_sc_hs__or3b_2_1/a_458_368#
+ fine_freq_track_1/sky130_fd_sc_hs__o21a_1_71/a_320_74# fine_freq_track_1/sky130_fd_sc_hs__a21oi_1_27/a_29_368#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_43/Q_N fine_freq_track_1/sky130_fd_sc_hs__nor2_1_37/Y
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_53/a_789_463# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_47/a_498_360#
+ fine_freq_track_1/sky130_fd_sc_hs__dfstp_2_1/a_767_384# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_49/a_1547_508#
+ fine_freq_track_1/sky130_fd_sc_hs__a22o_1_17/a_222_392# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_35/Q_N
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_73/a_1678_395# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_35/a_834_355#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_91/a_37_78# fine_freq_track_1/sky130_fd_sc_hs__fa_2_7/a_27_79#
+ fine_freq_track_1/sky130_fd_sc_hs__xnor2_1_7/Y fine_freq_track_1/sky130_fd_sc_hs__a21oi_1_9/a_29_368#
+ fine_freq_track_1/sky130_fd_sc_hs__a21oi_1_71/a_29_368# fine_freq_track_1/sky130_fd_sc_hs__xor2_1_5/a_455_87#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_25/Q_N fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_43/D
+ fine_freq_track_1/sky130_fd_sc_hs__inv_4_85/Y fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_73/a_834_355#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_39/a_922_127# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_27/a_1350_392#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_21/D fine_freq_track_1/sky130_fd_sc_hs__maj3_1_3/a_598_384#
+ fine_freq_track_1/sky130_fd_sc_hs__nor2_1_47/B fine_freq_track_1/sky130_fd_sc_hs__o21a_1_15/A1
+ fine_freq_track_1/sky130_fd_sc_hs__inv_4_65/A fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_33/a_33_74#
+ fine_freq_track_1/sky130_fd_sc_hs__a22oi_1_15/Y fine_freq_track_1/sky130_fd_sc_hs__o21a_1_9/a_83_244#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_23/a_1678_395# fine_freq_track_1/sky130_fd_sc_hs__o21a_1_27/a_376_387#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_41/a_2026_424# fine_freq_track_1/sky130_fd_sc_hs__inv_4_37/A
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_23/a_832_118# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_29/a_890_138#
+ fine_freq_track_1/sky130_fd_sc_hs__a22oi_1_21/Y fine_freq_track_1/sky130_fd_sc_hs__o21a_1_67/a_376_387#
+ fine_freq_track_1/sky130_fd_sc_hs__maj3_1_1/a_595_136# fine_freq_track_1/sky130_fd_sc_hs__or2_1_3/A
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_25/a_1465_471# fine_freq_track_1/sky130_fd_sc_hs__a21oi_1_17/Y
+ fine_freq_track_1/sky130_fd_sc_hs__inv_4_45/Y fine_freq_track_1/sky130_fd_sc_hs__nor3_1_5/A
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_67/a_890_138# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_13/D
+ fine_freq_track_1/sky130_fd_sc_hs__xor2_1_11/B fine_freq_track_1/sky130_fd_sc_hs__o21a_1_35/X
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_57/a_2010_409# fine_freq_track_1/sky130_fd_sc_hs__nor4_1_1/C
+ fine_freq_track_1/sky130_fd_sc_hs__a21oi_1_57/a_117_74# fine_freq_track_1/sky130_fd_sc_hs__or3b_2_1/B
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_37/a_817_508# fine_freq_track_1/sky130_fd_sc_hs__a211oi_1_1/Y
+ fine_freq_track_1/sky130_fd_sc_hs__nor2_1_97/A fine_freq_track_1/sky130_fd_sc_hs__inv_4_79/Y
+ fine_freq_track_1/sky130_fd_sc_hs__dfxtp_4_9/a_27_74# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_41/a_910_118#
+ fine_freq_track_1/sky130_fd_sc_hs__nor2_1_33/a_116_368# fine_freq_track_1/sky130_fd_sc_hs__inv_4_43/Y
+ fine_freq_track_1/sky130_fd_sc_hs__nor2_1_71/a_116_368# fine_freq_track_1/sky130_fd_sc_hs__nand2_2_3/A
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_7/a_699_463# fine_freq_track_1/sky130_fd_sc_hs__nand2_2_3/a_27_74#
+ fine_freq_track_1/sky130_fd_sc_hs__inv_4_41/Y fine_freq_track_1/sky130_fd_sc_hs__o21ai_2_1/B1
+ fine_freq_track_1/sky130_fd_sc_hs__a31oi_2_1/A1 fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_71/a_699_463#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_31/a_300_74# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_59/D
+ fine_freq_track_1/sky130_fd_sc_hs__a21oi_1_105/a_29_368# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_73/a_313_74#
+ fine_freq_track_1/sky130_fd_sc_hs__nor2_1_87/Y fine_freq_track_1/sky130_fd_sc_hs__nand2_1_117/a_117_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_37/a_1624_74# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_1/a_319_360#
+ fine_freq_track_1/sky130_fd_sc_hs__nor3_1_9/Y fine_freq_track_1/sky130_fd_sc_hs__inv_4_129/A
+ fine_freq_track_1/sky130_fd_sc_hs__dfstp_2_5/a_27_74# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_3/a_1736_119#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_35/a_812_138# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_41/a_313_74#
+ fine_freq_track_1/sky130_fd_sc_hs__inv_4_69/A fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_37/D
+ fine_freq_track_1/sky130_fd_sc_hs__inv_4_129/Y fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_3/a_1266_119#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_73/a_812_138# fine_freq_track_1/sky130_fd_sc_hs__nor2_1_35/Y
+ fine_freq_track_1/sky130_fd_sc_hs__fa_2_3/a_27_378# fine_freq_track_1/sky130_fd_sc_hs__o21a_1_15/a_83_244#
+ fine_freq_track_1/sky130_fd_sc_hs__or2_1_1/A fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_9/a_124_78#
+ fine_freq_track_1/sky130_fd_sc_hs__xor2_1_9/A fine_freq_track_1/sky130_fd_sc_hs__inv_4_77/Y
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_19/a_1647_81# fine_freq_track_1/sky130_fd_sc_hs__maj3_1_1/A
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_87/a_1627_493# fine_freq_track_1/sky130_fd_sc_hs__o21a_1_23/A1
+ fine_freq_track_1/sky130_fd_sc_hs__nor4_1_3/Y fine_freq_track_1/sky130_fd_sc_hs__nor2_2_1/Y
+ fine_freq_track_1/sky130_fd_sc_hs__inv_4_55/A fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_45/a_37_78#
+ fine_freq_track_1/sky130_fd_sc_hs__inv_4_113/Y fine_freq_track_1/sky130_fd_sc_hs__maj3_1_3/A
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_19/a_1224_74# fine_freq_track_1/sky130_fd_sc_hs__fa_2_3/CIN
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_31/a_507_368# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_77/a_1350_392#
+ fine_freq_track_1/sky130_fd_sc_hs__nor4_1_1/a_342_368# fine_freq_track_1/sky130_fd_sc_hs__o21a_1_65/B1
+ fine_freq_track_1/sky130_fd_sc_hs__xor2_1_11/a_455_87# fine_freq_track_1/sky130_fd_sc_hs__xor2_1_9/a_158_392#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_47/a_1547_508# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_83/a_789_463#
+ fine_freq_track_1/sky130_fd_sc_hs__a22oi_1_5/Y fine_freq_track_1/sky130_fd_sc_hs__inv_4_11/A
+ fine_freq_track_1/sky130_fd_sc_hs__nand2_1_15/a_117_74# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_35/a_706_463#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_25/a_319_360# fine_freq_track_1/sky130_fd_sc_hs__inv_4_49/Y
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_63/a_834_355# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_49/a_494_366#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_85/a_124_78# fine_freq_track_1/sky130_fd_sc_hs__and2_2_5/a_31_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_7/a_1934_94# fine_freq_track_1/sky130_fd_sc_hs__nand2_4_9/Y
+ fine_freq_track_1/sky130_fd_sc_hs__fa_2_3/a_701_79# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_29/a_922_127#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_9/a_1598_93# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_25/a_1350_392#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_89/a_494_366# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_7/D
+ fine_freq_track_1/sky130_fd_sc_hs__o211ai_1_9/a_116_368# fine_freq_track_1/sky130_fd_sc_hs__o21a_1_75/a_320_74#
+ fine_freq_track_1/sky130_fd_sc_hs__nor2_1_31/B fine_freq_track_1/sky130_fd_sc_hs__fa_2_11/SUM
+ fine_freq_track_1/sky130_fd_sc_hs__dfxtp_2_1/a_1217_314# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_43/a_1434_74#
+ fine_freq_track_1/sky130_fd_sc_hs__xnor2_1_3/A fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_3/a_1624_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfxtp_4_3/a_206_368# fine_freq_track_1/sky130_fd_sc_hs__nor2_1_27/B
+ fine_freq_track_1/sky130_fd_sc_hs__a22o_1_29/X fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_21/a_1678_395#
+ fine_freq_track_1/sky130_fd_sc_hs__xnor2_1_3/a_112_119# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_13/a_832_118#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_19/a_890_138# fine_freq_track_1/sky130_fd_sc_hs__a21oi_1_75/a_29_368#
+ fine_freq_track_1/sky130_fd_sc_hs__xor2_1_9/a_455_87# fine_freq_track_1/sky130_fd_sc_hs__o21a_1_57/a_376_387#
+ fine_freq_track_1/sky130_fd_sc_hs__a31oi_2_1/a_200_74# fine_freq_track_1/sky130_fd_sc_hs__inv_4_63/A
+ fine_freq_track_1/sky130_fd_sc_hs__xor2_1_9/X fine_freq_track_1/sky130_fd_sc_hs__o21a_1_65/X
+ fine_freq_track_1/sky130_fd_sc_hs__a32oi_1_7/B1 fine_freq_track_1/sky130_fd_sc_hs__fa_2_5/a_992_347#
+ fine_freq_track_1/sky130_fd_sc_hs__or2_1_3/X fine_freq_track_1/sky130_fd_sc_hs__dfxtp_4_5/a_696_458#
+ fine_freq_track_1/sky130_fd_sc_hs__nor2_1_7/Y fine_freq_track_1/sky130_fd_sc_hs__o21ai_1_3/B1
+ fine_freq_track_1/sky130_fd_sc_hs__inv_2_1/A fine_freq_track_1/sky130_fd_sc_hs__nor2_1_23/a_116_368#
+ fine_freq_track_1/sky130_fd_sc_hs__o21a_1_3/a_376_387# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_21/a_699_463#
+ fine_freq_track_1/sky130_fd_sc_hs__nor2b_1_5/a_278_368# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_7/D
+ fine_freq_track_1/sky130_fd_sc_hs__nand2_4_9/a_27_74# fine_freq_track_1/sky130_fd_sc_hs__o21a_1_73/A2
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_61/a_699_463# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_37/a_1550_119#
+ fine_freq_track_1/sky130_fd_sc_hs__nor2_1_107/a_116_368# fine_freq_track_1/sky130_fd_sc_hs__nor2_1_65/Y
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_23/a_841_401# fine_freq_track_1/sky130_fd_sc_hs__nand2_1_59/Y
+ fine_freq_track_1/sky130_fd_sc_hs__fa_2_15/a_336_347# fine_freq_track_1/sky130_fd_sc_hs__nor2_1_63/B
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_1/a_1736_119# fine_freq_track_1/sky130_fd_sc_hs__inv_4_3/A
+ fine_freq_track_1/sky130_fd_sc_hs__inv_4_105/A fine_freq_track_1/sky130_fd_sc_hs__dfxtp_2_9/a_708_101#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_1/a_1266_119# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_63/a_812_138#
+ fine_freq_track_1/sky130_fd_sc_hs__nor2_1_25/B fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_41/a_856_304#
+ fine_freq_track_1/sky130_fd_sc_hs__a32oi_1_9/Y fine_freq_track_1/sky130_fd_sc_hs__o21a_1_25/A1
+ fine_freq_track_1/sky130_fd_sc_hs__fa_2_15/a_27_79# fine_freq_track_1/sky130_fd_sc_hs__o21a_1_27/X
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_41/a_850_127# fine_freq_track_1/sky130_fd_sc_hs__o31ai_1_1/B1
+ fine_freq_track_1/sky130_fd_sc_hs__a21oi_1_109/a_29_368# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_7/a_125_78#
+ fine_freq_track_1/sky130_fd_sc_hs__inv_4_81/Y fine_freq_track_1/sky130_fd_sc_hs__o22ai_1_11/a_340_368#
+ fine_freq_track_1/sky130_fd_sc_hs__fa_2_7/a_683_347# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_47/a_1647_81#
+ fine_freq_track_1/sky130_fd_sc_hs__o22ai_1_1/a_340_368# fine_freq_track_1/sky130_fd_sc_hs__fa_2_19/CIN
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_43/a_1827_81# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_21/a_507_368#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_87/a_1647_81# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_47/a_1224_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfxtp_4_7/D fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_45/a_313_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_9/a_789_463# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_27/a_498_360#
+ fine_freq_track_1/sky130_fd_sc_hs__nor3_1_11/a_114_368# fine_freq_track_1/sky130_fd_sc_hs__nor2_1_27/Y
+ fine_freq_track_1/sky130_fd_sc_hs__xnor2_1_11/a_112_119# fine_freq_track_1/sky130_fd_sc_hs__a222oi_1_3/a_116_392#
+ fine_freq_track_1/sky130_fd_sc_hs__xnor2_1_1/A fine_freq_track_1/sky130_fd_sc_hs__fa_2_7/a_27_378#
+ fine_freq_track_1/sky130_fd_sc_hs__o21a_1_19/a_83_244# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_35/a_1627_493#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_15/a_319_360# fine_freq_track_1/sky130_fd_sc_hs__maj3_1_1/C
+ fine_freq_track_1/sky130_fd_sc_hs__clkbuf_8_1/A fine_freq_track_1/sky130_fd_sc_hs__nor2_1_17/Y
+ fine_freq_track_1/sky130_fd_sc_hs__a21oi_1_121/a_29_368# fine_freq_track_1/sky130_fd_sc_hs__fa_2_17/a_683_347#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_53/a_834_355# fine_freq_track_1/sky130_fd_sc_hs__maj3_1_3/B
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_85/a_37_78# fine_freq_track_1/sky130_fd_sc_hs__nor3_1_3/A
+ fine_freq_track_1/sky130_fd_sc_hs__nor4_1_1/a_144_368# fine_freq_track_1/sky130_fd_sc_hs__fa_2_21/a_1205_79#
+ fine_freq_track_1/sky130_fd_sc_hs__o21a_1_59/A1 fine_freq_track_1/sky130_fd_sc_hs__o21ai_1_7/a_162_368#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_19/a_922_127# fine_freq_track_1/sky130_fd_sc_hs__o21a_1_63/a_83_244#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_79/a_494_366# fine_freq_track_1/sky130_fd_sc_hs__maj3_1_1/a_223_120#
+ fine_freq_track_1/sky130_fd_sc_hs__inv_4_79/A fine_freq_track_1/sky130_fd_sc_hs__inv_4_21/Y
+ fine_freq_track_1/sky130_fd_sc_hs__nand4_1_3/a_373_74# fine_freq_track_1/sky130_fd_sc_hs__fa_2_21/a_487_79#
+ fine_freq_track_1/sky130_fd_sc_hs__nor2_1_9/Y fine_freq_track_1/sky130_fd_sc_hs__inv_4_13/A
+ fine_freq_track_1/sky130_fd_sc_hs__nand2_1_19/a_117_74# fine_freq_track_1/sky130_fd_sc_hs__dfstp_2_1/a_612_74#
+ fine_freq_track_1/sky130_fd_sc_hs__nor3_1_1/Y fine_freq_track_1/sky130_fd_sc_hs__o21a_1_47/a_376_387#
+ fine_freq_track_1/sky130_fd_sc_hs__o21ai_1_3/a_27_74# fine_freq_track_1/sky130_fd_sc_hs__inv_4_125/Y
+ fine_freq_track_1/sky130_fd_sc_hs__dfxtp_4_3/a_437_503# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_23/a_1465_471#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_47/a_890_138# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_89/a_124_78#
+ fine_freq_track_1/sky130_fd_sc_hs__nor2b_1_31/a_27_112# fine_freq_track_1/sky130_fd_sc_hs__nor2_4_1/B
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_55/a_2010_409# fine_freq_track_1/sky130_fd_sc_hs__fa_2_7/a_701_79#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_87/a_890_138# fine_freq_track_1/sky130_fd_sc_hs__nor3_1_9/B
+ fine_freq_track_1/sky130_fd_sc_hs__o21a_1_73/B1 fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_37/D
+ fine_freq_track_1/sky130_fd_sc_hs__nor2_1_13/a_116_368# fine_freq_track_1/sky130_fd_sc_hs__nor4_1_3/B
+ fine_freq_track_1/sky130_fd_sc_hs__or3b_2_1/X fine_freq_track_1/sky130_fd_sc_hs__nor3_1_11/B
+ fine_freq_track_1/sky130_fd_sc_hs__inv_4_39/A fine_freq_track_1/sky130_fd_sc_hs__nor2_1_83/B
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_23/a_124_78# fine_freq_track_1/sky130_fd_sc_hs__dfsbp_2_1/a_2221_74#
+ fine_freq_track_1/sky130_fd_sc_hs__fa_2_19/SUM fine_freq_track_1/sky130_fd_sc_hs__nor2b_1_7/Y
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_51/a_699_463# fine_freq_track_1/sky130_fd_sc_hs__nor2_1_91/a_116_368#
+ fine_freq_track_1/sky130_fd_sc_hs__inv_4_67/Y fine_freq_track_1/sky130_fd_sc_hs__nand2_4_7/Y
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_13/a_841_401# fine_freq_track_1/sky130_fd_sc_hs__a32oi_1_7/A1
+ fine_freq_track_1/sky130_fd_sc_hs__a22o_1_13/a_132_392# fine_freq_track_1/sky130_fd_sc_hs__o31ai_1_1/a_203_368#
+ fine_freq_track_1/sky130_fd_sc_hs__o21a_1_75/B1 fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_3/D
+ fine_freq_track_1/sky130_fd_sc_hs__nor2_1_45/Y fine_freq_track_1/sky130_fd_sc_hs__a21oi_1_13/a_29_368#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_41/a_33_74# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_53/a_812_138#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_31/a_856_304# fine_freq_track_1/sky130_fd_sc_hs__nor2_1_5/Y
+ fine_freq_track_1/sky130_fd_sc_hs__nor4_1_1/a_228_368# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_31/a_850_127#
+ fine_freq_track_1/sky130_fd_sc_hs__nor3_1_1/B fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_85/a_1627_493#
+ fine_freq_track_1/sky130_fd_sc_hs__or3b_2_1/a_542_368# fine_freq_track_1/sky130_fd_sc_hs__o21a_1_53/B1
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_37/a_1647_81# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_3/a_1647_81#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_33/a_1827_81# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_39/a_714_127#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_11/a_507_368# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_77/a_1647_81#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_39/a_37_78# fine_freq_track_1/sky130_fd_sc_hs__inv_2_5/Y
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_75/a_1350_392# fine_freq_track_1/sky130_fd_sc_hs__a32oi_1_1/Y
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_17/a_498_360# fine_freq_track_1/sky130_fd_sc_hs__fa_2_11/B
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_31/a_796_463# fine_freq_track_1/sky130_fd_sc_hs__o211ai_1_3/Y
+ fine_freq_track_1/sky130_fd_sc_hs__nor2_1_25/Y fine_freq_track_1/sky130_fd_sc_hs__dfstp_2_1/a_2022_94#
+ fine_freq_track_1/sky130_fd_sc_hs__o22ai_1_11/a_142_368# fine_freq_track_1/sky130_fd_sc_hs__o22ai_1_1/a_142_368#
+ fine_freq_track_1/sky130_fd_sc_hs__nor2_1_1/a_116_368# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_71/a_1678_395#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_39/a_300_74# fine_freq_track_1/sky130_fd_sc_hs__nor2_1_87/B
+ fine_freq_track_1/sky130_fd_sc_hs__fa_2_13/B fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_83/a_834_355#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_69/a_494_366# fine_freq_track_1/sky130_fd_sc_hs__a21oi_1_1/Y
+ fine_freq_track_1/sky130_fd_sc_hs__inv_4_53/Y fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_49/a_922_127#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_23/a_1434_74# fine_freq_track_1/sky130_fd_sc_hs__a21oi_1_43/a_117_74#
+ fine_freq_track_1/sky130_fd_sc_hs__o22ai_1_1/Y fine_freq_track_1/sky130_fd_sc_hs__a32oi_1_3/a_469_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_15/a_313_74# fine_freq_track_1/sky130_fd_sc_hs__dfxtp_4_9/CLK
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_39/a_1678_395# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_33/a_832_118#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_37/a_890_138# fine_freq_track_1/sky130_fd_sc_hs__dfxtp_2_7/a_206_368#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_53/a_37_78# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_15/a_125_78#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_3/a_890_138# fine_freq_track_1/sky130_fd_sc_hs__inv_4_87/A
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_53/a_2010_409# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_77/a_890_138#
+ fine_freq_track_1/sky130_fd_sc_hs__o21a_1_67/a_83_244# fine_freq_track_1/sky130_fd_sc_hs__nand4_2_1/C
+ fine_freq_track_1/sky130_fd_sc_hs__inv_4_59/Y fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_41/D
+ fine_freq_track_1/sky130_fd_sc_hs__nand2_2_1/Y fine_freq_track_1/sky130_fd_sc_hs__nand2_1_103/a_117_74#
+ fine_freq_track_1/sky130_fd_sc_hs__o21a_1_63/A1 fine_freq_track_1/sky130_fd_sc_hs__maj3_1_1/B
+ fine_freq_track_1/sky130_fd_sc_hs__fa_2_3/B fine_freq_track_1/sky130_fd_sc_hs__nor2_1_41/a_116_368#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_7/a_796_463# fine_freq_track_1/sky130_fd_sc_hs__dfsbp_2_1/a_1339_74#
+ fine_freq_track_1/sky130_fd_sc_hs__o21a_1_67/B1 fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_41/a_699_463#
+ fine_freq_track_1/sky130_fd_sc_hs__nand2_1_99/a_117_74# fine_freq_track_1/sky130_fd_sc_hs__nor2_1_81/a_116_368#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_35/a_1550_119# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_5/a_37_78#
+ fine_freq_track_1/sky130_fd_sc_hs__nor2_4_3/a_27_368# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_29/Q_N
+ fine_freq_track_1/sky130_fd_sc_hs__nand2_1_67/a_117_74# fine_freq_track_1/sky130_fd_sc_hs__o21a_1_59/X
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_45/a_1624_74# fine_freq_track_1/sky130_fd_sc_hs__nor2_1_29/Y
+ fine_freq_track_1/sky130_fd_sc_hs__or2_1_3/B fine_freq_track_1/sky130_fd_sc_hs__xnor2_1_5/B
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_27/a_124_78# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_21/a_856_304#
+ fine_freq_track_1/sky130_fd_sc_hs__fa_2_15/B fine_freq_track_1/sky130_fd_sc_hs__dfxtp_2_5/a_431_508#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_83/a_812_138# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_21/a_850_127#
+ fine_freq_track_1/sky130_fd_sc_hs__a22oi_1_3/a_159_74# fine_freq_track_1/sky130_fd_sc_hs__o21a_1_17/a_320_74#
+ fine_freq_track_1/sky130_fd_sc_hs__inv_4_33/Y fine_freq_track_1/sky130_fd_sc_hs__xnor2_1_3/a_138_385#
+ fine_freq_track_1/sky130_fd_sc_hs__nand3_1_1/A fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_23/a_1827_81#
+ fine_freq_track_1/sky130_fd_sc_hs__a21oi_1_49/a_29_368# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_29/a_714_127#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_3/D fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_71/a_124_78#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_9/a_832_118# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_27/a_1224_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_73/a_1350_392# fine_freq_track_1/sky130_fd_sc_hs__nor2_1_99/Y
+ fine_freq_track_1/sky130_fd_sc_hs__o21a_1_61/a_320_74# fine_freq_track_1/sky130_fd_sc_hs__a21oi_1_17/a_29_368#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_21/a_796_463# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_19/a_38_78#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_45/a_1547_508# fine_freq_track_1/sky130_fd_sc_hs__o21a_1_17/X
+ fine_freq_track_1/sky130_fd_sc_hs__inv_4_83/Y fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_33/a_1627_493#
+ fine_freq_track_1/sky130_fd_sc_hs__inv_4_61/A fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_31/D
+ fine_freq_track_1/sky130_fd_sc_hs__xnor2_1_13/A fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_43/a_706_463#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_35/a_319_360# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_9/a_834_355#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_89/a_1678_395# fine_freq_track_1/sky130_fd_sc_hs__fa_2_11/a_27_378#
+ fine_freq_track_1/sky130_fd_sc_hs__a21oi_1_61/a_29_368# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_23/a_1350_392#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_59/a_494_366# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_79/a_37_78#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_13/a_1434_74# fine_freq_track_1/sky130_fd_sc_hs__maj3_1_1/a_598_384#
+ fine_freq_track_1/sky130_fd_sc_hs__and2_2_5/X fine_freq_track_1/sky130_fd_sc_hs__o21a_1_17/A1
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_39/a_1482_48# fine_freq_track_1/sky130_fd_sc_hs__fa_2_3/A
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_37/a_1678_395# fine_freq_track_1/sky130_fd_sc_hs__o22ai_1_7/A1
+ fine_freq_track_1/sky130_fd_sc_hs__nor3_1_15/A fine_freq_track_1/sky130_fd_sc_hs__fa_2_21/CIN
+ fine_freq_track_1/sky130_fd_sc_hs__a21oi_1_79/a_117_74# fine_freq_track_1/sky130_fd_sc_hs__fa_2_19/B
+ fine_freq_track_1/sky130_fd_sc_hs__dfxtp_4_5/a_544_485# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_7/a_38_78#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_27/a_120_74# fine_freq_track_1/sky130_fd_sc_hs__nand2_2_1/B
+ fine_freq_track_1/sky130_fd_sc_hs__a21oi_1_47/a_117_74# fine_freq_track_1/sky130_fd_sc_hs__o21a_1_33/X
+ fine_freq_track_1/sky130_fd_sc_hs__inv_4_25/A fine_freq_track_1/sky130_fd_sc_hs__fa_2_11/a_701_79#
+ fine_freq_track_1/sky130_fd_sc_hs__a32oi_1_7/a_469_74# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_31/a_699_463#
+ fine_freq_track_1/sky130_fd_sc_hs__xnor2_1_11/a_138_385# fine_freq_track_1/sky130_fd_sc_hs__a21oi_1_91/a_117_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_23/a_37_78# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_21/a_300_74#
+ fine_freq_track_1/sky130_fd_sc_hs__nor2_1_117/a_116_368# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_7/Q
+ fine_freq_track_1/sky130_fd_sc_hs__a211oi_1_1/a_159_74# fine_freq_track_1/sky130_fd_sc_hs__dfxtp_4_3/a_27_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_63/a_313_74# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_33/a_841_401#
+ fine_freq_track_1/sky130_fd_sc_hs__o21a_1_63/X fine_freq_track_1/sky130_fd_sc_hs__o21a_1_63/A2
+ fine_freq_track_1/sky130_fd_sc_hs__nand2_1_107/a_117_74# fine_freq_track_1/sky130_fd_sc_hs__nor2_1_33/Y
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_39/a_1934_94# fine_freq_track_1/sky130_fd_sc_hs__xnor2_1_1/a_376_368#
+ fine_freq_track_1/sky130_fd_sc_hs__nor2b_1_47/a_278_368# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_1/a_120_74#
+ fine_freq_track_1/sky130_fd_sc_hs__inv_2_3/A fine_freq_track_1/sky130_fd_sc_hs__nand4_1_5/A
+ fine_freq_track_1/sky130_fd_sc_hs__o21a_1_37/a_83_244# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_31/a_313_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_9/a_812_138# fine_freq_track_1/sky130_fd_sc_hs__nor2_1_7/B
+ fine_freq_track_1/sky130_fd_sc_hs__nand4_1_1/C fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_11/a_856_304#
+ fine_freq_track_1/sky130_fd_sc_hs__inv_4_123/Y fine_freq_track_1/sky130_fd_sc_hs__o21a_1_71/B1
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_11/a_850_127# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_83/a_1627_493#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_31/a_125_78# fine_freq_track_1/sky130_fd_sc_hs__nor2b_1_19/Y
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_17/a_1647_81# fine_freq_track_1/sky130_fd_sc_hs__fa_2_5/a_1119_79#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_13/a_1827_81# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_9/a_1547_508#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_19/a_714_127# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_57/a_1647_81#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_17/a_1224_74# fine_freq_track_1/sky130_fd_sc_hs__inv_4_19/A
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_1/Q_N fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_9/a_2010_409#
+ fine_freq_track_1/sky130_fd_sc_hs__nor2_1_57/Y fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_3/a_817_508#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_11/a_796_463# fine_freq_track_1/sky130_fd_sc_hs__fa_2_9/SUM
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_43/a_789_463# fine_freq_track_1/sky130_fd_sc_hs__o22ai_1_9/Y
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_91/a_1827_81# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_37/a_498_360#
+ fine_freq_track_1/sky130_fd_sc_hs__nor2b_2_1/Y fine_freq_track_1/sky130_fd_sc_hs__nor3_1_3/Y
+ fine_freq_track_1/sky130_fd_sc_hs__xor2_1_7/a_158_392# fine_freq_track_1/sky130_fd_sc_hs__a22oi_1_7/a_159_74#
+ fine_freq_track_1/sky130_fd_sc_hs__nand2_2_5/a_27_74# fine_freq_track_1/sky130_fd_sc_hs__nor2_1_69/B
+ fine_freq_track_1/sky130_fd_sc_hs__o21ai_1_3/Y fine_freq_track_1/sky130_fd_sc_hs__nor2_1_5/B
+ fine_freq_track_1/sky130_fd_sc_hs__nand3_1_1/B fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_41/D
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_21/a_1350_392# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_75/a_124_78#
+ fine_freq_track_1/sky130_fd_sc_hs__inv_4_41/A fine_freq_track_1/sky130_fd_sc_hs__fa_2_5/SUM
+ fine_freq_track_1/sky130_fd_sc_hs__o21a_1_27/A1 fine_freq_track_1/sky130_fd_sc_hs__nor2_1_99/A
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_7/a_1598_93# fine_freq_track_1/sky130_fd_sc_hs__o21a_1_65/a_320_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_9/a_841_401# fine_freq_track_1/sky130_fd_sc_hs__a22oi_1_1/a_339_74#
+ fine_freq_track_1/sky130_fd_sc_hs__fa_2_23/B fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_1/a_1624_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfxtp_4_2/a_206_368# fine_freq_track_1/sky130_fd_sc_hs__sdlclkp_4_1/a_1292_74#
+ fine_freq_track_1/sky130_fd_sc_hs__o21a_1_17/a_376_387# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_21/a_1465_471#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_17/a_890_138# fine_freq_track_1/sky130_fd_sc_hs__a21oi_1_65/a_29_368#
+ fine_freq_track_1/sky130_fd_sc_hs__or2_1_1/X fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_39/a_1465_471#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_57/a_890_138# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_47/a_37_78#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_9/a_507_368# fine_freq_track_1/sky130_fd_sc_hs__fa_2_3/a_336_347#
+ fine_freq_track_1/sky130_fd_sc_hs__inv_4_29/A fine_freq_track_1/sky130_fd_sc_hs__nand2_2_5/B
+ fine_freq_track_1/sky130_fd_sc_hs__o21a_1_3/A1 fine_freq_track_1/sky130_fd_sc_hs__dfstp_2_5/a_1566_92#
+ fine_freq_track_1/sky130_fd_sc_hs__nor4_1_1/A fine_freq_track_1/sky130_fd_sc_hs__nand4_2_1/a_304_74#
+ fine_freq_track_1/sky130_fd_sc_hs__nor2_1_21/Y fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_31/a_910_118#
+ fine_freq_track_1/sky130_fd_sc_hs__a32oi_1_1/a_391_74# fine_freq_track_1/sky130_fd_sc_hs__maj3_1_3/C
+ fine_freq_track_1/sky130_fd_sc_hs__nor2_1_63/Y fine_freq_track_1/sky130_fd_sc_hs__inv_4_91/A
+ fine_freq_track_1/sky130_fd_sc_hs__nor2_1_61/a_116_368# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_33/a_1550_119#
+ fine_freq_track_1/sky130_fd_sc_hs__nor2b_1_3/a_278_368# fine_freq_track_1/sky130_fd_sc_hs__fa_2_9/B
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_3/a_498_360# fine_freq_track_1/sky130_fd_sc_hs__nor3_1_9/C
+ fine_freq_track_1/sky130_fd_sc_hs__nor2_1_73/Y fine_freq_track_1/sky130_fd_sc_hs__o31ai_1_3/a_114_74#
+ fine_freq_track_1/sky130_fd_sc_hs__inv_4_109/A fine_freq_track_1/sky130_fd_sc_hs__a22o_1_23/a_132_392#
+ fine_freq_track_1/sky130_fd_sc_hs__fa_2_5/CIN fine_freq_track_1/sky130_fd_sc_hs__inv_4_39/Y
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_29/a_1934_94# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_25/a_1624_74#
+ fine_freq_track_1/sky130_fd_sc_hs__fa_2_15/a_992_347# fine_freq_track_1/sky130_fd_sc_hs__nor2b_1_37/a_278_368#
+ fine_freq_track_1/sky130_fd_sc_hs__dfxtp_2_7/a_708_101# fine_freq_track_1/sky130_fd_sc_hs__a21oi_1_95/a_117_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfxtp_4_5/D fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_7/a_1547_508#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_67/a_313_74# fine_freq_track_1/sky130_fd_sc_hs__xnor2_1_5/Y
+ fine_freq_track_1/sky130_fd_sc_hs__nand2_1_89/Y fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_43/a_120_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_49/a_714_127# fine_freq_track_1/sky130_fd_sc_hs__o31ai_1_3/Y
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_43/a_1547_508# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_35/a_313_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_9/a_2026_424# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_33/a_789_463#
+ fine_freq_track_1/sky130_fd_sc_hs__o21a_1_1/A1 fine_freq_track_1/sky130_fd_sc_hs__nand4_1_1/D
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_81/a_1827_81# fine_freq_track_1/sky130_fd_sc_hs__xor2_1_5/a_355_368#
+ fine_freq_track_1/sky130_fd_sc_hs__inv_2_5/A fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_31/a_1627_493#
+ fine_freq_track_1/sky130_fd_sc_hs__inv_4_99/A fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_7/a_910_118#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_35/a_125_78# fine_freq_track_1/sky130_fd_sc_hs__o21a_1_25/X
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_23/a_706_463# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_87/a_1678_395#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_49/a_1627_493# fine_freq_track_1/sky130_fd_sc_hs__a21oi_1_111/a_29_368#
+ fine_freq_track_1/sky130_fd_sc_hs__inv_4_89/Y fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_19/a_1736_119#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_39/a_494_366# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_19/a_1266_119#
+ fine_freq_track_1/sky130_fd_sc_hs__o21a_1_53/a_83_244# fine_freq_track_1/sky130_fd_sc_hs__inv_4_23/A
+ fine_freq_track_1/sky130_fd_sc_hs__o21a_1_61/A2 fine_freq_track_1/sky130_fd_sc_hs__o21a_1_59/A2
+ fine_freq_track_1/sky130_fd_sc_hs__inv_4_117/Y fine_freq_track_1/sky130_fd_sc_hs__o21ai_1_11/Y
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_33/a_1434_74# fine_freq_track_1/sky130_fd_sc_hs__nor2_1_49/Y
+ fine_freq_track_1/sky130_fd_sc_hs__fa_2_17/a_27_79# fine_freq_track_1/sky130_fd_sc_hs__nor3_1_13/B
+ fine_freq_track_1/sky130_fd_sc_hs__nand3_1_1/C fine_freq_track_1/sky130_fd_sc_hs__xnor2_1_9/Y
+ fine_freq_track_1/sky130_fd_sc_hs__dfxtp_4_2/a_437_503# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_51/a_2010_409#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_41/a_832_118# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_79/a_124_78#
+ fine_freq_track_1/sky130_fd_sc_hs__nor2b_1_21/a_27_112# fine_freq_track_1/sky130_fd_sc_hs__nor2_1_99/B
+ fine_freq_track_1/sky130_fd_sc_hs__o21a_1_75/A2 fine_freq_track_1/sky130_fd_sc_hs__nand2_1_53/a_117_74#
+ fine_freq_track_1/sky130_fd_sc_hs__o21a_1_69/a_320_74# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_27/a_38_78#
+ fine_freq_track_1/sky130_fd_sc_hs__o21a_1_9/X fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_21/a_910_118#
+ fine_freq_track_1/sky130_fd_sc_hs__inv_4_69/Y fine_freq_track_1/sky130_fd_sc_hs__nor3_1_5/a_114_368#
+ fine_freq_track_1/sky130_fd_sc_hs__o21a_1_35/a_320_74# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_11/a_699_463#
+ fine_freq_track_1/sky130_fd_sc_hs__nor2_1_51/a_116_368# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_31/a_1550_119#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_13/a_124_78# fine_freq_track_1/sky130_fd_sc_hs__fa_2_19/a_27_378#
+ fine_freq_track_1/sky130_fd_sc_hs__a21oi_1_69/a_29_368# fine_freq_track_1/sky130_fd_sc_hs__inv_4_133/A
+ fine_freq_track_1/sky130_fd_sc_hs__a22oi_1_21/a_71_368# fine_freq_track_1/sky130_fd_sc_hs__nand2b_1_3/a_27_112#
+ fine_freq_track_1/sky130_fd_sc_hs__o21a_1_7/X fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_19/a_2010_409#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_19/a_1934_94# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_15/a_1624_74#
+ fine_freq_track_1/sky130_fd_sc_hs__a21oi_1_35/a_29_368# fine_freq_track_1/sky130_fd_sc_hs__nor2b_1_27/a_278_368#
+ fine_freq_track_1/sky130_fd_sc_hs__nor2_1_1/Y fine_freq_track_1/sky130_fd_sc_hs__nor4_1_1/B
+ fine_freq_track_1/sky130_fd_sc_hs__a32oi_1_5/a_391_74# fine_freq_track_1/sky130_fd_sc_hs__fa_2_15/SUM
+ fine_freq_track_1/sky130_fd_sc_hs__nand2_1_71/Y fine_freq_track_1/sky130_fd_sc_hs__o21a_1_71/X
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_81/a_1627_493# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_9/a_1434_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_29/a_33_74# fine_freq_track_1/sky130_fd_sc_hs__inv_4_71/A
+ fine_freq_track_1/sky130_fd_sc_hs__nor2_1_101/Y fine_freq_track_1/sky130_fd_sc_hs__o21a_1_9/B1
+ fine_freq_track_1/sky130_fd_sc_hs__sdlclkp_1_1/a_1166_94# fine_freq_track_1/sky130_fd_sc_hs__inv_2_3/Y
+ fine_freq_track_1/sky130_fd_sc_hs__o31ai_1_7/a_114_74# fine_freq_track_1/sky130_fd_sc_hs__a32oi_1_1/a_27_368#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_71/a_1350_392# fine_freq_track_1/sky130_fd_sc_hs__o31ai_1_1/Y
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_7/a_1827_81# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_7/a_2010_409#
+ fine_freq_track_1/sky130_fd_sc_hs__o21a_1_19/X fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_37/a_1224_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_41/a_1547_508# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_23/a_789_463#
+ fine_freq_track_1/sky130_fd_sc_hs__fa_2_19/a_701_79# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_71/a_1827_81#
+ fine_freq_track_1/sky130_fd_sc_hs__o31ai_1_7/Y fine_freq_track_1/sky130_fd_sc_hs__a22oi_1_23/Y
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_7/a_313_74# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_13/a_706_463#
+ fine_freq_track_1/sky130_fd_sc_hs__a22o_1_25/a_222_392# fine_freq_track_1/sky130_fd_sc_hs__a21oi_1_99/a_117_74#
+ fine_freq_track_1/sky130_fd_sc_hs__inv_4_89/A fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_29/a_300_74#
+ fine_freq_track_1/sky130_fd_sc_hs__inv_4_7/Y fine_freq_track_1/sky130_fd_sc_hs__inv_4_51/Y
+ fine_freq_track_1/sky130_fd_sc_hs__nand2_1_91/A fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_43/a_319_360#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_29/a_494_366# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_43/a_834_355#
+ fine_freq_track_1/sky130_fd_sc_hs__o21a_1_7/A2 fine_freq_track_1/sky130_fd_sc_hs__xor2_1_9/a_194_125#
+ fine_freq_track_1/sky130_fd_sc_hs__nor3_1_15/a_198_368# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_67/a_494_366#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_39/a_1350_392# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_39/a_313_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfstp_2_1/a_781_74# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_13/a_120_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_47/a_922_127# fine_freq_track_1/sky130_fd_sc_hs__o21a_1_75/A1
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_45/a_33_74# fine_freq_track_1/sky130_fd_sc_hs__inv_4_97/A
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_9/a_856_304# fine_freq_track_1/sky130_fd_sc_hs__fa_2_5/B
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_35/a_1678_395# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_9/a_850_127#
+ fine_freq_track_1/sky130_fd_sc_hs__inv_4_99/Y fine_freq_track_1/sky130_fd_sc_hs__inv_4_1/A
+ fine_freq_track_1/sky130_fd_sc_hs__xnor2_1_11/Y fine_freq_track_1/sky130_fd_sc_hs__o21a_1_35/a_376_387#
+ fine_freq_track_1/sky130_fd_sc_hs__a21oi_1_115/a_29_368# fine_freq_track_1/sky130_fd_sc_hs__inv_4_75/Y
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_83/a_313_74# fine_freq_track_1/sky130_fd_sc_hs__inv_4_15/Y
+ fine_freq_track_1/sky130_fd_sc_hs__o31ai_1_1/A3 fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_19/D
+ fine_freq_track_1/sky130_fd_sc_hs__o21a_1_75/a_376_387# fine_freq_track_1/sky130_fd_sc_hs__o21a_1_57/a_83_244#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_69/a_2010_409# fine_freq_track_1/sky130_fd_sc_hs__nand2_2_7/Y
+ fine_freq_track_1/sky130_fd_sc_hs__xnor2_1_7/B fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_11/a_910_118#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_45/a_817_508# fine_freq_track_1/sky130_fd_sc_hs__fa_2_15/a_487_79#
+ fine_freq_track_1/sky130_fd_sc_hs__inv_4_13/Y fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_3/a_1224_74#
+ fine_freq_track_1/sky130_fd_sc_hs__o21a_1_57/X fine_freq_track_1/sky130_fd_sc_hs__dfstp_2_7/a_1356_74#
+ fine_freq_track_1/sky130_fd_sc_hs__nor2b_1_25/a_27_112# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_17/a_2010_409#
+ fine_freq_track_1/sky130_fd_sc_hs__inv_4_107/Y fine_freq_track_1/sky130_fd_sc_hs__nor2b_1_17/a_278_368#
+ fine_freq_track_1/sky130_fd_sc_hs__nand2_1_57/a_117_74# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_41/a_841_401#
+ fine_freq_track_1/sky130_fd_sc_hs__nand2_2_13/Y fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_49/a_124_78#
+ fine_freq_track_1/sky130_fd_sc_hs__a22o_1_1/a_222_392# fine_freq_track_1/sky130_fd_sc_hs__a22oi_1_9/a_339_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_49/a_1934_94# fine_freq_track_1/sky130_fd_sc_hs__o21a_1_1/X
+ fine_freq_track_1/sky130_fd_sc_hs__fa_2_1/SUM fine_freq_track_1/sky130_fd_sc_hs__nand3_1_1/a_233_74#
+ fine_freq_track_1/sky130_fd_sc_hs__o21a_1_49/X fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_43/a_812_138#
+ fine_freq_track_1/sky130_fd_sc_hs__dfxtp_2_3/a_431_508# fine_freq_track_1/sky130_fd_sc_hs__o21a_1_67/A2
+ fine_freq_track_1/sky130_fd_sc_hs__o211ai_1_9/C1 fine_freq_track_1/sky130_fd_sc_hs__a22oi_1_25/a_71_368#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_27/a_1647_81# fine_freq_track_1/sky130_fd_sc_hs__nand2b_1_7/a_27_112#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_57/a_37_78# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_21/a_1827_81#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_61/a_124_78# fine_freq_track_1/sky130_fd_sc_hs__dfxtp_2_1/a_695_459#
+ fine_freq_track_1/sky130_fd_sc_hs__xor2_1_1/X fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_13/a_789_463#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_7/a_2026_424# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_61/a_1827_81#
+ fine_freq_track_1/sky130_fd_sc_hs__a32oi_1_9/a_391_74# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_89/a_1350_392#
+ fine_freq_track_1/sky130_fd_sc_hs__o21a_1_51/a_320_74# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_45/a_498_360#
+ fine_freq_track_1/sky130_fd_sc_hs__a22o_1_15/a_222_392# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_91/a_789_463#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_85/a_1678_395# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_47/a_1627_493#
+ fine_freq_track_1/sky130_fd_sc_hs__conb_1_1/HI fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_3/a_33_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_17/a_1736_119# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_33/a_834_355#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_19/a_494_366# fine_freq_track_1/sky130_fd_sc_hs__o21a_1_31/X
+ fine_freq_track_1/sky130_fd_sc_hs__a32oi_1_5/a_27_368# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_17/a_1266_119#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_37/a_1350_392# fine_freq_track_1/sky130_fd_sc_hs__o21a_1_57/B1
+ fine_freq_track_1/sky130_fd_sc_hs__inv_4_135/A fine_freq_track_1/sky130_fd_sc_hs__inv_4_113/A
+ fine_freq_track_1/sky130_fd_sc_hs__o22ai_1_5/a_27_74# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_27/a_890_138#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_37/a_1465_471# fine_freq_track_1/sky130_fd_sc_hs__inv_4_31/Y
+ fine_freq_track_1/sky130_fd_sc_hs__o211ai_1_1/a_31_74# fine_freq_track_1/sky130_fd_sc_hs__o22ai_1_1/A2
+ fine_freq_track_1/sky130_fd_sc_hs__dfxtp_4_3/a_651_503# fine_freq_track_1/sky130_fd_sc_hs__o21a_1_65/a_376_387#
+ fine_freq_track_1/sky130_fd_sc_hs__o21a_1_77/B1 fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_67/a_2010_409#
+ fine_freq_track_1/sky130_fd_sc_hs__o21a_1_9/A1 fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_5/Q_N
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_17/a_120_74# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_35/a_817_508#
+ fine_freq_track_1/sky130_fd_sc_hs__nor2b_1_33/Y fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_13/a_33_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfxtp_2_9/a_27_74# fine_freq_track_1/sky130_fd_sc_hs__nor2_1_31/a_116_368#
+ fine_freq_track_1/sky130_fd_sc_hs__o21a_1_1/a_83_244# fine_freq_track_1/sky130_fd_sc_hs__o21a_1_21/X
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_45/a_300_74# fine_freq_track_1/sky130_fd_sc_hs__nor2_1_75/B
+ fine_freq_track_1/sky130_fd_sc_hs__nand2_1_91/B fine_freq_track_1/sky130_fd_sc_hs__o21a_1_61/X
+ fine_freq_track_1/sky130_fd_sc_hs__nor2_2_1/a_35_368# fine_freq_track_1/sky130_fd_sc_hs__a21oi_1_119/a_29_368#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_5/a_699_463# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_7/a_300_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_87/a_313_74# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_49/a_1550_119#
+ fine_freq_track_1/sky130_fd_sc_hs__nor2b_1_41/A fine_freq_track_1/sky130_fd_sc_hs__inv_4_5/Y
+ fine_freq_track_1/sky130_fd_sc_hs__fa_2_9/a_484_347# fine_freq_track_1/sky130_fd_sc_hs__a21oi_1_82/a_117_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_11/a_300_74# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_53/a_313_74#
+ fine_freq_track_1/sky130_fd_sc_hs__fa_2_23/a_336_347# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_35/a_1624_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_5/a_922_127# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_39/a_1598_93#
+ fine_freq_track_1/sky130_fd_sc_hs__o21a_1_27/a_83_244# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_33/a_812_138#
+ fine_freq_track_1/sky130_fd_sc_hs__fa_2_3/a_27_79# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_21/a_125_78#
+ fine_freq_track_1/sky130_fd_sc_hs__fa_2_19/a_484_347# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_5/a_1547_508#
+ fine_freq_track_1/sky130_fd_sc_hs__nor2b_1_29/a_27_112# fine_freq_track_1/sky130_fd_sc_hs__nor2b_1_1/a_27_112#
+ fine_freq_track_1/sky130_fd_sc_hs__a22o_1_25/a_230_79# fine_freq_track_1/sky130_fd_sc_hs__nor4_1_3/C
+ fine_freq_track_1/sky130_fd_sc_hs__nor2_2_3/Y fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_5/a_1482_48#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_5/a_2010_409# fine_freq_track_1/sky130_fd_sc_hs__o2bb2ai_1_1/a_114_74#
+ fine_freq_track_1/sky130_fd_sc_hs__fa_2_7/CIN fine_freq_track_1/sky130_fd_sc_hs__o21ai_1_1/Y
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_37/a_38_78# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_51/a_1827_81#
+ fine_freq_track_1/sky130_fd_sc_hs__nand2_4_5/Y fine_freq_track_1/sky130_fd_sc_hs__inv_4_37/Y
+ fine_freq_track_1/sky130_fd_sc_hs__inv_4_17/A fine_freq_track_1/sky130_fd_sc_hs__o21ai_1_5/B1
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_1/a_817_508# fine_freq_track_1/sky130_fd_sc_hs__inv_4_35/A
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_1/a_124_78# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_31/D
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_81/a_789_463# fine_freq_track_1/sky130_fd_sc_hs__fa_2_13/SUM
+ fine_freq_track_1/sky130_fd_sc_hs__a222oi_1_1/Y fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_33/a_706_463#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_23/a_319_360# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_23/a_834_355#
+ fine_freq_track_1/sky130_fd_sc_hs__fa_2_15/a_1119_79# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_25/a_37_78#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_65/a_124_78# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_47/a_494_366#
+ fine_freq_track_1/sky130_fd_sc_hs__dfxtp_4_5/a_27_74# fine_freq_track_1/sky130_fd_sc_hs__dfxtp_4_9/a_1178_124#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_27/a_922_127# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_87/a_494_366#
+ fine_freq_track_1/sky130_fd_sc_hs__o211ai_1_7/a_116_368# fine_freq_track_1/sky130_fd_sc_hs__o21a_1_55/a_320_74#
+ fine_freq_track_1/sky130_fd_sc_hs__a222o_1_1/X fine_freq_track_1/sky130_fd_sc_hs__a32oi_1_1/a_119_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_41/a_1434_74# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_33/a_1678_395#
+ fine_freq_track_1/sky130_fd_sc_hs__o21a_1_21/A1 fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_29/a_1482_48#
+ fine_freq_track_1/sky130_fd_sc_hs__inv_4_127/A fine_freq_track_1/sky130_fd_sc_hs__xnor2_1_1/a_112_119#
+ fine_freq_track_1/sky130_fd_sc_hs__nor2b_1_21/Y fine_freq_track_1/sky130_fd_sc_hs__a22oi_1_5/a_71_368#
+ fine_freq_track_1/sky130_fd_sc_hs__o21a_1_55/a_376_387# fine_freq_track_1/sky130_fd_sc_hs__a21oi_1_55/a_29_368#
+ fine_freq_track_1/sky130_fd_sc_hs__a32oi_1_9/a_27_368# fine_freq_track_1/sky130_fd_sc_hs__nor2_1_61/Y
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_7/a_507_368# fine_freq_track_1/sky130_fd_sc_hs__fa_2_3/a_992_347#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_25/a_817_508# fine_freq_track_1/sky130_fd_sc_hs__dfstp_2_4/a_1566_92#
+ fine_freq_track_1/sky130_fd_sc_hs__nor2_1_95/A fine_freq_track_1/sky130_fd_sc_hs__nor2_1_65/A
+ fine_freq_track_1/sky130_fd_sc_hs__nor2_1_21/a_116_368# fine_freq_track_1/sky130_fd_sc_hs__o21a_1_1/a_376_387#
+ fine_freq_track_1/sky130_fd_sc_hs__nor2_1_3/Y fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_41/a_37_78#
+ fine_freq_track_1/sky130_fd_sc_hs__nor2_1_21/B fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_1/a_498_360#
+ fine_freq_track_1/sky130_fd_sc_hs__nand2_2_9/a_27_74# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_47/a_1550_119#
+ fine_freq_track_1/sky130_fd_sc_hs__sdlclkp_4_1/a_116_395# fine_freq_track_1/sky130_fd_sc_hs__a22oi_1_1/Y
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_15/a_2010_409# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_9/a_706_463#
+ fine_freq_track_1/sky130_fd_sc_hs__a22o_1_21/a_132_392# fine_freq_track_1/sky130_fd_sc_hs__fa_2_13/a_336_347#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_29/a_1598_93# fine_freq_track_1/sky130_fd_sc_hs__nor2b_1_35/a_278_368#
+ fine_freq_track_1/sky130_fd_sc_hs__inv_2_7/A fine_freq_track_1/sky130_fd_sc_hs__xnor2_1_1/a_293_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_23/a_812_138# fine_freq_track_1/sky130_fd_sc_hs__o21a_1_5/a_83_244#
+ fine_freq_track_1/sky130_fd_sc_hs__dfstp_2_5/a_716_456# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_49/a_300_74#
+ fine_freq_track_1/sky130_fd_sc_hs__o21a_1_53/X fine_freq_track_1/sky130_fd_sc_hs__nor2_1_49/B
+ fine_freq_track_1/sky130_fd_sc_hs__and2_2_1/a_31_74# fine_freq_track_1/sky130_fd_sc_hs__inv_4_1/Y
+ fine_freq_track_1/sky130_fd_sc_hs__nand2_1_67/Y fine_freq_track_1/sky130_fd_sc_hs__a21oi_1_85/a_117_74#
+ fine_freq_track_1/sky130_fd_sc_hs__fa_2_15/CIN fine_freq_track_1/sky130_fd_sc_hs__inv_2_9/A
+ fine_freq_track_1/sky130_fd_sc_hs__fa_2_5/a_683_347# fine_freq_track_1/sky130_fd_sc_hs__fa_2_23/CIN
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_33/a_120_74# fine_freq_track_1/sky130_fd_sc_hs__inv_4_51/A
+ fine_freq_track_1/sky130_fd_sc_hs__a21oi_1_51/a_117_74# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_41/a_1827_81#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_47/a_714_127# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_87/a_1350_392#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_85/a_1647_81# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_45/a_1224_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_7/a_789_463# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_25/a_498_360#
+ fine_freq_track_1/sky130_fd_sc_hs__fa_2_13/CIN fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_71/a_789_463#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_83/a_1678_395# fine_freq_track_1/sky130_fd_sc_hs__a222oi_1_1/a_116_392#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_31/Q_N fine_freq_track_1/sky130_fd_sc_hs__dfxtp_2_9/a_644_504#
+ fine_freq_track_1/sky130_fd_sc_hs__a22o_1_27/X fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_13/a_319_360#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_13/a_834_355# fine_freq_track_1/sky130_fd_sc_hs__a21oi_1_101/a_29_368#
+ fine_freq_track_1/sky130_fd_sc_hs__a22o_1_29/a_230_79# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_37/a_494_366#
+ fine_freq_track_1/sky130_fd_sc_hs__nand2_1_111/a_117_74# fine_freq_track_1/sky130_fd_sc_hs__a21oi_1_1/a_117_74#
+ fine_freq_track_1/sky130_fd_sc_hs__sdlclkp_4_1/a_792_48# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_3/a_494_366#
+ fine_freq_track_1/sky130_fd_sc_hs__inv_4_53/A fine_freq_track_1/sky130_fd_sc_hs__o21ai_1_5/a_162_368#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_17/a_922_127# fine_freq_track_1/sky130_fd_sc_hs__o21a_1_43/a_83_244#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_77/a_494_366# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_91/a_834_355#
+ fine_freq_track_1/sky130_fd_sc_hs__dfxtp_2_11/a_206_368# fine_freq_track_1/sky130_fd_sc_hs__nor2_1_91/Y
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_33/D fine_freq_track_1/sky130_fd_sc_hs__a21oi_1_19/Y
+ fine_freq_track_1/sky130_fd_sc_hs__nand2_4_5/a_27_74# fine_freq_track_1/sky130_fd_sc_hs__a22o_1_9/a_132_392#
+ fine_freq_track_1/sky130_fd_sc_hs__dfxtp_2_11/a_1125_508# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_19/a_1482_48#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_35/a_1465_471# fine_freq_track_1/sky130_fd_sc_hs__o21a_1_45/a_376_387#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_69/a_124_78# fine_freq_track_1/sky130_fd_sc_hs__nor2b_1_11/a_27_112#
+ fine_freq_track_1/sky130_fd_sc_hs__nor2b_1_29/Y fine_freq_track_1/sky130_fd_sc_hs__nor2_1_51/B
+ fine_freq_track_1/sky130_fd_sc_hs__nand2_4_7/A fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_85/a_890_138#
+ fine_freq_track_1/sky130_fd_sc_hs__o21a_1_59/a_320_74# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_15/a_817_508#
+ fine_freq_track_1/sky130_fd_sc_hs__a32oi_1_5/a_119_74# fine_freq_track_1/sky130_fd_sc_hs__dfxtp_4_9/a_735_102#
+ fine_freq_track_1/sky130_fd_sc_hs__nor2_1_11/a_116_368# fine_freq_track_1/sky130_fd_sc_hs__o21a_1_71/A2
+ fine_freq_track_1/sky130_fd_sc_hs__o211ai_1_5/a_311_74# fine_freq_track_1/sky130_fd_sc_hs__conb_1_1/LO
+ fine_freq_track_1/sky130_fd_sc_hs__fa_2_21/SUM fine_freq_track_1/sky130_fd_sc_hs__nor2b_1_13/Y
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_19/a_2026_424# fine_freq_track_1/sky130_fd_sc_hs__a21oi_1_59/a_29_368#
+ fine_freq_track_1/sky130_fd_sc_hs__nor2_1_23/Y fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_21/a_38_78#
+ fine_freq_track_1/sky130_fd_sc_hs__a22oi_1_11/a_71_368# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_19/a_1598_93#
+ fine_freq_track_1/sky130_fd_sc_hs__inv_4_67/A fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_13/a_812_138#
+ fine_freq_track_1/sky130_fd_sc_hs__inv_4_3/Y fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_29/D
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_81/a_37_78# fine_freq_track_1/sky130_fd_sc_hs__fa_2_21/a_27_378#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_3/a_1547_508# fine_freq_track_1/sky130_fd_sc_hs__xnor2_1_9/B
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_91/a_812_138# fine_freq_track_1/sky130_fd_sc_hs__fa_2_9/a_1205_79#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_1/a_1647_81# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_5/a_2026_424#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_31/a_1827_81# fine_freq_track_1/sky130_fd_sc_hs__xnor2_1_5/a_293_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_75/a_1647_81# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_21/a_789_463#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_23/a_33_74# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_15/a_498_360#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_39/a_796_463# fine_freq_track_1/sky130_fd_sc_hs__fa_2_1/A
+ fine_freq_track_1/sky130_fd_sc_hs__a22o_1_25/a_52_123# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_61/a_789_463#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_45/a_1627_493# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_15/a_1736_119#
+ fine_freq_track_1/sky130_fd_sc_hs__maj3_1_1/X fine_freq_track_1/sky130_fd_sc_hs__a21oi_1_89/a_117_74#
+ fine_freq_track_1/sky130_fd_sc_hs__xor2_1_11/a_355_368# fine_freq_track_1/sky130_fd_sc_hs__a222oi_1_3/a_461_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_19/a_300_74# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_15/a_1266_119#
+ fine_freq_track_1/sky130_fd_sc_hs__fa_2_19/a_1205_79# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_1/Q
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_35/a_1350_392# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_37/a_120_74#
+ fine_freq_track_1/sky130_fd_sc_hs__inv_4_81/A fine_freq_track_1/sky130_fd_sc_hs__xor2_1_7/a_194_125#
+ fine_freq_track_1/sky130_fd_sc_hs__dfxtp_4_7/a_1178_124# fine_freq_track_1/sky130_fd_sc_hs__nor2_1_15/Y
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_81/a_834_355# fine_freq_track_1/sky130_fd_sc_hs__o21a_1_23/X
+ fine_freq_track_1/sky130_fd_sc_hs__fa_2_21/a_701_79# fine_freq_track_1/sky130_fd_sc_hs__inv_4_97/Y
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_29/a_313_74# fine_freq_track_1/sky130_fd_sc_hs__xnor2_1_7/A
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_31/a_1678_395# fine_freq_track_1/sky130_fd_sc_hs__a21oi_1_23/a_117_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_7/a_856_304# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_29/a_125_78#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_7/a_850_127# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_49/a_1678_395#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_47/a_1482_48# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_3/a_125_78#
+ fine_freq_track_1/sky130_fd_sc_hs__o21ai_1_9/a_27_74# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_31/a_832_118#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_65/a_2010_409# fine_freq_track_1/sky130_fd_sc_hs__a21oi_1_5/a_117_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_1/a_890_138# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_45/a_38_78#
+ fine_freq_track_1/sky130_fd_sc_hs__sdlclkp_4_1/a_324_79# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_5/a_714_127#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_75/a_890_138# fine_freq_track_1/sky130_fd_sc_hs__fa_2_17/CIN
+ fine_freq_track_1/sky130_fd_sc_hs__o21a_1_47/a_83_244# fine_freq_track_1/sky130_fd_sc_hs__a22o_1_1/a_230_79#
+ fine_freq_track_1/sky130_fd_sc_hs__o21a_1_13/a_83_244# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_1/a_1224_74#
+ fine_freq_track_1/sky130_fd_sc_hs__o21a_1_3/a_320_74# fine_freq_track_1/sky130_fd_sc_hs__nor2_1_43/B
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_17/a_2026_424# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_49/a_699_463#
+ fine_freq_track_1/sky130_fd_sc_hs__or3b_2_1/C_N fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_35/a_37_78#
+ fine_freq_track_1/sky130_fd_sc_hs__and2_2_1/a_118_74# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_89/a_699_463#
+ fine_freq_track_1/sky130_fd_sc_hs__nor2b_1_15/a_27_112# fine_freq_track_1/sky130_fd_sc_hs__inv_4_35/Y
+ fine_freq_track_1/sky130_fd_sc_hs__o21a_1_47/X fine_freq_track_1/sky130_fd_sc_hs__a22o_1_11/a_230_79#
+ fine_freq_track_1/sky130_fd_sc_hs__nor3_1_9/a_198_368# fine_freq_track_1/sky130_fd_sc_hs__nand2_1_47/a_117_74#
+ fine_freq_track_1/sky130_fd_sc_hs__inv_4_47/Y fine_freq_track_1/sky130_fd_sc_hs__inv_4_9/A
+ fine_freq_track_1/sky130_fd_sc_hs__nand2_4_11/a_27_74# fine_freq_track_1/sky130_fd_sc_hs__a32oi_1_9/a_119_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_47/a_1934_94# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_43/a_1624_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_49/a_1598_93# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_47/a_33_74#
+ fine_freq_track_1/sky130_fd_sc_hs__sdlclkp_4_1/a_354_105# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_1/a_1547_508#
+ fine_freq_track_1/sky130_fd_sc_hs__nand2_1_91/a_117_74# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_81/a_812_138#
+ fine_freq_track_1/sky130_fd_sc_hs__a32oi_1_7/Y fine_freq_track_1/sky130_fd_sc_hs__a21oi_1_9/Y
+ fine_freq_track_1/sky130_fd_sc_hs__nand2_1_99/A fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_3/a_2010_409#
+ fine_freq_track_1/sky130_fd_sc_hs__a22oi_1_15/a_71_368# fine_freq_track_1/sky130_fd_sc_hs__xnor2_1_1/a_138_385#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_25/a_1647_81# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_27/a_714_127#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_85/a_1350_392# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_7/a_832_118#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_51/a_124_78# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_65/a_1647_81#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_25/a_1224_74# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_7/Q_N
+ fine_freq_track_1/sky130_fd_sc_hs__nor2_1_3/B fine_freq_track_1/sky130_fd_sc_hs__maj3_1_1/a_84_74#
+ fine_freq_track_1/sky130_fd_sc_hs__o21a_1_41/a_320_74# fine_freq_track_1/sky130_fd_sc_hs__inv_4_31/A
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_81/a_1678_395# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_85/D
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_51/a_789_463# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_13/a_1736_119#
+ fine_freq_track_1/sky130_fd_sc_hs__xor2_1_7/a_455_87# fine_freq_track_1/sky130_fd_sc_hs__a22o_1_13/a_222_392#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_13/a_1266_119# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_41/a_706_463#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_7/a_834_355# fine_freq_track_1/sky130_fd_sc_hs__o21a_1_19/A1
+ fine_freq_track_1/sky130_fd_sc_hs__o21a_1_5/A1 fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_33/a_319_360#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_17/a_494_366# fine_freq_track_1/sky130_fd_sc_hs__a21oi_1_41/a_29_368#
+ fine_freq_track_1/sky130_fd_sc_hs__inv_4_111/A fine_freq_track_1/sky130_fd_sc_hs__inv_4_9/Y
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_57/a_494_366# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_71/a_834_355#
+ fine_freq_track_1/sky130_fd_sc_hs__xnor2_1_9/a_293_74# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_37/a_922_127#
+ fine_freq_track_1/sky130_fd_sc_hs__nand2_2_1/A fine_freq_track_1/sky130_fd_sc_hs__a22o_1_29/a_52_123#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_33/a_1465_471# fine_freq_track_1/sky130_fd_sc_hs__o21a_1_25/a_376_387#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_25/a_890_138# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_21/a_832_118#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_63/a_2010_409# fine_freq_track_1/sky130_fd_sc_hs__dfxtp_4_2/a_651_503#
+ fine_freq_track_1/sky130_fd_sc_hs__nor2_1_7/A fine_freq_track_1/sky130_fd_sc_hs__inv_4_121/Y
+ fine_freq_track_1/sky130_fd_sc_hs__o31ai_1_3/B1 fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_65/a_890_138#
+ fine_freq_track_1/sky130_fd_sc_hs__nor2b_1_11/Y fine_freq_track_1/sky130_fd_sc_hs__nor2_1_73/B
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_31/D fine_freq_track_1/sky130_fd_sc_hs__o21a_1_77/X
+ fine_freq_track_1/sky130_fd_sc_hs__a21oi_1_27/a_117_74# fine_freq_track_1/sky130_fd_sc_hs__fa_2_19/a_1094_347#
+ fine_freq_track_1/sky130_fd_sc_hs__nor2_1_89/A fine_freq_track_1/sky130_fd_sc_hs__inv_4_61/Y
+ fine_freq_track_1/sky130_fd_sc_hs__nor2_1_75/Y fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_45/a_1550_119#
+ fine_freq_track_1/sky130_fd_sc_hs__nand4_2_1/D fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_35/a_300_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfxtp_2_9/a_538_429# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_13/a_2010_409#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_77/a_313_74# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_79/a_699_463#
+ fine_freq_track_1/sky130_fd_sc_hs__a21oi_1_71/a_117_74# fine_freq_track_1/sky130_fd_sc_hs__a21oi_1_9/a_117_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfxtp_2_11/a_708_101# fine_freq_track_1/sky130_fd_sc_hs__nor2_1_115/a_116_368#
+ fine_freq_track_1/sky130_fd_sc_hs__dfxtp_2_1/a_27_74# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_9/a_319_360#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_31/a_841_401# fine_freq_track_1/sky130_fd_sc_hs__nor2_1_77/Y
+ fine_freq_track_1/sky130_fd_sc_hs__fa_2_23/a_992_347# fine_freq_track_1/sky130_fd_sc_hs__a22o_1_5/a_230_79#
+ fine_freq_track_1/sky130_fd_sc_hs__nor2b_1_45/a_278_368# fine_freq_track_1/sky130_fd_sc_hs__inv_4_137/Y
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_11/a_313_74# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_7/a_812_138#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_43/a_125_78# fine_freq_track_1/sky130_fd_sc_hs__nor4_1_3/A
+ fine_freq_track_1/sky130_fd_sc_hs__o21a_1_7/a_320_74# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_71/a_812_138#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_75/a_37_78# fine_freq_track_1/sky130_fd_sc_hs__o21a_1_75/X
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_11/a_125_78# fine_freq_track_1/sky130_fd_sc_hs__and2_2_5/a_118_74#
+ fine_freq_track_1/sky130_fd_sc_hs__nor2b_1_19/a_27_112# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_15/a_1647_81#
+ fine_freq_track_1/sky130_fd_sc_hs__o21a_1_29/X fine_freq_track_1/sky130_fd_sc_hs__a22o_1_15/a_230_79#
+ fine_freq_track_1/sky130_fd_sc_hs__fa_2_3/a_1119_79# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_3/a_2026_424#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_11/a_1827_81# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_17/a_714_127#
+ fine_freq_track_1/sky130_fd_sc_hs__o22ai_1_1/A1 fine_freq_track_1/sky130_fd_sc_hs__and2_2_1/X
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_55/a_1647_81# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_15/a_1224_74#
+ fine_freq_track_1/sky130_fd_sc_hs__fa_2_17/B fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_39/a_507_368#
+ fine_freq_track_1/sky130_fd_sc_hs__dfxtp_2_5/D fine_freq_track_1/sky130_fd_sc_hs__nand2b_4_1/a_243_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_41/a_789_463# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_43/a_1627_493#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_35/a_498_360# fine_freq_track_1/sky130_fd_sc_hs__a22oi_1_21/a_159_74#
+ fine_freq_track_1/sky130_fd_sc_hs__nand2_1_95/a_117_74# fine_freq_track_1/sky130_fd_sc_hs__a32oi_1_5/Y
+ fine_freq_track_1/sky130_fd_sc_hs__fa_2_5/A fine_freq_track_1/sky130_fd_sc_hs__a22oi_1_19/a_71_368#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_21/a_834_355# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_33/a_1350_392#
+ fine_freq_track_1/sky130_fd_sc_hs__inv_4_71/Y fine_freq_track_1/sky130_fd_sc_hs__dfxtp_4_5/a_1178_124#
+ fine_freq_track_1/sky130_fd_sc_hs__a21oi_1_105/a_117_74# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_55/a_124_78#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_61/a_834_355# fine_freq_track_1/sky130_fd_sc_hs__sdlclkp_1_1/a_722_492#
+ fine_freq_track_1/sky130_fd_sc_hs__a222oi_1_3/a_369_392# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_5/a_1934_94#
+ fine_freq_track_1/sky130_fd_sc_hs__o211ai_1_5/a_116_368# fine_freq_track_1/sky130_fd_sc_hs__o21a_1_45/a_320_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_7/a_841_401# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_21/a_124_78#
+ fine_freq_track_1/sky130_fd_sc_hs__inv_4_101/A fine_freq_track_1/sky130_fd_sc_hs__a21oi_1_77/a_29_368#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_47/a_1678_395# fine_freq_track_1/sky130_fd_sc_hs__o21a_1_11/a_320_74#
+ fine_freq_track_1/sky130_fd_sc_hs__o21a_1_15/a_376_387# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_27/a_1482_48#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_15/a_890_138# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_11/a_832_118#
+ fine_freq_track_1/sky130_fd_sc_hs__a21oi_1_45/a_29_368# fine_freq_track_1/sky130_fd_sc_hs__inv_4_85/A
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_55/a_890_138# fine_freq_track_1/sky130_fd_sc_hs__a21oi_1_11/a_29_368#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_39/a_38_78# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_9/a_1550_119#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_31/a_33_74# fine_freq_track_1/sky130_fd_sc_hs__fa_2_1/a_336_347#
+ fine_freq_track_1/sky130_fd_sc_hs__dfxtp_4_3/a_696_458# fine_freq_track_1/sky130_fd_sc_hs__dfstp_2_1/a_1566_92#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_39/a_910_118# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_35/D
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_15/a_2026_424# fine_freq_track_1/sky130_fd_sc_hs__nor2b_1_1/a_278_368#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_69/a_699_463# fine_freq_track_1/sky130_fd_sc_hs__a22o_1_1/a_52_123#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_29/a_37_78# fine_freq_track_1/sky130_fd_sc_hs__nor2_1_105/a_116_368#
+ fine_freq_track_1/sky130_fd_sc_hs__dfxtp_4_2/D fine_freq_track_1/sky130_fd_sc_hs__fa_2_1/a_487_79#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_21/a_841_401# fine_freq_track_1/sky130_fd_sc_hs__o21a_1_51/X
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_23/a_1624_74# fine_freq_track_1/sky130_fd_sc_hs__fa_2_11/a_336_347#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_27/a_1934_94# fine_freq_track_1/sky130_fd_sc_hs__fa_2_13/a_992_347#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_15/Q_N fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_11/D
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_21/a_812_138# fine_freq_track_1/sky130_fd_sc_hs__a22o_1_11/a_52_123#
+ fine_freq_track_1/sky130_fd_sc_hs__dfstp_2_4/a_716_456# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_61/a_812_138#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_1/a_2010_409# fine_freq_track_1/sky130_fd_sc_hs__a21oi_1_75/a_117_74#
+ fine_freq_track_1/sky130_fd_sc_hs__o22ai_1_9/a_340_368# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_1/a_2026_424#
+ fine_freq_track_1/sky130_fd_sc_hs__dfstp_2_4/a_27_74# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_83/a_1350_392#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_47/a_313_74# fine_freq_track_1/sky130_fd_sc_hs__nand2_1_85/Y
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_45/a_1647_81# fine_freq_track_1/sky130_fd_sc_hs__a222o_1_1/a_27_390#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_23/a_120_74# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_29/a_507_368#
+ fine_freq_track_1/sky130_fd_sc_hs__nor2b_1_3/Y fine_freq_track_1/sky130_fd_sc_hs__a22o_1_9/a_230_79#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_31/a_789_463# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_47/a_125_78#
+ fine_freq_track_1/sky130_fd_sc_hs__xor2_1_3/a_355_368# fine_freq_track_1/sky130_fd_sc_hs__inv_4_109/Y
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_11/a_1736_119# fine_freq_track_1/sky130_fd_sc_hs__a21oi_1_123/a_29_368#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_11/a_1266_119# fine_freq_track_1/sky130_fd_sc_hs__dfxtp_2_7/a_644_504#
+ fine_freq_track_1/sky130_fd_sc_hs__or2_1_3/a_63_368# fine_freq_track_1/sky130_fd_sc_hs__a22o_1_19/a_230_79#
+ fine_freq_track_1/sky130_fd_sc_hs__fa_2_15/a_683_347# fine_freq_track_1/sky130_fd_sc_hs__a31oi_1_1/a_145_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_51/a_834_355# fine_freq_track_1/sky130_fd_sc_hs__maj3_1_3/X
+ fine_freq_track_1/sky130_fd_sc_hs__o21a_1_33/a_83_244# fine_freq_track_1/sky130_fd_sc_hs__dfstp_2_7/D
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_31/a_1434_74# fine_freq_track_1/sky130_fd_sc_hs__o21a_1_3/X
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_31/a_1465_471# fine_freq_track_1/sky130_fd_sc_hs__a22oi_1_25/a_159_74#
+ fine_freq_track_1/sky130_fd_sc_hs__nand2b_1_3/Y fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_17/a_1482_48#
+ fine_freq_track_1/sky130_fd_sc_hs__nand3b_2_1/a_403_54# fine_freq_track_1/sky130_fd_sc_hs__o22ai_1_3/Y
+ fine_freq_track_1/sky130_fd_sc_hs__a21oi_1_109/a_117_74# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_45/a_890_138#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_59/a_124_78# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_7/a_1550_119#
+ fine_freq_track_1/sky130_fd_sc_hs__nand2_1_33/a_117_74# fine_freq_track_1/sky130_fd_sc_hs__o21a_1_49/a_320_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_13/a_817_508# fine_freq_track_1/sky130_fd_sc_hs__fa_2_17/a_1094_347#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_25/a_124_78# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_43/a_1550_119#
+ fine_freq_track_1/sky130_fd_sc_hs__nor3_1_3/a_114_368# fine_freq_track_1/sky130_fd_sc_hs__xnor2_1_11/a_293_74#
+ fine_freq_track_1/sky130_fd_sc_hs__o22ai_1_9/A1 fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_11/a_2010_409#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_59/a_699_463# fine_freq_track_1/sky130_fd_sc_hs__nor2_1_99/a_116_368#
+ fine_freq_track_1/sky130_fd_sc_hs__nor2_1_59/A fine_freq_track_1/sky130_fd_sc_hs__a21oi_1_121/a_117_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_11/a_841_401# fine_freq_track_1/sky130_fd_sc_hs__a22o_1_11/a_132_392#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_17/a_1934_94# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_13/a_1624_74#
+ fine_freq_track_1/sky130_fd_sc_hs__clkbuf_2_1/a_43_192# fine_freq_track_1/sky130_fd_sc_hs__nor2b_1_25/a_278_368#
+ fine_freq_track_1/sky130_fd_sc_hs__o21a_1_15/X fine_freq_track_1/sky130_fd_sc_hs__a21oi_1_93/a_29_368#
+ fine_freq_track_1/sky130_fd_sc_hs__nand2_4_7/a_27_74# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_51/a_812_138#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_39/a_856_304# fine_freq_track_1/sky130_fd_sc_hs__nor3_1_1/C
+ fine_freq_track_1/sky130_fd_sc_hs__nor2_1_9/B fine_freq_track_1/sky130_fd_sc_hs__maj3_1_3/a_226_384#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_7/a_1434_74# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_39/a_850_127#
+ fine_freq_track_1/sky130_fd_sc_hs__a22o_1_5/a_52_123# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_69/a_37_78#
+ fine_freq_track_1/sky130_fd_sc_hs__fa_2_5/a_487_79# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_35/a_1647_81#
+ fine_freq_track_1/sky130_fd_sc_hs__nor2_1_83/Y fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_19/a_507_368#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_5/a_1827_81# fine_freq_track_1/sky130_fd_sc_hs__nand4_1_1/Y
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_37/a_714_127# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_73/a_1647_81#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_35/a_1224_74# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_41/a_1627_493#
+ fine_freq_track_1/sky130_fd_sc_hs__a22o_1_15/a_52_123# fine_freq_track_1/sky130_fd_sc_hs__o22ai_1_9/a_142_368#
+ fine_freq_track_1/sky130_fd_sc_hs__dfstp_2_5/a_1278_74# fine_freq_track_1/sky130_fd_sc_hs__a22o_1_23/a_222_392#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_29/a_1736_119# fine_freq_track_1/sky130_fd_sc_hs__inv_4_95/Y
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_31/a_1350_392# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_23/a_38_78#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_41/a_319_360# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_27/a_494_366#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_41/a_834_355# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_29/a_1266_119#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_49/a_1350_392# fine_freq_track_1/sky130_fd_sc_hs__a21oi_1_82/Y
+ fine_freq_track_1/sky130_fd_sc_hs__nor3_1_13/a_198_368# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_19/a_313_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_21/a_1434_74# fine_freq_track_1/sky130_fd_sc_hs__a21oi_1_13/a_117_74#
+ fine_freq_track_1/sky130_fd_sc_hs__o2bb2ai_1_1/a_131_383# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_19/a_125_78#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_13/a_37_78# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_61/a_2010_409#
+ fine_freq_track_1/sky130_fd_sc_hs__nand4_1_1/a_259_74# fine_freq_track_1/sky130_fd_sc_hs__dfxtp_2_5/a_206_368#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_35/a_890_138# fine_freq_track_1/sky130_fd_sc_hs__a31oi_1_1/A2
+ fine_freq_track_1/sky130_fd_sc_hs__o21a_1_73/a_376_387# fine_freq_track_1/sky130_fd_sc_hs__nor4_1_3/D
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_73/a_890_138# fine_freq_track_1/sky130_fd_sc_hs__nor3_1_9/A
+ fine_freq_track_1/sky130_fd_sc_hs__nor2b_1_1/Y fine_freq_track_1/sky130_fd_sc_hs__dfsbp_2_1/Q
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_43/a_817_508# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_41/a_1550_119#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_13/a_2026_424# fine_freq_track_1/sky130_fd_sc_hs__nor2_1_41/B
+ fine_freq_track_1/sky130_fd_sc_hs__o21a_1_45/X fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_5/a_796_463#
+ fine_freq_track_1/sky130_fd_sc_hs__nor2_1_89/a_116_368# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_29/a_2010_409#
+ fine_freq_track_1/sky130_fd_sc_hs__nor2b_1_15/a_278_368# fine_freq_track_1/sky130_fd_sc_hs__nand2_1_37/a_117_74#
+ fine_freq_track_1/sky130_fd_sc_hs__a22oi_1_23/a_339_74# fine_freq_track_1/sky130_fd_sc_hs__dfsbp_2_1/a_1501_92#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_47/a_1598_93# fine_freq_track_1/sky130_fd_sc_hs__dfsbp_2_1/a_1521_508#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_91/a_1627_493# fine_freq_track_1/sky130_fd_sc_hs__a22oi_1_5/a_159_74#
+ fine_freq_track_1/sky130_fd_sc_hs__xnor2_1_15/a_293_74# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_41/a_812_138#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_29/a_856_304# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_29/a_850_127#
+ fine_freq_track_1/sky130_fd_sc_hs__dfxtp_2_1/a_431_508# fine_freq_track_1/sky130_fd_sc_hs__nand2_1_81/a_117_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_73/a_124_78# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_81/a_1350_392#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_83/D fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_41/a_124_78#
+ fine_freq_track_1/sky130_fd_sc_hs__o21a_1_13/A1 fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_63/a_1647_81#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_11/a_789_463# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_49/a_507_368#
+ fine_freq_track_1/sky130_fd_sc_hs__a21oi_1_97/a_29_368# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_29/a_796_463#
+ fine_freq_track_1/sky130_fd_sc_hs__o21a_1_31/a_320_74# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_43/a_498_360#
+ fine_freq_track_1/sky130_fd_sc_hs__dfstp_2_5/a_398_74# fine_freq_track_1/sky130_fd_sc_hs__a2bb2oi_1_1/Y
+ fine_freq_track_1/sky130_fd_sc_hs__fa_2_15/a_27_378# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_59/a_1627_493#
+ fine_freq_track_1/sky130_fd_sc_hs__a22o_1_9/a_52_123# fine_freq_track_1/sky130_fd_sc_hs__dfxtp_4_3/a_1178_124#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_37/a_37_78# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_31/a_834_355#
+ fine_freq_track_1/sky130_fd_sc_hs__fa_2_9/a_487_79# fine_freq_track_1/sky130_fd_sc_hs__a21oi_1_31/a_29_368#
+ fine_freq_track_1/sky130_fd_sc_hs__fa_2_23/a_1119_79# fine_freq_track_1/sky130_fd_sc_hs__o211ai_1_5/Y
+ fine_freq_track_1/sky130_fd_sc_hs__nand2_1_23/Y fine_freq_track_1/sky130_fd_sc_hs__nand2_4_15/a_27_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_19/a_1547_508# fine_freq_track_1/sky130_fd_sc_hs__nor2_1_13/Y
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_11/a_1434_74# fine_freq_track_1/sky130_fd_sc_hs__a22o_1_19/a_52_123#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_45/a_1678_395# fine_freq_track_1/sky130_fd_sc_hs__o21ai_1_9/Y
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_37/a_1482_48# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_47/a_1465_471#
+ fine_freq_track_1/sky130_fd_sc_hs__o21a_1_63/a_376_387# fine_freq_track_1/sky130_fd_sc_hs__nor2_2_1/A
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_79/a_2010_409# fine_freq_track_1/sky130_fd_sc_hs__a21oi_1_49/a_117_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_63/a_890_138# fine_freq_track_1/sky130_fd_sc_hs__dfxtp_4_3/a_544_485#
+ fine_freq_track_1/sky130_fd_sc_hs__fa_2_15/a_701_79# fine_freq_track_1/sky130_fd_sc_hs__a21oi_1_17/a_117_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_3/a_313_74# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_33/a_817_508#
+ fine_freq_track_1/sky130_fd_sc_hs__nor2_1_79/a_116_368# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_39/a_699_463#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_25/a_300_74# fine_freq_track_1/sky130_fd_sc_hs__dfxtp_2_7/a_538_429#
+ fine_freq_track_1/sky130_fd_sc_hs__nand4_1_5/a_259_74# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_41/a_120_74#
+ fine_freq_track_1/sky130_fd_sc_hs__fa_2_7/a_484_347# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_5/D
+ fine_freq_track_1/sky130_fd_sc_hs__a21oi_1_61/a_117_74# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_5/a_120_74#
+ fine_freq_track_1/sky130_fd_sc_hs__xnor2_1_9/a_376_368# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_37/a_1934_94#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_33/a_1624_74# fine_freq_track_1/sky130_fd_sc_hs__inv_2_1/Y
+ fine_freq_track_1/sky130_fd_sc_hs__fa_2_21/a_336_347# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_3/a_922_127#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_19/a_856_304# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_31/a_812_138#
+ fine_freq_track_1/sky130_fd_sc_hs__a32oi_1_5/A1 fine_freq_track_1/sky130_fd_sc_hs__o21a_1_37/X
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_19/a_850_127# fine_freq_track_1/sky130_fd_sc_hs__nand2_1_121/a_117_74#
+ fine_freq_track_1/sky130_fd_sc_hs__fa_2_17/a_484_347# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_3/a_1482_48#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_53/a_1647_81# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_19/a_796_463#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_45/Q_N fine_freq_track_1/sky130_fd_sc_hs__o22ai_1_1/a_27_74#
+ fine_freq_track_1/sky130_fd_sc_hs__a22oi_1_11/a_159_74# fine_freq_track_1/sky130_fd_sc_hs__dfxtp_2_9/a_1125_508#
+ fine_freq_track_1/sky130_fd_sc_hs__xor2_1_5/a_158_392# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_27/a_1736_119#
+ fine_freq_track_1/sky130_fd_sc_hs__nand2_1_85/a_117_74# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_37/Q_N
+ fine_freq_track_1/sky130_fd_sc_hs__nand3b_2_1/a_206_74# fine_freq_track_1/sky130_fd_sc_hs__dfxtp_4_2/a_1178_124#
+ fine_freq_track_1/sky130_fd_sc_hs__conb_1_1/a_21_290# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_9/a_33_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_31/a_706_463# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_27/a_1266_119#
+ fine_freq_track_1/sky130_fd_sc_hs__fa_2_13/a_1119_79# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_27/Q_N
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_47/a_1350_392# fine_freq_track_1/sky130_fd_sc_hs__sdlclkp_4_1/a_119_143#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_17/a_38_78# fine_freq_track_1/sky130_fd_sc_hs__nor2_1_11/Y
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_45/a_124_78# fine_freq_track_1/sky130_fd_sc_hs__dfxtp_2_5/a_27_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_5/a_1598_93# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_19/Q_N
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_85/a_494_366# fine_freq_track_1/sky130_fd_sc_hs__o31ai_1_5/Y
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_9/a_1624_74# fine_freq_track_1/sky130_fd_sc_hs__dfstp_2_7/a_398_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfxtp_4_9/a_206_368# fine_freq_track_1/sky130_fd_sc_hs__o21a_1_13/a_376_387#
+ fine_freq_track_1/sky130_fd_sc_hs__sdlclkp_4_1/a_1289_368# fine_freq_track_1/sky130_fd_sc_hs__nand2_2_3/Y
+ fine_freq_track_1/sky130_fd_sc_hs__o21a_1_53/a_376_387# fine_freq_track_1/sky130_fd_sc_hs__o211ai_1_7/a_31_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_5/a_1550_119# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_53/a_890_138#
+ fine_freq_track_1/sky130_fd_sc_hs__fa_2_15/a_1094_347# fine_freq_track_1/sky130_fd_sc_hs__fa_2_23/a_27_79#
+ fine_freq_track_1/sky130_fd_sc_hs__fa_2_1/a_992_347# fine_freq_track_1/sky130_fd_sc_hs__dfxtp_4_2/a_696_458#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_23/a_817_508# fine_freq_track_1/sky130_fd_sc_hs__o21a_1_9/a_376_387#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_19/a_33_74# fine_freq_track_1/sky130_fd_sc_hs__o31ai_1_5/a_114_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_29/a_699_463# fine_freq_track_1/sky130_fd_sc_hs__nor2_1_69/a_116_368#
+ fine_freq_track_1/sky130_fd_sc_hs__inv_4_73/Y fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_27/a_2010_409#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_33/a_38_78# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_67/a_699_463#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_15/D fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_7/a_706_463#
+ fine_freq_track_1/sky130_fd_sc_hs__fa_2_11/a_992_347# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_27/a_1598_93#
+ fine_freq_track_1/sky130_fd_sc_hs__o21ai_1_1/B1 fine_freq_track_1/sky130_fd_sc_hs__dfxtp_2_5/a_708_101#
+ fine_freq_track_1/sky130_fd_sc_hs__fa_2_9/a_27_79# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_21/a_37_78#
+ fine_freq_track_1/sky130_fd_sc_hs__dfstp_2_1/a_716_456# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_49/a_856_304#
+ fine_freq_track_1/sky130_fd_sc_hs__dfxtp_4_2/a_27_74# fine_freq_track_1/sky130_fd_sc_hs__dfxtp_4_7/Q
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_49/a_850_127# fine_freq_track_1/sky130_fd_sc_hs__a21oi_1_65/a_117_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_9/a_120_74# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_37/a_313_74#
+ fine_freq_track_1/sky130_fd_sc_hs__fa_2_3/a_683_347# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_49/a_1827_81#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_35/a_33_74# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_83/a_1647_81#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_43/a_1224_74# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_89/a_1827_81#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_5/a_789_463# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_23/a_498_360#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_47/a_796_463# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_57/a_1627_493#
+ fine_freq_track_1/sky130_fd_sc_hs__a21oi_1_113/a_29_368# fine_freq_track_1/sky130_fd_sc_hs__dfxtp_2_7/a_1125_508#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_3/a_300_74# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_5/a_910_118#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_21/a_706_463# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_11/a_834_355#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_17/a_1547_508# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_1/a_494_366#
+ fine_freq_track_1/sky130_fd_sc_hs__nand2_2_15/a_27_74# fine_freq_track_1/sky130_fd_sc_hs__o21ai_1_3/a_162_368#
+ fine_freq_track_1/sky130_fd_sc_hs__o21a_1_23/a_83_244# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_75/a_494_366#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_43/a_1678_395# fine_freq_track_1/sky130_fd_sc_hs__fa_2_9/A
+ fine_freq_track_1/sky130_fd_sc_hs__a222oi_1_3/a_697_74# fine_freq_track_1/sky130_fd_sc_hs__a22oi_1_15/a_159_74#
+ fine_freq_track_1/sky130_fd_sc_hs__a22o_1_7/a_132_392# fine_freq_track_1/sky130_fd_sc_hs__nand2_1_89/a_117_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_45/a_1465_471# fine_freq_track_1/sky130_fd_sc_hs__dfxtp_4_9/a_437_503#
+ fine_freq_track_1/sky130_fd_sc_hs__o21a_1_43/a_376_387# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_77/a_2010_409#
+ fine_freq_track_1/sky130_fd_sc_hs__xnor2_1_1/Y fine_freq_track_1/sky130_fd_sc_hs__nor2_1_95/B
+ fine_freq_track_1/sky130_fd_sc_hs__nand2b_1_3/a_269_74# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_83/a_890_138#
+ fine_freq_track_1/sky130_fd_sc_hs__nand2_1_23/a_117_74# fine_freq_track_1/sky130_fd_sc_hs__o21a_1_39/a_320_74#
+ fine_freq_track_1/sky130_fd_sc_hs__fa_2_7/B fine_freq_track_1/sky130_fd_sc_hs__nor2_1_47/Y
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_11/a_2026_424# fine_freq_track_1/sky130_fd_sc_hs__dfsbp_2_1/a_1531_118#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_29/a_910_118# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_15/a_124_78#
+ fine_freq_track_1/sky130_fd_sc_hs__nor3_1_3/B fine_freq_track_1/sky130_fd_sc_hs__dfxtp_4_7/a_735_102#
+ fine_freq_track_1/sky130_fd_sc_hs__nor2_1_91/B fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_19/a_699_463#
+ fine_freq_track_1/sky130_fd_sc_hs__nor2_1_59/a_116_368# fine_freq_track_1/sky130_fd_sc_hs__fa_2_9/a_1094_347#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_25/a_2010_409# fine_freq_track_1/sky130_fd_sc_hs__a21oi_1_39/a_29_368#
+ fine_freq_track_1/sky130_fd_sc_hs__a21oi_1_111/a_117_74# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_25/D
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_17/a_1598_93# fine_freq_track_1/sky130_fd_sc_hs__fa_2_1/B
+ fine_freq_track_1/sky130_fd_sc_hs__dfxtp_4_9/a_1034_424# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_11/a_812_138#
+ fine_freq_track_1/sky130_fd_sc_hs__a22oi_1_13/Y fine_freq_track_1/sky130_fd_sc_hs__inv_4_83/A
+ fine_freq_track_1/sky130_fd_sc_hs__nand4_1_3/a_181_74# fine_freq_track_1/sky130_fd_sc_hs__maj3_1_1/a_226_384#
+ fine_freq_track_1/sky130_fd_sc_hs__a22oi_1_1/a_71_368# fine_freq_track_1/sky130_fd_sc_hs__fa_2_7/a_1205_79#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_9/a_1647_81# fine_freq_track_1/sky130_fd_sc_hs__nand2_4_1/a_27_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_79/a_1827_81# fine_freq_track_1/sky130_fd_sc_hs__o21a_1_13/X
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_13/a_498_360# fine_freq_track_1/sky130_fd_sc_hs__sdlclkp_1_1/a_1238_94#
+ fine_freq_track_1/sky130_fd_sc_hs__nor2_1_9/a_116_368# fine_freq_track_1/sky130_fd_sc_hs__dfstp_2_4/a_1278_74#
+ fine_freq_track_1/sky130_fd_sc_hs__inv_4_5/A fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_11/a_706_463#
+ fine_freq_track_1/sky130_fd_sc_hs__a22o_1_21/a_222_392# fine_freq_track_1/sky130_fd_sc_hs__a21oi_1_69/a_117_74#
+ fine_freq_track_1/sky130_fd_sc_hs__nor2_1_43/Y fine_freq_track_1/sky130_fd_sc_hs__fa_2_17/a_1205_79#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_25/a_494_366# fine_freq_track_1/sky130_fd_sc_hs__a211oi_4_1/a_901_368#
+ fine_freq_track_1/sky130_fd_sc_hs__a21oi_1_35/a_117_74# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_65/a_494_366#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_45/a_922_127# fine_freq_track_1/sky130_fd_sc_hs__nand4_2_1/a_515_74#
+ fine_freq_track_1/sky130_fd_sc_hs__nor3_1_7/A fine_freq_track_1/sky130_fd_sc_hs__o21a_1_33/a_376_387#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_45/a_1482_48# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_39/a_832_118#
+ fine_freq_track_1/sky130_fd_sc_hs__fa_2_21/B fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_3/a_1550_119#
+ fine_freq_track_1/sky130_fd_sc_hs__dfxtp_2_3/a_206_368# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_9/a_890_138#
+ fine_freq_track_1/sky130_fd_sc_hs__fa_2_13/a_1094_347# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_3/a_714_127#
+ fine_freq_track_1/sky130_fd_sc_hs__o21a_1_43/X fine_freq_track_1/sky130_fd_sc_hs__fa_2_17/a_487_79#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_19/a_910_118# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_41/a_817_508#
+ fine_freq_track_1/sky130_fd_sc_hs__a22oi_1_19/a_159_74# fine_freq_track_1/sky130_fd_sc_hs__nor2_1_49/a_116_368#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_29/a_2026_424# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_47/a_699_463#
+ fine_freq_track_1/sky130_fd_sc_hs__o21a_1_71/a_83_244# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_5/D
+ fine_freq_track_1/sky130_fd_sc_hs__nand2b_1_7/a_269_74# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_87/a_699_463#
+ fine_freq_track_1/sky130_fd_sc_hs__nor2_1_123/a_116_368# fine_freq_track_1/sky130_fd_sc_hs__a222oi_1_3/a_119_74#
+ fine_freq_track_1/sky130_fd_sc_hs__nor2b_1_13/a_278_368# fine_freq_track_1/sky130_fd_sc_hs__nand2_1_27/a_117_74#
+ fine_freq_track_1/sky130_fd_sc_hs__a22oi_1_13/a_339_74# fine_freq_track_1/sky130_fd_sc_hs__nor3_1_7/a_198_368#
+ fine_freq_track_1/sky130_fd_sc_hs__a22o_1_9/a_222_392# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_41/a_1624_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfstp_2_7/a_1521_508# fine_freq_track_1/sky130_fd_sc_hs__o31ai_1_7/a_119_368#
+ fine_freq_track_1/sky130_fd_sc_hs__inv_4_19/Y fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_87/a_37_78#
+ fine_freq_track_1/sky130_fd_sc_hs__nand2_1_71/a_117_74# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_15/a_37_78#
+ fine_freq_track_1/sky130_fd_sc_hs__a21oi_1_115/a_117_74# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_63/a_124_78#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_31/a_124_78# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_23/a_1224_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_69/a_1827_81# fine_freq_track_1/sky130_fd_sc_hs__o211ai_1_1/a_311_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_47/a_507_368# fine_freq_track_1/sky130_fd_sc_hs__a21oi_1_87/a_29_368#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_27/a_796_463# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_55/a_1627_493#
+ fine_freq_track_1/sky130_fd_sc_hs__o21a_1_21/a_320_74# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_25/a_1736_119#
+ fine_freq_track_1/sky130_fd_sc_hs__o21ai_1_5/a_27_74# fine_freq_track_1/sky130_fd_sc_hs__dfstp_2_7/a_767_384#
+ fine_freq_track_1/sky130_fd_sc_hs__a21oi_1_53/a_29_368# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_25/a_1266_119#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_41/a_38_78# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_45/a_1350_392#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_31/a_319_360# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_15/a_494_366#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_5/a_834_355# fine_freq_track_1/sky130_fd_sc_hs__a21oi_1_21/a_29_368#
+ fine_freq_track_1/sky130_fd_sc_hs__inv_4_93/A fine_freq_track_1/sky130_fd_sc_hs__o21ai_1_7/Y
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_55/a_494_366# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_41/a_1678_395#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_35/a_922_127# fine_freq_track_1/sky130_fd_sc_hs__o21a_1_73/X
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_31/a_37_78# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_43/a_1465_471#
+ fine_freq_track_1/sky130_fd_sc_hs__a21oi_1_3/a_29_368# fine_freq_track_1/sky130_fd_sc_hs__o21a_1_23/a_376_387#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_75/a_2010_409# fine_freq_track_1/sky130_fd_sc_hs__fa_2_19/a_1202_368#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_1/a_1550_119# fine_freq_track_1/sky130_fd_sc_hs__fa_2_11/a_1094_347#
+ fine_freq_track_1/sky130_fd_sc_hs__dfxtp_4_2/a_544_485# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_47/a_300_74#
+ fine_freq_track_1/sky130_fd_sc_hs__nor2_2_3/a_35_368# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_31/a_817_508#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_47/a_910_118# fine_freq_track_1/sky130_fd_sc_hs__nor2_1_39/a_116_368#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_27/a_2026_424# fine_freq_track_1/sky130_fd_sc_hs__o21a_1_5/B1
+ fine_freq_track_1/sky130_fd_sc_hs__fa_2_7/a_1094_347# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_39/Q_N
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_37/a_699_463# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_15/a_300_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_3/a_699_463# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_57/a_313_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_77/a_699_463# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_31/a_120_74#
+ fine_freq_track_1/sky130_fd_sc_hs__nor2_1_113/a_116_368# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_39/a_841_401#
+ fine_freq_track_1/sky130_fd_sc_hs__a222o_1_1/a_386_74# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_7/a_319_360#
+ fine_freq_track_1/sky130_fd_sc_hs__dfxtp_4_7/a_1034_424# fine_freq_track_1/sky130_fd_sc_hs__fa_2_21/a_992_347#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_1/a_922_127# fine_freq_track_1/sky130_fd_sc_hs__nor2b_1_43/a_278_368#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_37/a_1598_93# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_23/a_125_78#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_5/a_812_138# fine_freq_track_1/sky130_fd_sc_hs__nor2b_1_5/a_27_112#
+ fine_freq_track_1/sky130_fd_sc_hs__o21a_1_75/a_83_244# fine_freq_track_1/sky130_fd_sc_hs__inv_4_115/Y
+ fine_freq_track_1/sky130_fd_sc_hs__a211oi_1_3/a_71_368# fine_freq_track_1/sky130_fd_sc_hs__nand2_1_51/Y
+ fine_freq_track_1/sky130_fd_sc_hs__o21a_1_69/A2 fine_freq_track_1/sky130_fd_sc_hs__fa_2_1/a_1119_79#
+ fine_freq_track_1/sky130_fd_sc_hs__dfstp_2_5/D fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_1/a_1482_48#
+ fine_freq_track_1/sky130_fd_sc_hs__a22oi_1_17/a_339_74# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_13/a_1224_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_59/a_1827_81# fine_freq_track_1/sky130_fd_sc_hs__dfxtp_2_11/a_644_504#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_17/a_796_463# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_91/a_1678_395#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_53/a_1627_493# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_49/a_789_463#
+ fine_freq_track_1/sky130_fd_sc_hs__dfxtp_2_5/a_1125_508# fine_freq_track_1/sky130_fd_sc_hs__nor2b_1_43/a_27_112#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_33/a_498_360# fine_freq_track_1/sky130_fd_sc_hs__nand2b_4_1/a_31_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_89/a_789_463# fine_freq_track_1/sky130_fd_sc_hs__dfsbp_2_1/a_757_401#
+ fine_freq_track_1/sky130_fd_sc_hs__nand2_1_75/a_117_74# fine_freq_track_1/sky130_fd_sc_hs__a21oi_1_119/a_117_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_67/a_124_78# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_21/a_319_360#
+ fine_freq_track_1/sky130_fd_sc_hs__fa_2_11/a_1119_79# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_15/a_1547_508#
+ fine_freq_track_1/sky130_fd_sc_hs__dfstp_2_5/a_225_74# fine_freq_track_1/sky130_fd_sc_hs__nand2_1_41/a_117_74#
+ fine_freq_track_1/sky130_fd_sc_hs__fa_2_23/a_683_347# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_45/a_494_366#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_35/a_124_78# fine_freq_track_1/sky130_fd_sc_hs__a222oi_1_1/a_369_392#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_3/a_1934_94# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_25/a_922_127#
+ fine_freq_track_1/sky130_fd_sc_hs__o21a_1_25/a_320_74# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_1/a_33_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_59/a_1678_395# fine_freq_track_1/sky130_fd_sc_hs__a22oi_1_9/a_71_368#
+ fine_freq_track_1/sky130_fd_sc_hs__o21a_1_67/X fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_7/a_37_78#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_11/a_38_78# fine_freq_track_1/sky130_fd_sc_hs__xnor2_1_9/a_112_119#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_25/a_1482_48# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_73/a_2010_409#
+ fine_freq_track_1/sky130_fd_sc_hs__inv_4_7/A fine_freq_track_1/sky130_fd_sc_hs__nand2_1_3/a_117_74#
+ fine_freq_track_1/sky130_fd_sc_hs__a21oi_1_25/a_29_368# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_5/a_507_368#
+ fine_freq_track_1/sky130_fd_sc_hs__xnor2_1_9/A fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_21/a_817_508#
+ fine_freq_track_1/sky130_fd_sc_hs__nor2_1_29/a_116_368# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_71/a_37_78#
+ fine_freq_track_1/sky130_fd_sc_hs__xor2_1_3/a_455_87# fine_freq_track_1/sky130_fd_sc_hs__a21oi_1_7/a_29_368#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_17/D fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_23/a_2010_409#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_9/a_498_360# fine_freq_track_1/sky130_fd_sc_hs__nand2_2_9/B
+ fine_freq_track_1/sky130_fd_sc_hs__nor2_1_103/a_116_368# fine_freq_track_1/sky130_fd_sc_hs__dfxtp_2_7/a_27_74#
+ fine_freq_track_1/sky130_fd_sc_hs__nor2b_1_33/a_278_368# fine_freq_track_1/sky130_fd_sc_hs__sdlclkp_1_1/a_709_54#
+ fine_freq_track_1/sky130_fd_sc_hs__inv_4_95/A fine_freq_track_1/sky130_fd_sc_hs__nand2_2_11/Y
+ fine_freq_track_1/sky130_fd_sc_hs__dfxtp_2_3/a_708_101# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_47/a_856_304#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_47/a_850_127# fine_freq_track_1/sky130_fd_sc_hs__a21oi_1_55/a_117_74#
+ fine_freq_track_1/sky130_fd_sc_hs__inv_4_29/Y fine_freq_track_1/sky130_fd_sc_hs__o22ai_1_7/a_340_368#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_43/a_1647_81# fine_freq_track_1/sky130_fd_sc_hs__a21oi_1_15/Y
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_27/a_507_368# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_45/a_714_127#
+ fine_freq_track_1/sky130_fd_sc_hs__dfxtp_2_3/a_1125_508# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_23/a_1736_119#
+ fine_freq_track_1/sky130_fd_sc_hs__a31oi_1_1/a_136_368# fine_freq_track_1/sky130_fd_sc_hs__o21a_1_77/A2
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_27/a_125_78# fine_freq_track_1/sky130_fd_sc_hs__xor2_1_1/a_355_368#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_79/a_789_463# fine_freq_track_1/sky130_fd_sc_hs__nor2b_1_9/a_27_112#
+ fine_freq_track_1/sky130_fd_sc_hs__a21oi_1_103/a_29_368# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_1/a_125_78#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_23/a_1266_119# fine_freq_track_1/sky130_fd_sc_hs__nand2_1_115/a_117_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_43/a_1350_392# fine_freq_track_1/sky130_fd_sc_hs__nor2_1_29/B
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_11/a_319_360# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_13/a_1547_508#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_9/a_38_78# fine_freq_track_1/sky130_fd_sc_hs__nand2_2_3/B
+ fine_freq_track_1/sky130_fd_sc_hs__nor2_1_19/B fine_freq_track_1/sky130_fd_sc_hs__fa_2_13/a_683_347#
+ fine_freq_track_1/sky130_fd_sc_hs__xor2_1_11/a_158_392# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_35/a_494_366#
+ fine_freq_track_1/sky130_fd_sc_hs__fa_2_1/a_27_378# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_15/a_922_127#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_73/a_494_366# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_7/a_124_78#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_39/a_1434_74# fine_freq_track_1/sky130_fd_sc_hs__nor2b_1_47/a_27_112#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_41/a_1465_471# fine_freq_track_1/sky130_fd_sc_hs__nor3_1_13/Y
+ fine_freq_track_1/sky130_fd_sc_hs__nand2_1_79/a_117_74# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_15/a_1482_48#
+ fine_freq_track_1/sky130_fd_sc_hs__fa_2_17/a_1202_368# fine_freq_track_1/sky130_fd_sc_hs__nor2b_1_13/a_27_112#
+ fine_freq_track_1/sky130_fd_sc_hs__o31ai_1_7/A1 fine_freq_track_1/sky130_fd_sc_hs__dfstp_2_7/a_225_74#
+ fine_freq_track_1/sky130_fd_sc_hs__nand2_1_45/a_117_74# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_43/a_890_138#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_39/a_124_78# fine_freq_track_1/sky130_fd_sc_hs__o211ai_1_9/a_311_74#
+ fine_freq_track_1/sky130_fd_sc_hs__nand2_1_13/a_117_74# fine_freq_track_1/sky130_fd_sc_hs__o21a_1_29/a_320_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_11/a_817_508# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_27/a_910_118#
+ fine_freq_track_1/sky130_fd_sc_hs__nor2_1_19/a_116_368# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_25/a_2026_424#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_9/a_1627_493# fine_freq_track_1/sky130_fd_sc_hs__a22oi_1_11/Y
+ fine_freq_track_1/sky130_fd_sc_hs__fa_2_5/a_1094_347# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_21/a_2010_409#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_17/a_699_463# fine_freq_track_1/sky130_fd_sc_hs__nor3_1_1/a_114_368#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_83/a_124_78# fine_freq_track_1/sky130_fd_sc_hs__fa_2_1/a_701_79#
+ fine_freq_track_1/sky130_fd_sc_hs__nand2_1_7/a_117_74# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_57/a_699_463#
+ fine_freq_track_1/sky130_fd_sc_hs__nor2_1_97/a_116_368# fine_freq_track_1/sky130_fd_sc_hs__o21a_1_73/a_320_74#
+ fine_freq_track_1/sky130_fd_sc_hs__a21oi_1_29/a_29_368# fine_freq_track_1/sky130_fd_sc_hs__a21oi_1_101/a_117_74#
+ fine_freq_track_1/sky130_fd_sc_hs__or2_1_1/B fine_freq_track_1/sky130_fd_sc_hs__o31ai_1_7/a_203_368#
+ fine_freq_track_1/sky130_fd_sc_hs__dfxtp_4_5/a_1034_424# fine_freq_track_1/sky130_fd_sc_hs__nor2b_1_23/a_278_368#
+ fine_freq_track_1/sky130_fd_sc_hs__a31oi_1_1/a_223_74# fine_freq_track_1/sky130_fd_sc_hs__a21oi_1_73/a_29_368#
+ fine_freq_track_1/sky130_fd_sc_hs__nor3_1_15/Y fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_33/a_1647_81#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_39/a_1827_81# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_17/a_507_368#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_35/a_714_127# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_33/a_1224_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_21/a_1736_119# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_37/a_796_463#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_69/a_789_463# fine_freq_track_1/sky130_fd_sc_hs__dfstp_2_7/a_2022_94#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_21/a_1266_119# fine_freq_track_1/sky130_fd_sc_hs__o22ai_1_7/a_142_368#
+ fine_freq_track_1/sky130_fd_sc_hs__nor2_1_7/a_116_368# fine_freq_track_1/sky130_fd_sc_hs__dfstp_2_1/a_1278_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_39/a_120_74# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_49/a_37_78#
+ fine_freq_track_1/sky130_fd_sc_hs__a21oi_1_59/a_117_74# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_49/a_834_355#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_89/a_834_355# fine_freq_track_1/sky130_fd_sc_hs__xor2_1_5/a_194_125#
+ fine_freq_track_1/sky130_fd_sc_hs__nor3_1_11/a_198_368# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_63/a_494_366#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_57/a_1678_395# fine_freq_track_1/sky130_fd_sc_hs__a21oi_1_107/a_29_368#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_5/a_856_304# fine_freq_track_1/sky130_fd_sc_hs__nand2_1_119/a_117_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_5/a_850_127# fine_freq_track_1/sky130_fd_sc_hs__o21a_1_41/X
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_43/a_313_74# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_33/a_890_138#
+ fine_freq_track_1/sky130_fd_sc_hs__a31oi_2_1/a_114_74# fine_freq_track_1/sky130_fd_sc_hs__o21a_1_71/a_376_387#
+ fine_freq_track_1/sky130_fd_sc_hs__nand2_4_3/a_27_74# fine_freq_track_1/sky130_fd_sc_hs__dfxtp_2_11/a_538_429#
+ fine_freq_track_1/sky130_fd_sc_hs__fa_2_5/a_27_378# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_1/a_714_127#
+ fine_freq_track_1/sky130_fd_sc_hs__o21a_1_17/a_83_244# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_17/a_910_118#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_3/D fine_freq_track_1/sky130_fd_sc_hs__nor2_1_47/a_116_368#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_9/a_1224_74# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_65/a_37_78#
+ fine_freq_track_1/sky130_fd_sc_hs__o21a_1_61/a_83_244# fine_freq_track_1/sky130_fd_sc_hs__a22o_1_13/a_230_79#
+ fine_freq_track_1/sky130_fd_sc_hs__nor2_1_87/a_116_368# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_3/a_796_463#
+ fine_freq_track_1/sky130_fd_sc_hs__nand4_1_1/a_373_74# fine_freq_track_1/sky130_fd_sc_hs__dfstp_2_5/a_1356_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_21/Q_N fine_freq_track_1/sky130_fd_sc_hs__nand2_1_17/a_117_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfstp_2_5/a_1521_508# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_45/a_1934_94#
+ fine_freq_track_1/sky130_fd_sc_hs__nor2_1_89/Y fine_freq_track_1/sky130_fd_sc_hs__dfxtp_2_11/a_1019_424#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_49/a_812_138# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_87/a_124_78#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_27/a_856_304# fine_freq_track_1/sky130_fd_sc_hs__o31ai_1_5/a_119_368#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_27/a_850_127# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_89/a_812_138#
+ fine_freq_track_1/sky130_fd_sc_hs__fa_2_5/a_701_79# fine_freq_track_1/sky130_fd_sc_hs__nand2_1_61/a_117_74#
+ fine_freq_track_1/sky130_fd_sc_hs__o21a_1_77/a_320_74# fine_freq_track_1/sky130_fd_sc_hs__nor3_1_3/C
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_53/a_124_78# fine_freq_track_1/sky130_fd_sc_hs__xnor2_1_9/a_138_385#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_23/a_1647_81# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_29/a_1827_81#
+ fine_freq_track_1/sky130_fd_sc_hs__dfxtp_2_9/a_695_459# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_25/a_714_127#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_5/a_832_118# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_51/a_1627_493#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_67/a_1827_81# fine_freq_track_1/sky130_fd_sc_hs__dfxtp_2_1/a_1125_508#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_59/a_789_463# fine_freq_track_1/sky130_fd_sc_hs__fa_2_19/a_27_79#
+ fine_freq_track_1/sky130_fd_sc_hs__sdlclkp_1_1/a_566_74# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_41/a_498_360#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_39/a_1736_119# fine_freq_track_1/sky130_fd_sc_hs__sdlclkp_1_1/a_318_74#
+ fine_freq_track_1/sky130_fd_sc_hs__o21ai_1_5/Y fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_41/a_1350_392#
+ fine_freq_track_1/sky130_fd_sc_hs__a22o_1_11/a_222_392# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_39/a_1266_119#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_11/a_1547_508# fine_freq_track_1/sky130_fd_sc_hs__clkbuf_8_1/a_125_368#
+ fine_freq_track_1/sky130_fd_sc_hs__fa_2_21/a_1119_79# fine_freq_track_1/sky130_fd_sc_hs__dfsbp_2_1/a_595_97#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_21/a_33_74# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_79/a_834_355#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_53/a_494_366# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_19/a_1627_493#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_71/a_2010_409# fine_freq_track_1/sky130_fd_sc_hs__dfxtp_2_11/a_27_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_19/a_37_78# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_35/a_1482_48#
+ fine_freq_track_1/sky130_fd_sc_hs__dfsbp_2_1/a_1453_118# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_29/a_832_118#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_23/a_890_138# fine_freq_track_1/sky130_fd_sc_hs__dfxtp_4_9/a_651_503#
+ fine_freq_track_1/sky130_fd_sc_hs__a21oi_1_93/Y fine_freq_track_1/sky130_fd_sc_hs__o21a_1_61/a_376_387#
+ fine_freq_track_1/sky130_fd_sc_hs__nor3_1_5/B fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_23/a_2026_424#
+ fine_freq_track_1/sky130_fd_sc_hs__dfsbp_2_1/a_731_97# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_7/a_1627_493#
+ fine_freq_track_1/sky130_fd_sc_hs__fa_2_3/a_1094_347# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_9/a_125_78#
+ fine_freq_track_1/sky130_fd_sc_hs__nor2_1_81/Y fine_freq_track_1/sky130_fd_sc_hs__nor2_1_77/a_116_368#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_39/a_2010_409# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_21/a_120_74#
+ fine_freq_track_1/sky130_fd_sc_hs__a21oi_1_41/a_117_74# fine_freq_track_1/sky130_fd_sc_hs__fa_2_5/a_484_347#
+ fine_freq_track_1/sky130_fd_sc_hs__a211oi_1_3/a_354_368# fine_freq_track_1/sky130_fd_sc_hs__fa_2_9/a_27_378#
+ fine_freq_track_1/sky130_fd_sc_hs__a32oi_1_1/a_469_74# fine_freq_track_1/sky130_fd_sc_hs__o21ai_2_1/a_27_74#
+ fine_freq_track_1/sky130_fd_sc_hs__xnor2_1_7/a_376_368# fine_freq_track_1/sky130_fd_sc_hs__dfstp_2_4/a_1521_508#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_31/a_1624_74# fine_freq_track_1/sky130_fd_sc_hs__o21a_1_9/a_320_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_35/a_1934_94# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_91/a_313_74#
+ fine_freq_track_1/sky130_fd_sc_hs__fa_2_3/SUM fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_19/a_1550_119#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_17/a_856_304# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_13/a_125_78#
+ fine_freq_track_1/sky130_fd_sc_hs__a222o_1_1/a_32_74# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_17/a_850_127#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_79/a_812_138# fine_freq_track_1/sky130_fd_sc_hs__o21a_1_65/a_83_244#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_91/a_1350_392# fine_freq_track_1/sky130_fd_sc_hs__nand2_1_101/a_117_74#
+ fine_freq_track_1/sky130_fd_sc_hs__nand4_1_5/a_373_74# fine_freq_track_1/sky130_fd_sc_hs__o211ai_1_11/a_116_368#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_13/a_1647_81# fine_freq_track_1/sky130_fd_sc_hs__dfsbp_2_1/a_27_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_19/a_1827_81# fine_freq_track_1/sky130_fd_sc_hs__fa_2_23/a_487_79#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_15/a_714_127# fine_freq_track_1/sky130_fd_sc_hs__dfstp_2_7/a_1266_341#
+ fine_freq_track_1/sky130_fd_sc_hs__dfstp_2_5/a_612_74# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_37/a_507_368#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_9/a_817_508# fine_freq_track_1/sky130_fd_sc_hs__nand2_1_97/a_117_74#
+ fine_freq_track_1/sky130_fd_sc_hs__conb_1_3/a_165_290# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_91/a_1647_81#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_69/a_1627_493# fine_freq_track_1/sky130_fd_sc_hs__dfsbp_2_1/a_1001_74#
+ fine_freq_track_1/sky130_fd_sc_hs__nor2b_1_33/a_27_112# fine_freq_track_1/sky130_fd_sc_hs__nor2_4_1/a_27_368#
+ fine_freq_track_1/sky130_fd_sc_hs__fa_2_9/a_701_79# fine_freq_track_1/sky130_fd_sc_hs__nand2_1_65/a_117_74#
+ fine_freq_track_1/sky130_fd_sc_hs__xor2_1_3/a_158_392# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_39/a_706_463#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_59/a_1350_392# fine_freq_track_1/sky130_fd_sc_hs__or3b_2_1/a_27_368#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_69/a_834_355# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_29/a_1547_508#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_1/a_1934_94# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_55/a_1678_395#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_3/a_1598_93# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_17/a_1627_493#
+ fine_freq_track_1/sky130_fd_sc_hs__a22oi_1_1/a_159_74# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_83/a_494_366#
+ fine_freq_track_1/sky130_fd_sc_hs__o211ai_1_3/a_116_368# fine_freq_track_1/sky130_fd_sc_hs__o21a_1_15/a_320_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_5/a_841_401# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_7/a_1624_74#
+ fine_freq_track_1/sky130_fd_sc_hs__fa_2_15/a_1202_368# fine_freq_track_1/sky130_fd_sc_hs__dfxtp_4_7/a_206_368#
+ fine_freq_track_1/sky130_fd_sc_hs__o21a_1_11/a_376_387# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_19/a_832_118#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_89/a_2010_409# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_13/a_890_138#
+ fine_freq_track_1/sky130_fd_sc_hs__a21oi_1_15/a_29_368# fine_freq_track_1/sky130_fd_sc_hs__o21a_1_51/a_376_387#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_15/D fine_freq_track_1/sky130_fd_sc_hs__xnor2_1_15/a_376_368#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_1/a_37_78# fine_freq_track_1/sky130_fd_sc_hs__fa_2_9/a_336_347#
+ fine_freq_track_1/sky130_fd_sc_hs__o211ai_1_11/a_31_74# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_91/a_890_138#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_37/a_910_118# fine_freq_track_1/sky130_fd_sc_hs__nor2_1_27/a_116_368#
+ fine_freq_track_1/sky130_fd_sc_hs__nand2_2_7/B fine_freq_track_1/sky130_fd_sc_hs__nor2_1_67/a_116_368#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_27/a_699_463# fine_freq_track_1/sky130_fd_sc_hs__fa_2_7/COUT
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_59/a_37_78# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_37/a_2010_409#
+ fine_freq_track_1/sky130_fd_sc_hs__dfxtp_4_3/a_1034_424# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_29/a_841_401#
+ fine_freq_track_1/sky130_fd_sc_hs__a22o_1_29/a_132_392# fine_freq_track_1/sky130_fd_sc_hs__nor3_1_5/C
+ fine_freq_track_1/sky130_fd_sc_hs__fa_2_19/a_336_347# fine_freq_track_1/sky130_fd_sc_hs__dfstp_2_1/a_1521_508#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_25/a_1934_94# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_21/a_1624_74#
+ fine_freq_track_1/sky130_fd_sc_hs__a22o_1_13/a_52_123# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_5/a_33_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_69/a_812_138# fine_freq_track_1/sky130_fd_sc_hs__a21oi_1_77/a_117_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_13/a_38_78# fine_freq_track_1/sky130_fd_sc_hs__a21oi_1_45/a_117_74#
+ fine_freq_track_1/sky130_fd_sc_hs__a32oi_1_5/a_469_74# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_17/a_313_74#
+ fine_freq_track_1/sky130_fd_sc_hs__fa_2_1/a_683_347# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_47/a_1827_81#
+ fine_freq_track_1/sky130_fd_sc_hs__a21oi_1_11/a_117_74# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_81/a_1647_81#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_39/a_789_463# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_41/a_1224_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_87/a_1827_81# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_67/a_1627_493#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_17/a_125_78# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_73/a_37_78#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_45/a_796_463# fine_freq_track_1/sky130_fd_sc_hs__o22ai_1_7/a_27_74#
+ fine_freq_track_1/sky130_fd_sc_hs__o21a_1_69/a_83_244# fine_freq_track_1/sky130_fd_sc_hs__o211ai_1_3/a_31_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_3/a_910_118# fine_freq_track_1/sky130_fd_sc_hs__nand2_1_105/a_117_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfxtp_2_5/a_644_504# fine_freq_track_1/sky130_fd_sc_hs__o21a_1_35/a_83_244#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_59/a_834_355# fine_freq_track_1/sky130_fd_sc_hs__fa_2_11/a_683_347#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_9/a_494_366# fine_freq_track_1/sky130_fd_sc_hs__dfstp_2_7/a_612_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_53/a_1678_395# fine_freq_track_1/sky130_fd_sc_hs__o21ai_1_1/a_162_368#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_13/a_922_127# fine_freq_track_1/sky130_fd_sc_hs__nor2b_1_9/Y
+ fine_freq_track_1/sky130_fd_sc_hs__nor2b_1_37/a_27_112# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_3/a_38_78#
+ fine_freq_track_1/sky130_fd_sc_hs__a22o_1_5/a_132_392# fine_freq_track_1/sky130_fd_sc_hs__nand2_1_69/a_117_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfxtp_4_7/a_437_503# fine_freq_track_1/sky130_fd_sc_hs__o21a_1_41/a_376_387#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_47/a_832_118# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_29/a_124_78#
+ fine_freq_track_1/sky130_fd_sc_hs__fa_2_9/a_1202_368# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_81/a_890_138#
+ fine_freq_track_1/sky130_fd_sc_hs__fa_2_5/a_27_79# fine_freq_track_1/sky130_fd_sc_hs__fa_2_1/a_1094_347#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_5/a_1627_493# fine_freq_track_1/sky130_fd_sc_hs__o21a_1_19/a_320_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfxtp_4_5/a_735_102# fine_freq_track_1/sky130_fd_sc_hs__a21oi_1_123/a_117_74#
+ fine_freq_track_1/sky130_fd_sc_hs__nor2_1_57/a_116_368# fine_freq_track_1/sky130_fd_sc_hs__a21oi_1_19/a_29_368#
+ fine_freq_track_1/sky130_fd_sc_hs__o21a_1_63/a_320_74# fine_freq_track_1/sky130_fd_sc_hs__dfxtp_4_2/a_1034_424#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_19/a_841_401# fine_freq_track_1/sky130_fd_sc_hs__a22o_1_19/a_132_392#
+ fine_freq_track_1/sky130_fd_sc_hs__o31ai_1_5/a_203_368# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_15/a_1934_94#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_11/a_1624_74# fine_freq_track_1/sky130_fd_sc_hs__dfstp_2_4/a_398_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_17/a_1550_119# fine_freq_track_1/sky130_fd_sc_hs__nor2b_1_17/Y
+ fine_freq_track_1/sky130_fd_sc_hs__a21oi_1_63/a_29_368# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_59/a_812_138#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_37/a_856_304# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_5/a_1434_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_37/a_850_127# fine_freq_track_1/sky130_fd_sc_hs__dfxtp_4_7/a_27_74#
+ fine_freq_track_1/sky130_fd_sc_hs__nand2_2_11/a_27_74# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_7/a_1647_81#
+ fine_freq_track_1/sky130_fd_sc_hs__nand2_2_1/a_27_74# fine_freq_track_1/sky130_fd_sc_hs__fa_2_5/a_1205_79#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_37/a_1827_81# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_3/a_1827_81#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_39/D fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_29/a_789_463#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_71/a_1647_81# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_77/a_1827_81#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_37/a_1736_119# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_41/Q_N
+ fine_freq_track_1/sky130_fd_sc_hs__o31ai_1_1/a_114_74# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_67/a_789_463#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_37/a_1266_119# fine_freq_track_1/sky130_fd_sc_hs__dfstp_2_1/a_27_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_33/Q_N fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_29/a_120_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_57/a_1350_392# fine_freq_track_1/sky130_fd_sc_hs__a32oi_1_9/a_469_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_27/a_1547_508# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_23/Q_N
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_15/a_1627_493# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_29/a_1434_74#
+ fine_freq_track_1/sky130_fd_sc_hs__a21oi_1_93/a_117_74# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_43/a_37_78#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_43/a_922_127# fine_freq_track_1/sky130_fd_sc_hs__fa_2_13/a_1202_368#
+ fine_freq_track_1/sky130_fd_sc_hs__a211oi_1_3/a_159_74# fine_freq_track_1/sky130_fd_sc_hs__nand2_1_109/a_117_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_87/a_2010_409# fine_freq_track_1/sky130_fd_sc_hs__o21a_1_31/a_376_387#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_43/a_1482_48# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_33/a_313_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfxtp_2_1/a_206_368# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_7/a_890_138#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_21/a_2026_424# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_71/a_890_138#
+ fine_freq_track_1/sky130_fd_sc_hs__xnor2_1_3/Y fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_33/a_125_78#
+ fine_freq_track_1/sky130_fd_sc_hs__and2_2_3/a_31_74# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_39/a_2026_424#
+ fine_freq_track_1/sky130_fd_sc_hs__nor3_1_1/A fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_1/a_796_463#
+ fine_freq_track_1/sky130_fd_sc_hs__o21a_1_51/a_83_244# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_85/a_699_463#
+ fine_freq_track_1/sky130_fd_sc_hs__dfstp_2_4/a_1356_74# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_47/a_841_401#
+ fine_freq_track_1/sky130_fd_sc_hs__nor2_1_121/a_116_368# fine_freq_track_1/sky130_fd_sc_hs__nor3_1_5/a_198_368#
+ fine_freq_track_1/sky130_fd_sc_hs__a22oi_1_9/a_159_74# fine_freq_track_1/sky130_fd_sc_hs__a22o_1_7/a_222_392#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_9/a_1678_395# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_45/a_1598_93#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_77/a_124_78# fine_freq_track_1/sky130_fd_sc_hs__nand2_1_51/a_117_74#
+ fine_freq_track_1/sky130_fd_sc_hs__o21a_1_67/a_320_74# fine_freq_track_1/sky130_fd_sc_hs__a22oi_1_3/a_339_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_21/a_1647_81# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_9/a_1465_471#
+ fine_freq_track_1/sky130_fd_sc_hs__dfxtp_2_7/a_695_459# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_11/a_124_78#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_19/a_789_463# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_61/a_1647_81#
+ fine_freq_track_1/sky130_fd_sc_hs__fa_2_17/a_27_378# fine_freq_track_1/sky130_fd_sc_hs__a21oi_1_67/a_29_368#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_25/a_796_463# fine_freq_track_1/sky130_fd_sc_hs__nor2_1_57/B
+ fine_freq_track_1/sky130_fd_sc_hs__nand2b_1_1/a_27_112# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_67/a_37_78#
+ fine_freq_track_1/sky130_fd_sc_hs__a21oi_1_33/a_29_368# fine_freq_track_1/sky130_fd_sc_hs__sdlclkp_4_1/a_744_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_39/a_834_355# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_39/a_319_360#
+ fine_freq_track_1/sky130_fd_sc_hs__a32oi_1_3/a_391_74# fine_freq_track_1/sky130_fd_sc_hs__fa_2_13/a_27_79#
+ fine_freq_track_1/sky130_fd_sc_hs__nand4_1_5/D fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_19/a_1434_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_33/a_922_127# fine_freq_track_1/sky130_fd_sc_hs__fa_2_11/a_1202_368#
+ fine_freq_track_1/sky130_fd_sc_hs__fa_2_7/SUM fine_freq_track_1/sky130_fd_sc_hs__xor2_1_11/a_194_125#
+ fine_freq_track_1/sky130_fd_sc_hs__o21a_1_21/a_376_387# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_27/a_832_118#
+ fine_freq_track_1/sky130_fd_sc_hs__dfsbp_2_1/a_706_463# fine_freq_track_1/sky130_fd_sc_hs__fa_2_23/a_1094_347#
+ fine_freq_track_1/sky130_fd_sc_hs__fa_2_17/a_701_79# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_21/a_890_138#
+ fine_freq_track_1/sky130_fd_sc_hs__fa_2_7/a_1202_368# fine_freq_track_1/sky130_fd_sc_hs__dfsbp_2_1/a_1261_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfxtp_2_11/a_1172_124# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_61/a_890_138#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_5/a_313_74# fine_freq_track_1/sky130_fd_sc_hs__nand2_4_9/A
+ fine_freq_track_1/sky130_fd_sc_hs__nor3_1_7/Y fine_freq_track_1/sky130_fd_sc_hs__a21oi_1_97/a_117_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_83/a_37_78# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_57/D
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_27/a_300_74# fine_freq_track_1/sky130_fd_sc_hs__nor2_1_37/a_116_368#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_45/a_910_118# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_35/a_2010_409#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_45/a_120_74# fine_freq_track_1/sky130_fd_sc_hs__nor2_1_75/a_116_368#
+ fine_freq_track_1/sky130_fd_sc_hs__dfxtp_2_5/a_538_429# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_7/a_120_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_1/a_699_463# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_11/a_120_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_75/a_699_463# fine_freq_track_1/sky130_fd_sc_hs__a21oi_1_31/a_117_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_25/a_33_74# fine_freq_track_1/sky130_fd_sc_hs__nor2_1_111/a_116_368#
+ fine_freq_track_1/sky130_fd_sc_hs__o21ai_1_1/a_27_74# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_37/a_125_78#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_35/a_1598_93# fine_freq_track_1/sky130_fd_sc_hs__nor2b_1_41/a_278_368#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_81/a_313_74# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_39/a_812_138#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_1/a_300_74# fine_freq_track_1/sky130_fd_sc_hs__o21a_1_55/a_83_244#
+ fine_freq_track_1/sky130_fd_sc_hs__fa_2_15/a_484_347# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_17/a_1827_81#
+ fine_freq_track_1/sky130_fd_sc_hs__dfstp_2_5/a_1266_341# fine_freq_track_1/sky130_fd_sc_hs__fa_2_13/a_487_79#
+ fine_freq_track_1/sky130_fd_sc_hs__dfxtp_4_9/a_1226_296# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_13/a_714_127#
+ fine_freq_track_1/sky130_fd_sc_hs__nor2_1_15/B fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_51/a_1647_81#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_57/a_1827_81# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_65/a_1627_493#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_9/Q_N fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_7/a_817_508#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_15/a_796_463# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_35/a_1736_119#
+ fine_freq_track_1/sky130_fd_sc_hs__nor3_1_15/B fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_47/a_789_463#
+ fine_freq_track_1/sky130_fd_sc_hs__nor2b_1_23/a_27_112# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_31/a_498_360#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_35/a_1266_119# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_87/a_789_463#
+ fine_freq_track_1/sky130_fd_sc_hs__inv_4_27/Y fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_55/a_1350_392#
+ fine_freq_track_1/sky130_fd_sc_hs__nand2_1_55/a_117_74# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_47/a_38_78#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_29/a_834_355# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_47/a_124_78#
+ fine_freq_track_1/sky130_fd_sc_hs__a22oi_1_7/a_339_74# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_67/a_834_355#
+ fine_freq_track_1/sky130_fd_sc_hs__fa_2_21/a_683_347# fine_freq_track_1/sky130_fd_sc_hs__o21a_1_37/a_320_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_51/a_1678_395# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_43/a_494_366#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_23/a_922_127# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_1/a_1598_93#
+ fine_freq_track_1/sky130_fd_sc_hs__a22oi_1_23/a_71_368# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_47/a_1434_74#
+ fine_freq_track_1/sky130_fd_sc_hs__nand2b_1_5/a_27_112# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_85/a_2010_409#
+ fine_freq_track_1/sky130_fd_sc_hs__a21oi_1_37/a_29_368# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_23/a_1482_48#
+ fine_freq_track_1/sky130_fd_sc_hs__xnor2_1_7/a_112_119# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_17/a_832_118#
+ fine_freq_track_1/sky130_fd_sc_hs__a32oi_1_7/a_391_74# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_51/a_890_138#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_3/a_1627_493# fine_freq_track_1/sky130_fd_sc_hs__a21oi_1_83/a_29_368#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_19/a_1678_395# fine_freq_track_1/sky130_fd_sc_hs__nand3b_2_1/a_27_94#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_3/a_507_368# fine_freq_track_1/sky130_fd_sc_hs__fa_2_9/a_992_347#
+ fine_freq_track_1/sky130_fd_sc_hs__dfxtp_4_9/a_696_458# fine_freq_track_1/sky130_fd_sc_hs__o21a_1_7/a_376_387#
+ fine_freq_track_1/sky130_fd_sc_hs__dfxtp_4_2/Q fine_freq_track_1/sky130_fd_sc_hs__a32oi_1_3/a_27_368#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_25/a_699_463# fine_freq_track_1/sky130_fd_sc_hs__nor2b_1_9/a_278_368#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_7/a_498_360# fine_freq_track_1/sky130_fd_sc_hs__or3b_2_1/a_190_260#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_65/a_699_463# fine_freq_track_1/sky130_fd_sc_hs__nor2_1_101/a_116_368#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_27/a_841_401# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_9/a_313_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_5/a_706_463# fine_freq_track_1/sky130_fd_sc_hs__fa_2_19/a_992_347#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_15/a_1550_119# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_7/a_1678_395#
+ fine_freq_track_1/sky130_fd_sc_hs__nor2b_1_31/a_278_368# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_25/a_1598_93#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_29/a_812_138# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_49/a_120_74#
+ fine_freq_track_1/sky130_fd_sc_hs__maj3_1_3/a_403_136# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_67/a_812_138#
+ fine_freq_track_1/sky130_fd_sc_hs__dfxtp_2_1/a_708_101# fine_freq_track_1/sky130_fd_sc_hs__dfstp_2_5/a_781_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_7/a_1465_471# fine_freq_track_1/sky130_fd_sc_hs__dfstp_2_4/a_1266_341#
+ fine_freq_track_1/sky130_fd_sc_hs__o22ai_1_5/a_340_368# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_41/a_1647_81#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_63/a_1627_493# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_43/a_300_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_43/a_714_127# fine_freq_track_1/sky130_fd_sc_hs__a21oi_1_117/a_29_368#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_37/a_789_463# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_85/a_313_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_3/a_789_463# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_21/a_498_360#
+ fine_freq_track_1/sky130_fd_sc_hs__nor3_1_15/a_114_368# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_77/a_789_463#
+ fine_freq_track_1/sky130_fd_sc_hs__xnor2_1_15/a_112_119# fine_freq_track_1/sky130_fd_sc_hs__o21a_1_59/a_83_244#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_53/a_1350_392# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_29/a_706_463#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_19/a_834_355# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_1/a_910_118#
+ fine_freq_track_1/sky130_fd_sc_hs__dfxtp_2_3/a_644_504# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_25/a_1547_508#
+ fine_freq_track_1/sky130_fd_sc_hs__a21oi_1_91/Y fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_13/a_1627_493#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_33/a_494_366# fine_freq_track_1/sky130_fd_sc_hs__dfstp_2_7/a_1489_118#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_69/a_1678_395# fine_freq_track_1/sky130_fd_sc_hs__nor2b_1_27/a_27_112#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_7/a_33_74# fine_freq_track_1/sky130_fd_sc_hs__a22o_1_23/a_230_79#
+ fine_freq_track_1/sky130_fd_sc_hs__inv_4_25/Y fine_freq_track_1/sky130_fd_sc_hs__nand2_1_59/a_117_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_13/a_1482_48# fine_freq_track_1/sky130_fd_sc_hs__dfxtp_2_3/a_27_74#
+ fine_freq_track_1/sky130_fd_sc_hs__fa_2_21/a_1094_347# fine_freq_track_1/sky130_fd_sc_hs__inv_4_57/Y
+ fine_freq_track_1/sky130_fd_sc_hs__fa_2_5/a_1202_368# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_41/a_890_138#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_19/a_124_78# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_17/a_1678_395#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_37/a_2026_424# fine_freq_track_1/sky130_fd_sc_hs__or2_1_3/a_152_368#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_25/a_910_118# fine_freq_track_1/sky130_fd_sc_hs__o21a_1_55/X
+ fine_freq_track_1/sky130_fd_sc_hs__nor2_1_17/a_116_368# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_33/a_2010_409#
+ fine_freq_track_1/sky130_fd_sc_hs__dfxtp_2_9/a_1019_424# fine_freq_track_1/sky130_fd_sc_hs__nand2b_1_9/a_27_112#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_77/a_37_78# fine_freq_track_1/sky130_fd_sc_hs__nor2b_1_5/Y
+ fine_freq_track_1/sky130_fd_sc_hs__a21oi_1_113/a_117_74# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_15/a_699_463#
+ fine_freq_track_1/sky130_fd_sc_hs__o211ai_1_5/a_31_74# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_55/a_699_463#
+ fine_freq_track_1/sky130_fd_sc_hs__nor2_1_95/a_116_368# fine_freq_track_1/sky130_fd_sc_hs__o21a_1_53/a_320_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_17/a_841_401# fine_freq_track_1/sky130_fd_sc_hs__nor2b_1_15/Y
+ fine_freq_track_1/sky130_fd_sc_hs__dfstp_2_7/a_1057_118# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_13/a_1550_119#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_13/a_1934_94# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_15/a_1598_93#
+ fine_freq_track_1/sky130_fd_sc_hs__nor2b_1_21/a_278_368# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_17/Q_N
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_19/a_812_138# fine_freq_track_1/sky130_fd_sc_hs__a32oi_1_7/a_27_368#
+ fine_freq_track_1/sky130_fd_sc_hs__dfstp_2_1/a_1266_341# fine_freq_track_1/sky130_fd_sc_hs__dfxtp_4_7/a_1226_296#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_31/a_1647_81# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_33/a_1736_119#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_33/a_714_127# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_31/a_1224_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_11/a_498_360# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_33/a_1266_119#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_35/a_796_463# fine_freq_track_1/sky130_fd_sc_hs__o22ai_1_5/a_142_368#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_19/a_706_463# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_19/a_120_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfstp_2_7/a_781_74# fine_freq_track_1/sky130_fd_sc_hs__a21oi_1_39/a_117_74#
+ fine_freq_track_1/sky130_fd_sc_hs__a2bb2oi_1_1/a_399_368# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_47/a_834_355#
+ fine_freq_track_1/sky130_fd_sc_hs__o21ai_1_11/a_162_368# fine_freq_track_1/sky130_fd_sc_hs__fa_2_15/a_1205_79#
+ fine_freq_track_1/sky130_fd_sc_hs__o21a_1_3/a_83_244# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_23/a_494_366#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_87/a_834_355# fine_freq_track_1/sky130_fd_sc_hs__xor2_1_3/a_194_125#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_67/a_1678_395# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_89/a_313_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_27/a_1434_74# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_41/a_922_127#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_13/a_300_74# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_83/a_2010_409#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_3/a_856_304# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_3/a_850_127#
+ fine_freq_track_1/sky130_fd_sc_hs__nand2_2_13/a_27_74# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_37/a_832_118#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_23/a_313_74# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_31/a_890_138#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_1/a_1627_493# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_15/a_910_118#
+ fine_freq_track_1/sky130_fd_sc_hs__dfxtp_2_7/a_1019_424# fine_freq_track_1/sky130_fd_sc_hs__nor2b_1_3/a_27_112#
+ fine_freq_track_1/sky130_fd_sc_hs__a22o_1_27/a_230_79# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_7/a_1224_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_45/a_699_463# fine_freq_track_1/sky130_fd_sc_hs__o21a_1_41/a_83_244#
+ fine_freq_track_1/sky130_fd_sc_hs__nor2_1_85/a_116_368# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_9/a_1350_392#
+ fine_freq_track_1/sky130_fd_sc_hs__dfxtp_2_11/a_1217_314# fine_freq_track_1/sky130_fd_sc_hs__dfstp_2_1/a_1356_74#
+ fine_freq_track_1/sky130_fd_sc_hs__nand4_2_1/a_27_74# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_3/a_124_78#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_5/a_1678_395# fine_freq_track_1/sky130_fd_sc_hs__nor2b_1_11/a_278_368#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_43/a_1934_94# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_77/D
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_47/a_812_138# fine_freq_track_1/sky130_fd_sc_hs__dfxtp_2_9/a_431_508#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_87/a_812_138# fine_freq_track_1/sky130_fd_sc_hs__dfstp_2_4/a_225_74#
+ fine_freq_track_1/sky130_fd_sc_hs__o21a_1_57/a_320_74# fine_freq_track_1/sky130_fd_sc_hs__a32oi_1_3/a_119_74#
+ fine_freq_track_1/sky130_fd_sc_hs__xnor2_1_7/a_138_385# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_27/a_1827_81#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_23/a_714_127# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_31/a_1736_119#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_3/a_832_118# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_17/a_789_463#
+ fine_freq_track_1/sky130_fd_sc_hs__a2bb2oi_1_1/a_488_74# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_21/a_1224_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_45/a_507_368# fine_freq_track_1/sky130_fd_sc_hs__a21oi_1_57/a_29_368#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_31/a_1266_119# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_57/a_789_463#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_23/a_1547_508# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_47/a_706_463#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_37/a_834_355# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_11/a_1627_493#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_13/a_494_366# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_3/a_834_355#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_77/a_834_355# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_61/a_37_78#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_17/a_1434_74# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_31/a_922_127#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_91/a_494_366# fine_freq_track_1/sky130_fd_sc_hs__a2bb2oi_1_1/a_126_112#
+ fine_freq_track_1/sky130_fd_sc_hs__xnor2_1_3/a_293_74# fine_freq_track_1/sky130_fd_sc_hs__fa_2_3/a_1202_368#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_33/a_1482_48# fine_freq_track_1/sky130_fd_sc_hs__dfxtp_4_7/a_651_503#
+ fine_freq_track_1/sky130_fd_sc_hs__o21a_1_7/a_83_244# fine_freq_track_1/sky130_fd_sc_hs__a22o_1_23/a_52_123#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_15/a_1678_395# fine_freq_track_1/sky130_fd_sc_hs__dfxtp_4_9/a_544_485#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_35/a_2026_424# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_31/a_2010_409#
+ fine_freq_track_1/sky130_fd_sc_hs__a21oi_1_87/a_117_74# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_39/a_817_508#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_19/a_1465_471# fine_freq_track_1/sky130_fd_sc_hs__a222oi_1_1/a_461_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_17/a_300_74# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_35/a_120_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_49/a_2010_409# fine_freq_track_1/sky130_fd_sc_hs__a21oi_1_53/a_117_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_35/a_699_463# fine_freq_track_1/sky130_fd_sc_hs__dfxtp_2_3/a_538_429#
+ fine_freq_track_1/sky130_fd_sc_hs__xnor2_1_15/a_138_385# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_27/a_313_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_73/a_699_463# fine_freq_track_1/sky130_fd_sc_hs__fa_2_3/a_484_347#
+ fine_freq_track_1/sky130_fd_sc_hs__a21oi_1_21/a_117_74# fine_freq_track_1/sky130_fd_sc_hs__a211oi_1_1/a_354_368#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_11/a_1550_119# fine_freq_track_1/sky130_fd_sc_hs__o2bb2ai_1_1/a_397_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_37/a_841_401# fine_freq_track_1/sky130_fd_sc_hs__o21ai_2_1/a_116_368#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_39/a_1624_74# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_5/a_319_360#
+ fine_freq_track_1/sky130_fd_sc_hs__xnor2_1_5/a_376_368# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_33/a_1934_94#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_71/a_313_74# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_37/a_812_138#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_19/D fine_freq_track_1/sky130_fd_sc_hs__a21oi_1_3/a_117_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_3/a_812_138# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_25/a_38_78#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_77/a_812_138# fine_freq_track_1/sky130_fd_sc_hs__o21a_1_45/a_83_244#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_5/a_1465_471# fine_freq_track_1/sky130_fd_sc_hs__dfxtp_4_5/a_1226_296#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_11/a_1647_81# fine_freq_track_1/sky130_fd_sc_hs__fa_2_9/a_1119_79#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_61/a_1627_493# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_9/a_1482_48#
+ fine_freq_track_1/sky130_fd_sc_hs__o21a_1_11/a_83_244# fine_freq_track_1/sky130_fd_sc_hs__nor2b_2_1/a_27_392#
+ fine_freq_track_1/sky130_fd_sc_hs__o21a_1_1/a_320_74# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_11/a_1224_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_35/a_507_368# fine_freq_track_1/sky130_fd_sc_hs__conb_1_1/a_165_290#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_51/a_1350_392# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_21/a_1547_508#
+ fine_freq_track_1/sky130_fd_sc_hs__xor2_1_1/a_158_392# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_37/a_124_78#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_29/a_319_360# fine_freq_track_1/sky130_fd_sc_hs__a32oi_1_7/a_119_74#
+ fine_freq_track_1/sky130_fd_sc_hs__fa_2_19/a_1119_79# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_27/a_33_74#
+ fine_freq_track_1/sky130_fd_sc_hs__o21a_1_27/a_320_74# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_29/a_1627_493#
+ fine_freq_track_1/sky130_fd_sc_hs__dfstp_2_7/a_1596_118# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_21/a_922_127#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_81/a_494_366# fine_freq_track_1/sky130_fd_sc_hs__o211ai_1_1/a_116_368#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_81/a_2010_409# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_3/a_841_401#
+ fine_freq_track_1/sky130_fd_sc_hs__a22oi_1_13/a_71_368# fine_freq_track_1/sky130_fd_sc_hs__dfxtp_4_5/a_206_368#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_19/a_1350_392# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_79/D
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_11/a_890_138# fine_freq_track_1/sky130_fd_sc_hs__xnor2_1_13/a_376_368#
+ fine_freq_track_1/sky130_fd_sc_hs__fa_2_23/a_27_378# fine_freq_track_1/sky130_fd_sc_hs__fa_2_7/a_336_347#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_1/a_507_368# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_17/a_1465_471#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_29/a_817_508# fine_freq_track_1/sky130_fd_sc_hs__dfstp_2_7/a_1566_92#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_35/a_910_118# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_7/a_1350_392#
+ fine_freq_track_1/sky130_fd_sc_hs__nor2_1_65/a_116_368# fine_freq_track_1/sky130_fd_sc_hs__xnor2_1_7/a_293_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_43/a_33_74# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_63/a_699_463#
+ fine_freq_track_1/sky130_fd_sc_hs__a22o_1_27/a_52_123# fine_freq_track_1/sky130_fd_sc_hs__maj3_1_3/a_406_384#
+ fine_freq_track_1/sky130_fd_sc_hs__a22o_1_27/a_132_392# fine_freq_track_1/sky130_fd_sc_hs__fa_2_17/a_336_347#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_23/a_1934_94# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_29/a_1550_119#
+ fine_freq_track_1/sky130_fd_sc_hs__maj3_1_1/a_403_136# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_45/a_856_304#
+ fine_freq_track_1/sky130_fd_sc_hs__fa_2_23/a_701_79# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_45/a_850_127#
+ fine_freq_track_1/sky130_fd_sc_hs__a21oi_1_25/a_117_74# fine_freq_track_1/sky130_fd_sc_hs__sdlclkp_1_1/a_667_80#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_33/a_300_74# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_25/a_507_368#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_79/a_1627_493# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_41/a_714_127#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_5/a_125_78# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_49/a_1736_119#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_75/a_313_74# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_47/Q_N
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_85/a_1827_81# fine_freq_track_1/sky130_fd_sc_hs__xor2_1_9/a_355_368#
+ fine_freq_track_1/sky130_fd_sc_hs__a21oi_1_7/a_117_74# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_43/a_796_463#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_49/a_1266_119# fine_freq_track_1/sky130_fd_sc_hs__o21a_1_49/a_83_244#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_69/a_1350_392# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_27/a_706_463#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_17/a_834_355# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_19/a_319_360#
+ fine_freq_track_1/sky130_fd_sc_hs__a22o_1_3/a_230_79# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_39/a_1547_508#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_57/a_834_355# fine_freq_track_1/sky130_fd_sc_hs__dfstp_2_5/a_1489_118#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_41/a_125_78# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_65/a_1678_395#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_7/a_494_366# fine_freq_track_1/sky130_fd_sc_hs__o21a_1_5/a_320_74#
+ fine_freq_track_1/sky130_fd_sc_hs__nor2b_1_49/a_27_112# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_11/a_922_127#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_71/a_494_366# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_55/a_37_78#
+ fine_freq_track_1/sky130_fd_sc_hs__and2_2_3/a_118_74# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_37/a_1434_74#
+ fine_freq_track_1/sky130_fd_sc_hs__nor2b_1_17/a_27_112# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_17/a_1350_392#
+ fine_freq_track_1/sky130_fd_sc_hs__a22o_1_3/a_132_392# fine_freq_track_1/sky130_fd_sc_hs__nand2_1_49/a_117_74#
+ fine_freq_track_1/sky130_fd_sc_hs__fa_2_1/a_1202_368# fine_freq_track_1/sky130_fd_sc_hs__a222o_1_1/a_119_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfxtp_4_5/a_437_503# fine_freq_track_1/sky130_fd_sc_hs__conb_1_3/LO
+ fine_freq_track_1/sky130_fd_sc_hs__nor2b_2_1/a_228_368# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_45/a_832_118#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_33/a_2026_424# fine_freq_track_1/sky130_fd_sc_hs__nand2_1_93/a_117_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfxtp_2_5/a_1019_424# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_19/a_817_508#
+ fine_freq_track_1/sky130_fd_sc_hs__a22oi_1_17/a_71_368# fine_freq_track_1/sky130_fd_sc_hs__sdlclkp_1_1/a_116_424#
+ fine_freq_track_1/sky130_fd_sc_hs__nand2_1_9/a_117_74# fine_freq_track_1/sky130_fd_sc_hs__nor3_1_9/a_114_368#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_47/a_2010_409# fine_freq_track_1/sky130_fd_sc_hs__a21oi_1_103/a_117_74#
+ fine_freq_track_1/sky130_fd_sc_hs__nor2_1_55/a_116_368# fine_freq_track_1/sky130_fd_sc_hs__a2bb2oi_1_1/a_117_392#
+ fine_freq_track_1/sky130_fd_sc_hs__nor2_1_53/Y fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_53/a_699_463#
+ fine_freq_track_1/sky130_fd_sc_hs__dfstp_2_5/a_1057_118# fine_freq_track_1/sky130_fd_sc_hs__o21a_1_43/a_320_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_3/a_1678_395# fine_freq_track_1/sky130_fd_sc_hs__a22o_1_17/a_132_392#
+ fine_freq_track_1/sky130_fd_sc_hs__o22ai_1_3/a_27_74# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_13/a_1598_93#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_17/a_812_138# fine_freq_track_1/sky130_fd_sc_hs__nor2b_1_27/Y
+ fine_freq_track_1/sky130_fd_sc_hs__a21oi_1_43/a_29_368# fine_freq_track_1/sky130_fd_sc_hs__nor2_1_13/B
+ fine_freq_track_1/sky130_fd_sc_hs__nor4_1_1/Y fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_57/a_812_138#
+ fine_freq_track_1/sky130_fd_sc_hs__dfxtp_2_11/a_695_459# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_3/a_1465_471#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_35/a_856_304# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_35/a_850_127#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_3/a_1434_74# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_11/a_33_74#
+ fine_freq_track_1/sky130_fd_sc_hs__fa_2_3/a_1205_79# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_5/a_1647_81#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_15/a_507_368# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_31/a_714_127#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_1/a_1827_81# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_27/a_789_463#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_47/a_1736_119# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_75/a_1827_81#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_47/a_1266_119# fine_freq_track_1/sky130_fd_sc_hs__o211ai_1_9/a_31_74#
+ fine_freq_track_1/sky130_fd_sc_hs__nor2_1_5/a_116_368# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_67/a_1350_392#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_17/a_706_463# fine_freq_track_1/sky130_fd_sc_hs__a22o_1_29/a_222_392#
+ fine_freq_track_1/sky130_fd_sc_hs__a21oi_1_29/a_117_74# fine_freq_track_1/sky130_fd_sc_hs__fa_2_1/a_27_79#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_47/a_319_360# fine_freq_track_1/sky130_fd_sc_hs__dfstp_2_4/a_1489_118#
+ fine_freq_track_1/sky130_fd_sc_hs__a211oi_4_1/a_77_368# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_21/a_494_366#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_63/a_1678_395# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_27/a_1627_493#
+ fine_freq_track_1/sky130_fd_sc_hs__dfxtp_2_9/a_1172_124# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_37/a_300_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_61/a_494_366# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_79/a_313_74#
+ fine_freq_track_1/sky130_fd_sc_hs__nor2_2_3/A fine_freq_track_1/sky130_fd_sc_hs__a21oi_1_73/a_117_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_35/a_38_78# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_1/a_856_304#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_1/a_850_127# fine_freq_track_1/sky130_fd_sc_hs__a22o_1_7/a_230_79#
+ fine_freq_track_1/sky130_fd_sc_hs__nor2b_1_43/Y fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_41/a_1482_48#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_13/a_1678_395# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_13/a_313_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_45/a_125_78# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_5/a_890_138#
+ fine_freq_track_1/sky130_fd_sc_hs__dfxtp_2_3/a_1019_424# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_15/a_1465_471#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_3/Q_N fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_49/a_817_508#
+ fine_freq_track_1/sky130_fd_sc_hs__a22o_1_17/a_230_79# fine_freq_track_1/sky130_fd_sc_hs__or2_1_1/a_63_368#
+ fine_freq_track_1/sky130_fd_sc_hs__nor2_1_45/a_116_368# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_5/a_1350_392#
+ fine_freq_track_1/sky130_fd_sc_hs__o21a_1_31/a_83_244# fine_freq_track_1/sky130_fd_sc_hs__dfstp_2_4/a_1057_118#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_37/a_33_74# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_83/a_699_463#
+ fine_freq_track_1/sky130_fd_sc_hs__dfstp_2_4/a_612_74# fine_freq_track_1/sky130_fd_sc_hs__a22oi_1_23/a_159_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_45/a_841_401# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_27/a_1550_119#
+ fine_freq_track_1/sky130_fd_sc_hs__nor3_1_3/a_198_368# fine_freq_track_1/sky130_fd_sc_hs__dfxtp_4_9/a_1141_508#
+ fine_freq_track_1/sky130_fd_sc_hs__a22o_1_5/a_222_392# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_41/a_1934_94#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_43/a_1598_93# fine_freq_track_1/sky130_fd_sc_hs__nand2_1_63/a_117_74#
+ fine_freq_track_1/sky130_fd_sc_hs__a21oi_1_107/a_117_74# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_57/a_124_78#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_1/a_1465_471# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_25/a_856_304#
+ fine_freq_track_1/sky130_fd_sc_hs__o31ai_1_3/a_119_368# fine_freq_track_1/sky130_fd_sc_hs__dfxtp_2_7/a_431_508#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_25/a_850_127# fine_freq_track_1/sky130_fd_sc_hs__dfxtp_4_3/a_1226_296#
+ fine_freq_track_1/sky130_fd_sc_hs__nand2_1_31/a_117_74# fine_freq_track_1/sky130_fd_sc_hs__o21a_1_47/a_320_74#
+ fine_freq_track_1/sky130_fd_sc_hs__fa_2_23/a_484_347# fine_freq_track_1/sky130_fd_sc_hs__a21oi_1_79/a_29_368#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_25/a_1827_81# fine_freq_track_1/sky130_fd_sc_hs__nand2_2_7/a_27_74#
+ fine_freq_track_1/sky130_fd_sc_hs__o21a_1_13/a_320_74# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_77/a_1627_493#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_21/a_714_127# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_1/a_832_118#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_65/a_1827_81# fine_freq_track_1/sky130_fd_sc_hs__a21oi_1_47/a_29_368#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_23/a_796_463# fine_freq_track_1/sky130_fd_sc_hs__dfstp_2_5/a_767_384#
+ fine_freq_track_1/sky130_fd_sc_hs__a22o_1_19/a_222_392# fine_freq_track_1/sky130_fd_sc_hs__dfstp_2_7/a_27_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfstp_2_1/a_1489_118# fine_freq_track_1/sky130_fd_sc_hs__a21oi_1_91/a_29_368#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_25/a_1627_493# fine_freq_track_1/sky130_fd_sc_hs__dfxtp_2_7/a_1172_124#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_51/a_494_366# fine_freq_track_1/sky130_fd_sc_hs__fa_2_23/a_1202_368#
+ fine_freq_track_1/sky130_fd_sc_hs__a222o_1_1/a_651_74# fine_freq_track_1/sky130_fd_sc_hs__a22o_1_3/a_52_123#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_15/a_1350_392# fine_freq_track_1/sky130_fd_sc_hs__fa_2_3/a_487_79#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_25/a_832_118# fine_freq_track_1/sky130_fd_sc_hs__o21a_1_69/a_376_387#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_31/a_2026_424# fine_freq_track_1/sky130_fd_sc_hs__nor2_2_3/B
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_43/a_910_118# fine_freq_track_1/sky130_fd_sc_hs__nor2_1_35/a_116_368#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_49/a_313_74# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_25/a_120_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_9/a_699_463# fine_freq_track_1/sky130_fd_sc_hs__nor2_1_73/a_116_368#
+ fine_freq_track_1/sky130_fd_sc_hs__dfstp_2_1/a_1057_118# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_1/a_1678_395#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_17/D fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_63/a_37_78#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_9/a_922_127# fine_freq_track_1/sky130_fd_sc_hs__nor2b_1_49/a_278_368#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_31/a_1934_94# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_33/a_1598_93#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_61/a_313_74# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_15/a_856_304#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_15/a_850_127# fine_freq_track_1/sky130_fd_sc_hs__dfxtp_4_2/a_1226_296#
+ fine_freq_track_1/sky130_fd_sc_hs__o21a_1_39/X fine_freq_track_1/sky130_fd_sc_hs__fa_2_13/a_484_347#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_15/a_1827_81# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_11/a_714_127#
+ fine_freq_track_1/sky130_fd_sc_hs__nor2b_1_35/a_27_112# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_55/a_1827_81#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_13/a_796_463# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_39/a_498_360#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_85/a_789_463# fine_freq_track_1/sky130_fd_sc_hs__a22oi_1_21/a_339_74#
+ fine_freq_track_1/sky130_fd_sc_hs__nand2_1_35/a_117_74# fine_freq_track_1/sky130_fd_sc_hs__o22ai_1_11/a_27_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_37/a_1547_508# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_37/a_706_463#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_27/a_834_355# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_27/a_319_360#
+ fine_freq_track_1/sky130_fd_sc_hs__xnor2_1_13/a_293_74# fine_freq_track_1/sky130_fd_sc_hs__dfstp_2_5/a_1596_118#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_41/a_494_366# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_11/Q_N
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_1/a_841_401# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_45/a_1434_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_5/a_1624_74# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_29/a_38_78#
+ fine_freq_track_1/sky130_fd_sc_hs__xnor2_1_5/a_112_119# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_15/a_832_118#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_11/a_1678_395# fine_freq_track_1/sky130_fd_sc_hs__a21oi_1_95/a_29_368#
+ fine_freq_track_1/sky130_fd_sc_hs__o21a_1_59/a_376_387# fine_freq_track_1/sky130_fd_sc_hs__dfxtp_2_1/a_1019_424#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_13/a_1465_471# fine_freq_track_1/sky130_fd_sc_hs__dfstp_2_1/a_398_74#
+ fine_freq_track_1/sky130_fd_sc_hs__fa_2_13/a_27_378# fine_freq_track_1/sky130_fd_sc_hs__fa_2_7/a_992_347#
+ fine_freq_track_1/sky130_fd_sc_hs__o21a_1_69/X fine_freq_track_1/sky130_fd_sc_hs__dfxtp_4_7/a_696_458#
+ fine_freq_track_1/sky130_fd_sc_hs__a22o_1_7/a_52_123# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_45/a_2010_409#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_89/a_37_78# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_17/a_37_78#
+ fine_freq_track_1/sky130_fd_sc_hs__nor2_1_25/a_116_368# fine_freq_track_1/sky130_fd_sc_hs__o21a_1_5/a_376_387#
+ fine_freq_track_1/sky130_fd_sc_hs__fa_2_7/a_487_79# fine_freq_track_1/sky130_fd_sc_hs__fa_2_17/SUM
+ fine_freq_track_1/sky130_fd_sc_hs__nor2b_1_7/a_278_368# fine_freq_track_1/sky130_fd_sc_hs__nor2_1_109/a_116_368#
+ fine_freq_track_1/sky130_fd_sc_hs__a22o_1_17/a_52_123# fine_freq_track_1/sky130_fd_sc_hs__maj3_1_1/a_406_384#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_25/a_841_401# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_3/a_706_463#
+ fine_freq_track_1/sky130_fd_sc_hs__dfxtp_4_7/a_1141_508# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_29/a_1624_74#
+ fine_freq_track_1/sky130_fd_sc_hs__fa_2_17/a_992_347# fine_freq_track_1/sky130_fd_sc_hs__nor2b_1_39/a_278_368#
+ fine_freq_track_1/sky130_fd_sc_hs__o21ai_1_7/a_27_74# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_21/a_1934_94#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_23/a_1598_93# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_27/a_812_138#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_43/a_38_78# fine_freq_track_1/sky130_fd_sc_hs__dfstp_2_7/a_716_456#
+ fine_freq_track_1/sky130_fd_sc_hs__fa_2_13/a_701_79# fine_freq_track_1/sky130_fd_sc_hs__a21oi_1_15/a_117_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_1/a_313_74# fine_freq_track_1/sky130_fd_sc_hs__fa_2_9/a_683_347#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_75/a_1627_493# fine_freq_track_1/sky130_fd_sc_hs__o22ai_1_3/a_340_368#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_49/a_1647_81# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_45/a_1736_119#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_45/a_1827_81# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_33/a_37_78#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_23/a_300_74# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_89/a_1647_81#
+ fine_freq_track_1/sky130_fd_sc_hs__nand4_1_3/a_259_74# fine_freq_track_1/sky130_fd_sc_hs__conb_1_3/HI
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_45/a_1266_119# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_65/a_313_74#
+ fine_freq_track_1/sky130_fd_sc_hs__xor2_1_7/a_355_368# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_1/a_789_463#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_65/a_1350_392# fine_freq_track_1/sky130_fd_sc_hs__nor3_1_13/a_114_368#
+ fine_freq_track_1/sky130_fd_sc_hs__sdlclkp_4_1/a_785_455# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_3/a_120_74#
+ fine_freq_track_1/sky130_fd_sc_hs__xnor2_1_13/a_112_119# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_75/a_789_463#
+ fine_freq_track_1/sky130_fd_sc_hs__o21a_1_39/a_83_244# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_17/a_319_360#
+ fine_freq_track_1/sky130_fd_sc_hs__dfxtp_2_1/a_644_504# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_61/a_1678_395#
+ fine_freq_track_1/sky130_fd_sc_hs__fa_2_19/a_683_347# fine_freq_track_1/sky130_fd_sc_hs__dfstp_2_4/a_1596_118#
+ fine_freq_track_1/sky130_fd_sc_hs__fa_2_23/a_1205_79# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_31/a_494_366#
+ fine_freq_track_1/sky130_fd_sc_hs__fa_2_21/a_1202_368# fine_freq_track_1/sky130_fd_sc_hs__nor2b_1_39/a_27_112#
+ fine_freq_track_1/sky130_fd_sc_hs__o21ai_1_9/a_162_368# fine_freq_track_1/sky130_fd_sc_hs__o21a_1_11/X
+ fine_freq_track_1/sky130_fd_sc_hs__a22oi_1_25/a_339_74# fine_freq_track_1/sky130_fd_sc_hs__nand2_1_39/a_117_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfsbp_2_1/a_398_74# fine_freq_track_1/sky130_fd_sc_hs__o21a_1_49/a_376_387#
+ fine_freq_track_1/sky130_fd_sc_hs__dfxtp_2_9/a_1217_314# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_49/a_890_138#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_29/a_1678_395# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_47/a_2026_424#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_89/a_890_138# fine_freq_track_1/sky130_fd_sc_hs__nand2_1_83/a_117_74#
+ fine_freq_track_1/sky130_fd_sc_hs__or2_1_1/a_152_368# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_23/a_910_118#
+ fine_freq_track_1/sky130_fd_sc_hs__nor2_1_15/a_116_368# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_3/a_1350_392#
+ fine_freq_track_1/sky130_fd_sc_hs__dfxtp_4_3/a_735_102# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_43/a_124_78#
+ fine_freq_track_1/sky130_fd_sc_hs__a21oi_1_99/a_29_368# fine_freq_track_1/sky130_fd_sc_hs__nor2_1_93/a_116_368#
+ fine_freq_track_1/sky130_fd_sc_hs__o21a_1_33/a_320_74# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_15/a_841_401#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_25/a_1550_119# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_19/a_1624_74#
+ fine_freq_track_1/sky130_fd_sc_hs__o31ai_1_3/a_203_368# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_11/a_1934_94#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_9/a_1736_119# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_1/a_1434_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_9/a_1266_119# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_73/a_1627_493#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_35/a_1827_81# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_13/a_507_368#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_79/a_1647_81# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_39/a_1224_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_9/a_37_78# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_25/a_789_463#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_73/a_1827_81# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_63/a_1350_392#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_33/a_796_463# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_65/a_789_463#
+ fine_freq_track_1/sky130_fd_sc_hs__dfstp_2_5/a_2022_94# fine_freq_track_1/sky130_fd_sc_hs__inv_2_9/Y
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_35/a_1547_508# fine_freq_track_1/sky130_fd_sc_hs__o22ai_1_3/a_142_368#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_23/a_1627_493# fine_freq_track_1/sky130_fd_sc_hs__a21oi_1_19/a_117_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfxtp_2_5/a_1172_124# fine_freq_track_1/sky130_fd_sc_hs__dfstp_2_1/a_1596_118#
+ fine_freq_track_1/sky130_fd_sc_hs__fa_2_13/a_1205_79# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_79/a_1678_395#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_85/a_834_355# fine_freq_track_1/sky130_fd_sc_hs__xor2_1_1/a_194_125#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_13/a_1350_392# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_69/a_313_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_25/a_1434_74# fine_freq_track_1/sky130_fd_sc_hs__a21oi_1_63/a_117_74#
+ fine_freq_track_1/sky130_fd_sc_hs__o21a_1_39/a_376_387# fine_freq_track_1/sky130_fd_sc_hs__dfsbp_2_1/a_1258_341#
+ fine_freq_track_1/sky130_fd_sc_hs__dfxtp_2_7/a_1217_314# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_15/a_33_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_35/a_832_118# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_9/a_714_127#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_79/a_890_138# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_1/a_38_78#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_43/a_2010_409# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_13/a_910_118#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_47/a_817_508# fine_freq_track_1/sky130_fd_sc_hs__fa_2_23/SUM
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_9/a_796_463# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_43/a_699_463#
+ fine_freq_track_1/sky130_fd_sc_hs__fa_2_11/a_487_79# fine_freq_track_1/sky130_fd_sc_hs__o21a_1_21/a_83_244#
+ fine_freq_track_1/sky130_fd_sc_hs__nor2_1_83/a_116_368# fine_freq_track_1/sky130_fd_sc_hs__a222oi_1_1/a_697_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfxtp_4_5/a_1141_508# fine_freq_track_1/sky130_fd_sc_hs__a22oi_1_13/a_159_74#
+ fine_freq_track_1/sky130_fd_sc_hs__nand2_1_87/a_117_74# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_47/a_1624_74#
+ fine_freq_track_1/sky130_fd_sc_hs__conb_1_3/a_21_290# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_41/a_1598_93#
+ fine_freq_track_1/sky130_fd_sc_hs__nand2b_1_1/a_269_74# fine_freq_track_1/sky130_fd_sc_hs__a22oi_1_5/a_339_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_7/a_1736_119# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_85/a_812_138#
+ fine_freq_track_1/sky130_fd_sc_hs__nand2_1_21/a_117_74# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_7/a_1266_119#
+ fine_freq_track_1/sky130_fd_sc_hs__xnor2_1_5/a_138_385# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_43/a_1736_119#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_91/a_124_78# fine_freq_track_1/sky130_fd_sc_hs__dfxtp_2_5/a_695_459#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_69/a_1647_81# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_43/a_1266_119#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_15/a_789_463# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_63/a_1827_81#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_27/a_37_78# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_43/a_507_368#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_55/a_789_463# fine_freq_track_1/sky130_fd_sc_hs__dfstp_2_4/a_767_384#
+ fine_freq_track_1/sky130_fd_sc_hs__inv_4_15/A fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_21/a_1627_493#
+ fine_freq_track_1/sky130_fd_sc_hs__dfxtp_2_3/a_1172_124# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_45/a_706_463#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_37/a_319_360# fine_freq_track_1/sky130_fd_sc_hs__a21oi_1_82/a_29_368#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_11/a_494_366# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_39/a_33_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_1/a_834_355# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_75/a_834_355#
+ fine_freq_track_1/sky130_fd_sc_hs__nand4_1_1/a_181_74# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_15/a_1434_74#
+ fine_freq_track_1/sky130_fd_sc_hs__o21a_1_29/a_376_387# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_31/a_1482_48#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_11/a_1465_471# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_27/a_1678_395#
+ fine_freq_track_1/sky130_fd_sc_hs__dfxtp_4_5/a_651_503# fine_freq_track_1/sky130_fd_sc_hs__maj3_1_3/a_595_136#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_45/a_2026_424# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_69/a_890_138#
+ fine_freq_track_1/sky130_fd_sc_hs__dfxtp_4_7/a_544_485# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_47/a_120_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_1/a_1350_392# fine_freq_track_1/sky130_fd_sc_hs__a21oi_1_67/a_117_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_15/a_120_74# fine_freq_track_1/sky130_fd_sc_hs__dfstp_2_4/a_781_74#
+ fine_freq_track_1/sky130_fd_sc_hs__a21oi_1_33/a_117_74# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_33/a_699_463#
+ fine_freq_track_1/sky130_fd_sc_hs__xnor2_1_13/a_138_385# fine_freq_track_1/sky130_fd_sc_hs__dfxtp_2_1/a_538_429#
+ fine_freq_track_1/sky130_fd_sc_hs__nand4_2_1/Y fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_23/a_1550_119#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_39/a_125_78# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_41/a_300_74#
+ fine_freq_track_1/sky130_fd_sc_hs__fa_2_1/a_484_347# fine_freq_track_1/sky130_fd_sc_hs__nor2_1_119/a_116_368#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_35/a_841_401# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_5/a_300_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_3/a_319_360# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_7/a_922_127#
+ fine_freq_track_1/sky130_fd_sc_hs__xnor2_1_3/a_376_368# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_13/Q_N
+ fine_freq_track_1/sky130_fd_sc_hs__o211ai_1_11/a_311_74# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_31/a_1598_93#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_51/a_313_74# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_13/a_856_304#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_1/a_812_138# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_75/a_812_138#
+ fine_freq_track_1/sky130_fd_sc_hs__o2bb2ai_1_1/a_490_368# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_13/a_850_127#
+ fine_freq_track_1/sky130_fd_sc_hs__o21a_1_25/a_83_244# fine_freq_track_1/sky130_fd_sc_hs__fa_2_11/a_484_347#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_41/a_1736_119# fine_freq_track_1/sky130_fd_sc_hs__fa_2_7/a_1119_79#
+ fine_freq_track_1/sky130_fd_sc_hs__a22oi_1_17/a_159_74# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_7/a_1482_48#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_59/a_1647_81# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_41/a_1266_119#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_53/a_1827_81# fine_freq_track_1/sky130_fd_sc_hs__a22o_1_21/a_230_79#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_33/a_507_368# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_5/a_817_508#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_45/a_789_463# fine_freq_track_1/sky130_fd_sc_hs__nor4_1_3/a_342_368#
+ fine_freq_track_1/sky130_fd_sc_hs__nand2b_1_5/a_269_74# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_33/a_1547_508#
+ fine_freq_track_1/sky130_fd_sc_hs__a222oi_1_1/a_119_74# fine_freq_track_1/sky130_fd_sc_hs__a22oi_1_11/a_339_74#
+ fine_freq_track_1/sky130_fd_sc_hs__nand2_1_25/a_117_74# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_25/a_834_355#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_17/a_124_78# fine_freq_track_1/sky130_fd_sc_hs__fa_2_17/a_1119_79#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_77/a_1678_395# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_65/a_834_355#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_9/a_1934_94# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_11/a_1350_392#
+ fine_freq_track_1/sky130_fd_sc_hs__o21a_1_19/a_376_387# fine_freq_track_1/sky130_fd_sc_hs__fa_2_11/a_27_79#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_21/a_1482_48# fine_freq_track_1/sky130_fd_sc_hs__nand2_1_15/Y
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_25/a_1678_395# fine_freq_track_1/sky130_fd_sc_hs__a21oi_1_85/a_29_368#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_59/a_890_138# fine_freq_track_1/sky130_fd_sc_hs__xnor2_1_11/a_376_368#
+ fine_freq_track_1/sky130_fd_sc_hs__nand4_1_5/a_181_74# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_41/a_2010_409#
+ fine_freq_track_1/sky130_fd_sc_hs__a22oi_1_3/a_71_368# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_29/a_1465_471#
+ fine_freq_track_1/sky130_fd_sc_hs__a21oi_1_51/a_29_368# fine_freq_track_1/sky130_fd_sc_hs__fa_2_5/a_336_347#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_27/a_817_508# fine_freq_track_1/sky130_fd_sc_hs__a211oi_4_1/a_92_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_33/a_910_118# fine_freq_track_1/sky130_fd_sc_hs__sdlclkp_1_1/a_288_48#
+ fine_freq_track_1/sky130_fd_sc_hs__a31oi_2_1/a_27_368# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_23/a_699_463#
+ fine_freq_track_1/sky130_fd_sc_hs__nor2_1_63/a_116_368# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_5/a_498_360#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_21/a_1550_119# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_11/a_37_78#
+ fine_freq_track_1/sky130_fd_sc_hs__a21oi_1_1/a_29_368# fine_freq_track_1/sky130_fd_sc_hs__a22o_1_25/a_132_392#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_1/a_706_463# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_27/a_1624_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_21/a_1598_93# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_25/a_812_138#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_65/a_812_138# fine_freq_track_1/sky130_fd_sc_hs__a21oi_1_37/a_117_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_43/a_856_304# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_71/a_1627_493#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_43/a_850_127# fine_freq_track_1/sky130_fd_sc_hs__o21ai_1_11/a_27_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_9/a_300_74# fine_freq_track_1/sky130_fd_sc_hs__a21oi_1_83/a_117_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_23/a_507_368# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_61/a_1350_392#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_35/a_789_463# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_55/a_313_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_29/a_498_360# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_83/a_1827_81#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_31/a_1547_508# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_41/a_796_463#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_73/a_789_463# fine_freq_track_1/sky130_fd_sc_hs__o21a_1_29/a_83_244#
+ fine_freq_track_1/sky130_fd_sc_hs__fa_2_19/a_487_79# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_9/a_910_118#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_21/a_313_74# fine_freq_track_1/sky130_fd_sc_hs__dfxtp_2_1/a_1172_124#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_25/a_706_463# fine_freq_track_1/sky130_fd_sc_hs__a222o_1_1/a_337_390#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_15/a_834_355# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_39/a_1627_493#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_55/a_834_355# fine_freq_track_1/sky130_fd_sc_hs__nor4_1_3/a_144_368#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_5/a_494_366# fine_freq_track_1/sky130_fd_sc_hs__o21a_1_73/a_83_244#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_91/a_2010_409# fine_freq_track_1/sky130_fd_sc_hs__maj3_1_3/a_223_120#
+ fine_freq_track_1/sky130_fd_sc_hs__nand2b_1_9/a_269_74# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_29/a_1350_392#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_35/a_1434_74# fine_freq_track_1/sky130_fd_sc_hs__a211oi_1_1/a_71_368#
+ fine_freq_track_1/sky130_fd_sc_hs__a22o_1_1/a_132_392# fine_freq_track_1/sky130_fd_sc_hs__dfxtp_2_5/a_1217_314#
+ fine_freq_track_1/sky130_fd_sc_hs__a22oi_1_15/a_339_74# fine_freq_track_1/sky130_fd_sc_hs__nand2_1_29/a_117_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_11/a_1482_48# fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_43/a_2026_424#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_43/a_832_118# fine_freq_track_1/sky130_fd_sc_hs__nor2b_1_41/a_27_112#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_27/a_1465_471# fine_freq_track_1/sky130_fd_sc_hs__nand2_1_73/a_117_74#
+ fine_freq_track_1/sky130_fd_sc_hs__a21oi_1_117/a_117_74# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_17/a_817_508#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_59/a_2010_409# fine_freq_track_1/sky130_fd_sc_hs__nor3_1_7/a_114_368#
+ fine_freq_track_1/sky130_fd_sc_hs__dfxtp_4_2/a_735_102# fine_freq_track_1/sky130_fd_sc_hs__dfstp_2_1/a_225_74#
+ fine_freq_track_1/sky130_fd_sc_hs__nand2_4_13/a_27_74# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_13/a_699_463#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_33/a_124_78# fine_freq_track_1/sky130_fd_sc_hs__nor2_1_53/a_116_368#
+ fine_freq_track_1/sky130_fd_sc_hs__o211ai_1_3/a_311_74# fine_freq_track_1/sky130_fd_sc_hs__a21oi_1_89/a_29_368#
+ fine_freq_track_1/sky130_fd_sc_hs__dfxtp_4_3/a_1141_508# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_49/a_33_74#
+ fine_freq_track_1/sky130_fd_sc_hs__o21a_1_23/a_320_74# fine_freq_track_1/sky130_fd_sc_hs__a22o_1_15/a_132_392#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_91/a_699_463# fine_freq_track_1/sky130_fd_sc_hs__dfxtp_2_11/a_431_508#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrbp_1_17/a_1624_74# fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_39/a_1550_119#
+ fine_freq_track_1/sky130_fd_sc_hs__a22oi_1_7/a_71_368# fine_freq_track_1/sky130_fd_sc_hs__nor2b_1_29/a_278_368#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_11/a_1598_93# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_15/a_812_138#
+ fine_freq_track_1/sky130_fd_sc_hs__nand2_1_1/a_117_74# fine_freq_track_1/sky130_fd_sc_hs__a21oi_1_23/a_29_368#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_5/a_1736_119# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_55/a_812_138#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_33/a_856_304# fine_freq_track_1/sky130_fd_sc_hs__maj3_1_3/a_84_74#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_5/a_1266_119# fine_freq_track_1/sky130_fd_sc_hs__nor4_1_3/a_228_368#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtn_1_33/a_850_127# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_51/a_37_78#
+ fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_39/a_1647_81# fine_freq_track_1/sky130_fd_sc_hs__xor2_1_1/a_455_87#
+ fine_freq_track_1/sky130_fd_sc_hs__a21oi_1_5/a_29_368# fine_freq_track_1/sky130_fd_sc_hs__dfrtp_4_89/a_1627_493#
+ fine_freq_track_1/sky130_fd_sc_hs__fa_2_1/a_1205_79# fine_freq_track
Xsky130_fd_sc_hs__clkbuf_16_90 DVSS: DVDD: DVDD: DVSS: prbs_generator_syn_19/inj_err
+ prbs_generator_syn_31/inj_err sky130_fd_sc_hs__clkbuf_16_91/a_114_74# sky130_fd_sc_hs__clkbuf_16
Xsky130_fd_sc_hs__buf_2_17 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__buf_2_17/A sky130_fd_sc_hs__buf_2_17/X
+ sky130_fd_sc_hs__buf_2_17/a_21_260# sky130_fd_sc_hs__buf_2
Xsky130_fd_sc_hs__buf_2_28 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__buf_2_31/A sky130_fd_sc_hs__buf_2_31/X
+ sky130_fd_sc_hs__buf_2_31/a_21_260# sky130_fd_sc_hs__buf_2
Xsky130_fd_sc_hs__buf_2_39 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__buf_2_39/A sky130_fd_sc_hs__buf_2_39/X
+ sky130_fd_sc_hs__buf_2_39/a_21_260# sky130_fd_sc_hs__buf_2
Xsky130_fd_sc_hs__o21bai_2_19 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__buf_2_77/A
+ sky130_fd_sc_hs__nand2_2_33/Y sky130_fd_sc_hs__dlrtp_1_79/D sky130_fd_sc_hs__buf_2_79/A
+ sky130_fd_sc_hs__o21bai_2_19/a_27_74# sky130_fd_sc_hs__o21bai_2_19/a_225_74# sky130_fd_sc_hs__o21bai_2_19/a_507_368#
+ sky130_fd_sc_hs__o21bai_2
Xsky130_fd_sc_hs__nand2_2_20 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__inv_4_25/A sky130_fd_sc_hs__nand2_2_21/B
+ sky130_fd_sc_hs__nand2_2_27/B sky130_fd_sc_hs__nand2_2_21/a_27_74# sky130_fd_sc_hs__nand2_2
Xsky130_fd_sc_hs__conb_1_206 DVSS: DVDD: DVDD: DVSS: prbs_generator_syn_19/eqn[31]
+ prbs_generator_syn_19/cke sky130_fd_sc_hs__conb_1_207/a_165_290# sky130_fd_sc_hs__conb_1_207/a_21_290#
+ sky130_fd_sc_hs__conb_1
Xsky130_fd_sc_hs__nand2_2_31 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__nand2_2_31/Y
+ sky130_fd_sc_hs__or4_2_1/C sky130_fd_sc_hs__or4_2_1/A sky130_fd_sc_hs__nand2_2_31/a_27_74#
+ sky130_fd_sc_hs__nand2_2
Xsky130_fd_sc_hs__conb_1_217 DVSS: DVDD: DVDD: DVSS: prbs_generator_syn_25/eqn[22]
+ prbs_generator_syn_25/eqn[20] sky130_fd_sc_hs__conb_1_217/a_165_290# sky130_fd_sc_hs__conb_1_217/a_21_290#
+ sky130_fd_sc_hs__conb_1
Xsky130_fd_sc_hs__conb_1_228 DVSS: DVDD: DVDD: DVSS: prbs_generator_syn_23/eqn[31]
+ prbs_generator_syn_23/cke sky130_fd_sc_hs__conb_1_229/a_165_290# sky130_fd_sc_hs__conb_1_229/a_21_290#
+ sky130_fd_sc_hs__conb_1
Xsky130_fd_sc_hs__conb_1_239 DVSS: DVDD: DVDD: DVSS: prbs_generator_syn_29/eqn[31]
+ prbs_generator_syn_29/cke sky130_fd_sc_hs__conb_1_239/a_165_290# sky130_fd_sc_hs__conb_1_239/a_21_290#
+ sky130_fd_sc_hs__conb_1
Xsky130_fd_sc_hs__o21bai_2_5 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__o21bai_2_5/A1
+ sky130_fd_sc_hs__nand2_2_3/B sky130_fd_sc_hs__dlrtp_1_55/D sky130_fd_sc_hs__buf_2_51/A
+ sky130_fd_sc_hs__o21bai_2_5/a_27_74# sky130_fd_sc_hs__o21bai_2_5/a_225_74# sky130_fd_sc_hs__o21bai_2_5/a_507_368#
+ sky130_fd_sc_hs__o21bai_2
Xsky130_fd_sc_hs__o21ai_2_10 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__inv_4_11/Y sky130_fd_sc_hs__nand2_2_3/B
+ sky130_fd_sc_hs__o21ai_2_55/A1 sky130_fd_sc_hs__o21ai_2_11/Y sky130_fd_sc_hs__o21ai_2_11/a_116_368#
+ sky130_fd_sc_hs__o21ai_2_11/a_27_74# sky130_fd_sc_hs__o21ai_2
Xsky130_fd_sc_hs__o21ai_2_21 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__inv_4_15/Y sky130_fd_sc_hs__or2b_4_5/X
+ sky130_fd_sc_hs__nand2_2_11/B sky130_fd_sc_hs__o21ai_2_21/Y sky130_fd_sc_hs__o21ai_2_21/a_116_368#
+ sky130_fd_sc_hs__o21ai_2_21/a_27_74# sky130_fd_sc_hs__o21ai_2
Xsky130_fd_sc_hs__o21ai_2_32 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__inv_4_19/Y sky130_fd_sc_hs__clkinv_4_7/Y
+ sky130_fd_sc_hs__o21ai_4_1/A1 sky130_fd_sc_hs__buf_2_89/A sky130_fd_sc_hs__o21ai_2_33/a_116_368#
+ sky130_fd_sc_hs__o21ai_2_33/a_27_74# sky130_fd_sc_hs__o21ai_2
Xsky130_fd_sc_hs__o21ai_2_43 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__inv_4_25/Y sky130_fd_sc_hs__or2b_2_3/A
+ sky130_fd_sc_hs__clkinv_4_7/Y sky130_fd_sc_hs__buf_2_129/A sky130_fd_sc_hs__o21ai_2_43/a_116_368#
+ sky130_fd_sc_hs__o21ai_2_43/a_27_74# sky130_fd_sc_hs__o21ai_2
Xsky130_fd_sc_hs__o21ai_2_54 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__inv_4_29/A sky130_fd_sc_hs__nand2_2_5/B
+ sky130_fd_sc_hs__o21ai_2_55/A1 sky130_fd_sc_hs__buf_2_149/A sky130_fd_sc_hs__o21ai_2_55/a_116_368#
+ sky130_fd_sc_hs__o21ai_2_55/a_27_74# sky130_fd_sc_hs__o21ai_2
Xsky130_fd_sc_hs__clkinv_4_13 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__o21bai_2_5/A1
+ sky130_fd_sc_hs__or4_2_1/C sky130_fd_sc_hs__clkinv_4
Xprbs_generator_syn_15 prbs_generator_syn_19/clk prbs_generator_syn_19/rst prbs_generator_syn_15/cke
+ sky130_fd_sc_hs__conb_1_145/LO sky130_fd_sc_hs__conb_1_145/LO sky130_fd_sc_hs__conb_1_145/HI
+ sky130_fd_sc_hs__conb_1_145/HI sky130_fd_sc_hs__conb_1_145/HI sky130_fd_sc_hs__conb_1_145/HI
+ sky130_fd_sc_hs__conb_1_145/HI sky130_fd_sc_hs__conb_1_145/LO sky130_fd_sc_hs__conb_1_145/LO
+ sky130_fd_sc_hs__conb_1_145/LO sky130_fd_sc_hs__conb_1_145/LO prbs_generator_syn_15/eqn[31]
+ sky130_fd_sc_hs__conb_1_147/HI prbs_generator_syn_17/eqn[13] sky130_fd_sc_hs__conb_1_147/HI
+ prbs_generator_syn_17/eqn[13] sky130_fd_sc_hs__conb_1_147/HI prbs_generator_syn_17/eqn[13]
+ prbs_generator_syn_15/eqn[1] prbs_generator_syn_15/eqn[2] prbs_generator_syn_15/eqn[2]
+ prbs_generator_syn_15/eqn[2] prbs_generator_syn_15/eqn[2] prbs_generator_syn_15/eqn[1]
+ sky130_fd_sc_hs__conb_1_151/HI sky130_fd_sc_hs__conb_1_151/LO sky130_fd_sc_hs__conb_1_151/LO
+ sky130_fd_sc_hs__conb_1_151/HI sky130_fd_sc_hs__conb_1_151/LO sky130_fd_sc_hs__conb_1_151/HI
+ sky130_fd_sc_hs__conb_1_151/LO sky130_fd_sc_hs__conb_1_151/HI prbs_generator_syn_15/eqn[31]
+ prbs_generator_syn_15/eqn[30] prbs_generator_syn_15/eqn[30] prbs_generator_syn_15/eqn[30]
+ prbs_generator_syn_15/eqn[30] prbs_generator_syn_15/eqn[30] prbs_generator_syn_15/eqn[30]
+ prbs_generator_syn_15/eqn[30] prbs_generator_syn_15/eqn[30] prbs_generator_syn_15/eqn[22]
+ prbs_generator_syn_15/eqn[22] prbs_generator_syn_15/eqn[20] prbs_generator_syn_15/eqn[22]
+ prbs_generator_syn_15/eqn[22] prbs_generator_syn_15/eqn[22] prbs_generator_syn_15/eqn[22]
+ prbs_generator_syn_15/eqn[22] prbs_generator_syn_15/eqn[22] prbs_generator_syn_15/eqn[13]
+ prbs_generator_syn_15/eqn[13] prbs_generator_syn_15/eqn[13] prbs_generator_syn_15/eqn[9]
+ prbs_generator_syn_15/eqn[9] prbs_generator_syn_15/eqn[9] prbs_generator_syn_15/eqn[9]
+ prbs_generator_syn_15/eqn[9] prbs_generator_syn_15/eqn[9] prbs_generator_syn_15/eqn[9]
+ prbs_generator_syn_15/eqn[9] prbs_generator_syn_15/eqn[2] prbs_generator_syn_15/eqn[1]
+ prbs_generator_syn_15/eqn[2] prbs_generator_syn_19/inj_err prbs_generator_syn_15/eqn[31]
+ prbs_generator_syn_15/eqn[31] hr_16t4_mux_top_1/din[1] DVSS: DVDD: prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_1/a_293_74#
+ prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_15/X prbs_generator_syn_15/sky130_fd_sc_hs__nand2_1_35/B
+ prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_51/Y prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_9/A
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_9/CLK prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_47/a_27_74#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_37/a_1226_296# prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_3/B
+ prbs_generator_syn_15/sky130_fd_sc_hs__nor2b_1_7/a_27_112# prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_29/B
+ prbs_generator_syn_15/sky130_fd_sc_hs__sdlclkp_2_1/a_580_74# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_1/a_1141_508#
+ prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_5/Y prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_41/a_230_79#
+ prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_61/a_138_385# prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_43/a_132_392#
+ prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_3/a_222_392# prbs_generator_syn_15/sky130_fd_sc_hs__nor2b_1_9/a_27_112#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_61/a_27_74# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_35/a_206_368#
+ prbs_generator_syn_15/sky130_fd_sc_hs__nand2_2_3/Y prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_25/B
+ prbs_generator_syn_15/sky130_fd_sc_hs__nand2_1_11/a_117_74# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_67/a_651_503#
+ prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_45/X prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_39/a_696_458#
+ prbs_generator_syn_15/sky130_fd_sc_hs__sdlclkp_2_1/a_1198_74# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_45/a_1034_424#
+ prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_17/a_222_392# prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_55/a_222_392#
+ prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_53/Y prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_35/A
+ prbs_generator_syn_15/m3_13600_1651# prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_59/a_52_123#
+ prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_5/a_293_74# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_35/a_1226_296#
+ prbs_generator_syn_15/sky130_fd_sc_hs__nand2_1_51/B prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_5/a_651_503#
+ prbs_generator_syn_15/sky130_fd_sc_hs__nand2_1_21/B prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_8/a_27_74#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_15/a_27_74# prbs_generator_syn_15/sky130_fd_sc_hs__and2b_2_1/X
+ prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_13/X prbs_generator_syn_15/sky130_fd_sc_hs__nand2_2_3/a_27_74#
+ prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_50/a_138_385# prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_33/a_132_392#
+ prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_1/a_376_368# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_25/a_206_368#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_35/a_437_503# prbs_generator_syn_15/sky130_fd_sc_hs__sdlclkp_2_1/a_708_451#
+ prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_45/a_230_79# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_29/a_696_458#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_32/a_27_74# prbs_generator_syn_15/sky130_fd_sc_hs__nor2b_1_4/Y
+ prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_59/a_293_74# prbs_generator_syn_15/sky130_fd_sc_hs__nand2_1_47/a_117_74#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_73/a_735_102# prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_21/a_112_119#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_23/a_1141_508# prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_25/a_293_74#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_7/Q prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_3/a_112_119#
+ prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_35/B prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_51/X
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_53/a_1178_124# prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_23/a_132_392#
+ prbs_generator_syn_15/sky130_fd_sc_hs__nand2_1_3/B prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_15/a_206_368#
+ prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_63/a_132_392# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_55/a_27_74#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_25/a_437_503# prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_41/a_52_123#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_47/a_651_503# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_73/a_1141_508#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_19/a_696_458# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_57/a_696_458#
+ prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_7/X prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_43/a_1034_424#
+ prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_55/A prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_11/a_112_119#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_21/a_1141_508# prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_35/a_222_392#
+ prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_49/a_230_79# prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_67/Y
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_71/a_27_74# prbs_generator_syn_15/sky130_fd_sc_hs__nand2_1_33/B
+ prbs_generator_syn_15/sky130_fd_sc_hs__conb_1_1/LO prbs_generator_syn_15/sky130_fd_sc_hs__nand2_1_19/a_117_74#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_51/a_1178_124# prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_33/X
+ prbs_generator_syn_15/sky130_fd_sc_hs__nand2_1_29/B prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_41/Y
+ prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_53/a_132_392# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_45/a_206_368#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_15/a_437_503# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_37/a_651_503#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_39/a_544_485# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_53/a_735_102#
+ prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_45/a_52_123# prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_1/B
+ prbs_generator_syn_15/sky130_fd_sc_hs__nand2_2_3/B prbs_generator_syn_15/sky130_fd_sc_hs__clkbuf_16_1/A
+ prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_21/X prbs_generator_syn_15/sky130_fd_sc_hs__nand2_1_25/B
+ prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_39/a_376_368# prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_63/X
+ prbs_generator_syn_15/m3_13600_3481# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_69/a_1178_124#
+ prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_21/a_138_385# prbs_generator_syn_15/sky130_fd_sc_hs__nor2b_1_8/Y
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_19/a_1178_124# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_49/a_27_74#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_45/a_437_503# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_27/a_651_503#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_71/a_1141_508# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_65/a_651_503#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_29/a_544_485# prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_3/a_138_385#
+ prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_55/X prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_43/a_735_102#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_41/a_1034_424# prbs_generator_syn_15/sky130_fd_sc_hs__nand2_1_9/B
+ prbs_generator_syn_15/sky130_fd_sc_hs__nor2b_1_9/Y prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_59/a_1034_424#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_39/a_1141_508# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_33/a_1226_296#
+ prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_49/a_52_123# prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_47/Y
+ prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_43/Y prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_4/a_651_503#
+ prbs_generator_syn_15/sky130_fd_sc_hs__nand2_1_49/B prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_19/A
+ prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_11/a_138_385# prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_5/X
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_63/a_206_368# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_17/a_651_503#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_19/a_544_485# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_55/a_651_503#
+ prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_9/Y prbs_generator_syn_15/sky130_fd_sc_hs__nand2_1_17/B
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_57/a_544_485# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_67/a_696_458#
+ prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_35/X prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_19/a_27_74#
+ prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_45/a_222_392# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_32/a_1226_296#
+ prbs_generator_syn_15/sky130_fd_sc_hs__nand2_1_43/B prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_25/A
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_1/a_206_368# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_49/a_1226_296#
+ prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_1/a_112_119# prbs_generator_syn_15/sky130_fd_sc_hs__or2_1_1/X
+ prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_59/a_376_368# prbs_generator_syn_15/sky130_fd_sc_hs__nand2_1_19/B
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_5/a_696_458# prbs_generator_syn_15/sky130_fd_sc_hs__nor2b_1_1/Y
+ prbs_generator_syn_15/sky130_fd_sc_hs__nor2b_1_5/a_278_368# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_17/a_1178_124#
+ prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_39/X prbs_generator_syn_15/m3_13600_5433#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_63/a_437_503# prbs_generator_syn_15/sky130_fd_sc_hs__nand2_2_5/B
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_23/a_735_102# prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_53/A
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_61/a_735_102# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_57/a_1034_424#
+ prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_63/B prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_37/a_1141_508#
+ prbs_generator_syn_15/sky130_fd_sc_hs__nand2_1_47/B prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_29/X
+ prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_65/Y prbs_generator_syn_15/m3_13600_4701#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_1/a_437_503# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_67/a_1178_124#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_9/a_735_102# prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_13/a_132_392#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_15/a_1178_124# prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_15/A
+ prbs_generator_syn_15/sky130_fd_sc_hs__nand2_1_1/B prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_43/B
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_35/a_651_503# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_8/D
+ prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_29/A prbs_generator_syn_15/sky130_fd_sc_hs__nand2_1_7/B
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_13/a_735_102# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_47/a_696_458#
+ prbs_generator_syn_15/sky130_fd_sc_hs__nand2_1_31/B prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_51/a_735_102#
+ prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_59/X prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_35/a_1141_508#
+ prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_25/a_222_392# prbs_generator_syn_15/sky130_fd_sc_hs__sdlclkp_2_1/a_288_48#
+ prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_55/B prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_17/B
+ prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_43/A prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_7/A
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_65/a_1178_124# prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_59/Y
+ prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_41/X prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_21/a_230_79#
+ prbs_generator_syn_15/sky130_fd_sc_hs__nand2_1_57/a_117_74# prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_1/a_222_392#
+ prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_19/B prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_35/a_293_74#
+ prbs_generator_syn_15/sky130_fd_sc_hs__nand2_1_23/a_117_74# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_73/a_206_368#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_25/a_651_503# prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_1/a_138_385#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_37/a_696_458# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_67/a_544_485#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_43/a_27_74# prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_9/X
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_55/a_1034_424# prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_39/a_112_119#
+ prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_15/a_222_392# prbs_generator_syn_15/sky130_fd_sc_hs__conb_1_1/HI
+ prbs_generator_syn_15/sky130_fd_sc_hs__nand2_1_23/B prbs_generator_syn_15/sky130_fd_sc_hs__nand2_1_53/B
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_9/a_1178_124# prbs_generator_syn_15/sky130_fd_sc_hs__nor2b_1_4/A
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_47/a_1226_296# prbs_generator_syn_15/m3_13600_11045#
+ prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_17/X prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_29/a_376_368#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_5/a_544_485# prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_3/X
+ prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_31/a_132_392# prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_61/A
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_15/a_651_503# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_73/a_437_503#
+ prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_25/a_230_79# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_27/a_696_458#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_65/a_696_458# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_33/a_735_102#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_71/a_735_102# prbs_generator_syn_15/m3_13600_7263#
+ prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_43/a_222_392# prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_50/Y
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_8/a_1178_124# prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_53/B
+ prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_19/a_376_368# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_63/a_1178_124#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_4/a_696_458# prbs_generator_syn_15/sky130_fd_sc_hs__nor2b_1_4/a_278_368#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_13/a_1178_124# prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_61/a_132_392#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_53/a_206_368# prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_21/a_52_123#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_45/a_651_503# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_17/a_696_458#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_47/a_544_485# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_55/a_696_458#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_21/a_735_102# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_37/a_27_74#
+ prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_61/B prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_61/X
+ prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_59/a_112_119# prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_31/A
+ prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_33/a_222_392# prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_29/a_230_79#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_45/a_1226_296# prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_9/a_132_392#
+ prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_5/A prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_57/Y
+ prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_31/X prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_51/a_27_74#
+ prbs_generator_syn_15/sky130_fd_sc_hs__nor2b_1_8/a_27_112# prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_47/a_376_368#
+ prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_53/a_293_74# prbs_generator_syn_15/sky130_fd_sc_hs__nand2_1_43/a_117_74#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_8/a_735_102# prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_21/a_293_74#
+ prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_39/a_138_385# prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_63/Y
+ prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_51/a_132_392# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_43/a_206_368#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_53/a_437_503# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_37/a_544_485#
+ prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_57/X prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_53/a_1034_424#
+ prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_25/a_52_123# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_33/a_1141_508#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_63/Q prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_23/a_222_392#
+ prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_63/a_222_392# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_7/a_1178_124#
+ prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_53/X prbs_generator_syn_15/sky130_fd_sc_hs__nand2_2_5/Y
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_61/a_1178_124# prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_1/a_230_79#
+ prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_43/a_230_79# prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_11/a_230_79#
+ prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_41/a_132_392# prbs_generator_syn_15/sky130_fd_sc_hs__nand2_1_13/a_117_74#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_43/a_437_503# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_27/a_544_485#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_63/a_651_503# prbs_generator_syn_15/sky130_fd_sc_hs__nand2_1_7/a_117_74#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_35/a_696_458# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_65/a_544_485#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_51/a_1034_424# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_41/a_735_102#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_32/a_1141_508# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_49/a_1141_508#
+ prbs_generator_syn_15/sky130_fd_sc_hs__nand2_1_55/B prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_53/a_222_392#
+ prbs_generator_syn_15/sky130_fd_sc_hs__sdlclkp_2_1/a_114_112# prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_9/a_293_74#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_43/a_1226_296# prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_29/a_52_123#
+ prbs_generator_syn_15/sky130_fd_sc_hs__nand2_1_37/B prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_1/a_651_503#
+ prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_27/a_376_368# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_4/a_544_485#
+ prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_67/a_376_368# prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_27/X
+ prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_1/X prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_59/a_138_385#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_29/a_1178_124# prbs_generator_syn_15/m3_13600_2871#
+ prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_5/a_230_79# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_23/a_206_368#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_61/a_206_368# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_17/a_544_485#
+ prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_15/a_230_79# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_25/a_696_458#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_55/a_544_485# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_32/a_735_102#
+ prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_29/a_293_74# prbs_generator_syn_15/sky130_fd_sc_hs__nand2_1_17/a_117_74#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_69/a_1034_424# prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_29/a_112_119#
+ prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_37/X prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_31/B
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_19/a_1034_424# prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_33/A
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_9/a_206_368# prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_57/a_376_368#
+ prbs_generator_syn_15/sky130_fd_sc_hs__sdlclkp_2_1/a_706_317# prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_11/B
+ prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_1/a_52_123# prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_39/B
+ prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_21/a_132_392# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_13/a_206_368#
+ prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_43/a_52_123# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_51/a_206_368#
+ prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_47/X prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_23/a_437_503#
+ prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_11/a_52_123# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_61/a_437_503#
+ prbs_generator_syn_15/sky130_fd_sc_hs__nor2b_1_7/Y prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_51/A
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_15/a_696_458# prbs_generator_syn_15/sky130_fd_sc_hs__nor2b_1_5/Y
+ prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_9/a_230_79# prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_25/X
+ prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_19/a_112_119# prbs_generator_syn_15/sky130_fd_sc_hs__nand2_1_45/B
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_5/a_1178_124# prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_19/a_230_79#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_41/a_1226_296# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_59/a_1226_296#
+ prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_63/a_230_79# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_51/Q
+ prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_7/a_132_392# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_9/a_437_503#
+ prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_46/a_376_368# prbs_generator_syn_15/sky130_fd_sc_hs__nand2_1_33/a_117_74#
+ prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_11/a_293_74# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_27/a_1178_124#
+ prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_11/a_132_392# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_13/a_437_503#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_51/a_437_503# prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_5/a_52_123#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_35/a_544_485# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_73/a_651_503#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_45/a_696_458# prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_15/a_52_123#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_47/a_1141_508# prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_47/a_112_119#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_4/a_1178_124# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_17/a_1034_424#
+ prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_23/B prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_37/a_376_368#
+ prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_15/B prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_7/Y
+ prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_29/a_138_385# prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_33/a_230_79#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_25/a_1178_124# prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_47/a_293_74#
+ prbs_generator_syn_15/sky130_fd_sc_hs__nand2_1_37/a_117_74# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_33/a_206_368#
+ prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_15/a_293_74# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_71/a_206_368#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_25/a_544_485# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_67/a_1034_424#
+ prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_13/a_222_392# prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_9/a_52_123#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_15/a_1034_424# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_57/a_1226_296#
+ prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_19/a_52_123# prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_23/X
+ prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_63/a_52_123# prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_19/a_138_385#
+ prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_9/a_376_368# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_21/a_206_368#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_33/a_437_503# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_71/a_437_503#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_53/a_651_503# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_15/a_544_485#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_63/a_696_458# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_65/a_1034_424#
+ prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_19/a_293_74# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_45/a_1141_508#
+ prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_27/a_112_119# prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_67/a_112_119#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_1/a_1178_124# prbs_generator_syn_15/sky130_fd_sc_hs__conb_1_1/a_21_290#
+ prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_63/a_293_74# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_8/a_206_368#
+ prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_17/a_376_368# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_63/a_27_74#
+ prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_21/A prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_55/a_376_368#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_1/a_696_458# prbs_generator_syn_15/sky130_fd_sc_hs__nor2b_1_1/a_278_368#
+ prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_47/a_138_385# prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_33/a_52_123#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_9/a_1034_424# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_21/a_437_503#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_1/a_27_74# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_43/a_651_503#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_1/Q prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_45/a_544_485#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_69/a_735_102# prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_57/a_112_119#
+ prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_31/a_222_392# prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_13/A
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_55/a_1226_296# prbs_generator_syn_15/sky130_fd_sc_hs__nand2_2_5/a_27_74#
+ prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_53/a_230_79# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_8/a_437_503#
+ prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_67/a_293_74# prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_33/a_293_74#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_7/a_735_102# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_23/a_1178_124#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_41/a_206_368# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_8/a_1034_424#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_63/a_1034_424# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_59/a_735_102#
+ prbs_generator_syn_15/sky130_fd_sc_hs__nand2_1_5/B prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_43/a_1141_508#
+ prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_46/a_112_119# prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_61/a_222_392#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_13/a_1034_424# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_73/a_1178_124#
+ prbs_generator_syn_15/sky130_fd_sc_hs__nand2_1_27/B prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_13/B
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_57/a_27_74# prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_57/a_230_79#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_21/a_1178_124# prbs_generator_syn_15/sky130_fd_sc_hs__nor2b_1_1/a_27_112#
+ prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_27/a_138_385# prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_23/a_230_79#
+ prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_67/a_138_385# prbs_generator_syn_15/sky130_fd_sc_hs__nand2_1_41/B
+ prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_9/a_222_392# prbs_generator_syn_15/sky130_fd_sc_hs__nand2_1_27/a_117_74#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_32/a_206_368# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_23/a_651_503#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_41/a_437_503# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_73/a_27_74#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_61/a_651_503# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_63/a_544_485#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_49/a_735_102# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_73/a_696_458#
+ prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_37/a_112_119# prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_51/a_222_392#
+ prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_43/X prbs_generator_syn_15/sky130_fd_sc_hs__nand2_2_1/B
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_9/a_651_503# prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_53/a_52_123#
+ prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_49/X prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_25/a_376_368#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_1/a_544_485# prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_65/a_376_368#
+ prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_57/a_138_385# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_27/a_27_74#
+ prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_39/a_132_392# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_7/a_1034_424#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_13/a_651_503# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_32/a_437_503#
+ prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_27/a_230_79# prbs_generator_syn_15/m3_13600_12265#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_51/a_651_503# prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_59/B
+ prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_47/A prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_61/a_1034_424#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_41/a_1141_508# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_59/a_1141_508#
+ prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_41/a_222_392# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_53/a_1226_296#
+ prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_3/A prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_71/a_1178_124#
+ prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_9/a_112_119# prbs_generator_syn_15/sky130_fd_sc_hs__nand2_1_3/a_117_74#
+ prbs_generator_syn_15/m3_13600_8483# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_39/a_1178_124#
+ prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_57/a_52_123# prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_46/a_138_385#
+ prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_23/a_52_123# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_67/a_27_74#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_53/a_696_458# prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_17/a_112_119#
+ prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_11/A prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_55/a_112_119#
+ prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_1/A prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_51/a_1226_296#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_29/a_1034_424# prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_59/A
+ prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_23/A prbs_generator_syn_15/sky130_fd_sc_hs__nand2_1_39/B
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_5/a_27_74# prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_57/a_293_74#
+ prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_37/a_138_385# prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_59/a_132_392#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_33/a_651_503# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_71/a_651_503#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_43/a_696_458# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_73/a_544_485#
+ prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_27/a_52_123# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_57/a_1141_508#
+ prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_21/a_222_392# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_35/a_27_74#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_69/a_1226_296# prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_37/B
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_19/a_1226_296# prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_35/a_376_368#
+ prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_47/a_230_79# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_37/a_1178_124#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_5/a_1034_424# prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_49/a_132_392#
+ prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_7/a_222_392# prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_27/a_293_74#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_21/a_651_503# prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_9/a_138_385#
+ prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_11/a_222_392# prbs_generator_syn_15/m3_13600_14095#
+ prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_50/A prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_27/a_1034_424#
+ prbs_generator_syn_15/sky130_fd_sc_hs__nand2_1_13/B prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_8/a_651_503#
+ prbs_generator_syn_15/m3_13600_9703# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_35/a_1178_124#
+ prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_17/a_138_385# prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_55/a_138_385#
+ prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_7/a_230_79# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_4/a_1034_424#
+ prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_7/a_376_368# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_69/a_206_368#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_23/a_696_458# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_53/a_544_485#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_39/a_735_102# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_61/a_696_458#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_55/a_1141_508# prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_25/a_112_119#
+ prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_65/a_112_119# prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_43/a_293_74#
+ prbs_generator_syn_15/sky130_fd_sc_hs__nand2_1_57/B prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_25/a_1034_424#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_7/a_206_368# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_17/a_1226_296#
+ prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_15/a_376_368# prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_53/a_376_368#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_9/a_696_458# prbs_generator_syn_15/m3_13600_431#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_45/a_27_74# prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_47/a_52_123#
+ prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_29/a_132_392# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_59/a_206_368#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_69/a_437_503# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_41/a_651_503#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_43/a_544_485# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_13/a_696_458#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_29/a_735_102# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_51/a_696_458#
+ prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_61/Y prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_67/a_1226_296#
+ prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_5/a_132_392# prbs_generator_syn_15/sky130_fd_sc_hs__and2b_2_1/a_198_48#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_7/a_437_503# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_15/a_1226_296#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_69/a_27_74# prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_46/a_293_74#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_1/a_1034_424# prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_19/a_132_392#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_49/a_206_368# prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_7/a_52_123#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_59/a_437_503# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_32/a_651_503#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_7/a_27_74# prbs_generator_syn_15/sky130_fd_sc_hs__nand2_2_1/a_27_74#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_19/a_735_102# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_57/a_735_102#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_65/a_1226_296# prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_37/A
+ prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_33/a_376_368# prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_37/a_230_79#
+ prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_25/a_138_385# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_39/a_27_74#
+ prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_65/a_138_385# prbs_generator_syn_15/sky130_fd_sc_hs__nor2b_1_9/a_278_368#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_49/a_437_503# prbs_generator_syn_15/sky130_fd_sc_hs__and2b_2_1/a_505_74#
+ prbs_generator_syn_15/sky130_fd_sc_hs__nand2_1_51/a_117_74# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_23/a_544_485#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_33/a_696_458# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_61/a_544_485#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_9/a_1226_296# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_53/a_1141_508#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_71/a_696_458# prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_35/a_112_119#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_23/a_1034_424# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_9/a_544_485#
+ prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_63/a_376_368# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_33/a_1178_124#
+ prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_5/a_376_368# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_13/a_544_485#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_73/a_1034_424# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_21/a_696_458#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_51/a_544_485# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_8/a_1226_296#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_51/a_1141_508# prbs_generator_syn_15/sky130_fd_sc_hs__nand2_1_55/a_117_74#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_21/a_1034_424# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_63/a_1226_296#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_23/a_27_74# prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_7/a_112_119#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_13/a_1226_296# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_8/a_696_458#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_32/a_1178_124# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_49/a_1178_124#
+ prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_37/a_52_123# prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_27/a_132_392#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_71/Q prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_67/a_735_102#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_69/a_1141_508# prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_15/a_112_119#
+ prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_53/a_112_119# prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_39/a_222_392#
+ prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_55/a_230_79# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_19/a_1141_508#
+ prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_37/a_293_74# prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_43/a_376_368#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_5/a_735_102# prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_35/a_138_385#
+ prbs_generator_syn_15/sky130_fd_sc_hs__sdlclkp_2_1/a_114_424# prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_57/a_132_392#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_71/a_1034_424# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_7/a_1226_296#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_33/a_544_485# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_41/a_696_458#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_71/a_544_485# prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_21/B
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_61/a_1226_296# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_39/a_1034_424#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_17/a_27_74# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_9/a_27_74#
+ prbs_generator_syn_15/sky130_fd_sc_hs__nor2b_1_5/a_27_112# prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_47/a_132_392#
+ prbs_generator_syn_15/sky130_fd_sc_hs__nor2b_1_8/a_278_368# prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_9/B
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_39/a_206_368# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_33/a_27_74#
+ prbs_generator_syn_15/sky130_fd_sc_hs__nand2_1_41/a_117_74# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_69/a_651_503#
+ prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_51/a_293_74# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_21/a_544_485#
+ prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_7/a_138_385# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_32/a_696_458#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_47/a_735_102# prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_33/a_112_119#
+ prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_59/a_222_392# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_17/a_1141_508#
+ prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_55/a_52_123# prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_3/a_293_74#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_7/a_651_503# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_29/a_1226_296#
+ prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_23/a_376_368# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_8/a_544_485#
+ prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_47/B prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_47/a_1178_124#
+ prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_15/a_138_385# prbs_generator_syn_15/sky130_fd_sc_hs__sdlclkp_2_1/a_1195_374#
+ prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_53/a_138_385# prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_37/a_132_392#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_29/a_206_368# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_39/a_437_503#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_59/a_651_503# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_37/a_735_102#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_67/a_1141_508# prbs_generator_syn_15/sky130_fd_sc_hs__and2b_2_1/a_27_74#
+ prbs_generator_syn_15/sky130_fd_sc_hs__conb_1_1/a_165_290# prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_55/a_293_74#
+ prbs_generator_syn_15/sky130_fd_sc_hs__nand2_1_45/a_117_74# prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_63/a_112_119#
+ prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_49/a_222_392# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_37/a_1034_424#
+ prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_23/a_293_74# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_15/a_1141_508#
+ prbs_generator_syn_15/sky130_fd_sc_hs__nand2_1_5/a_117_74# prbs_generator_syn_15/m3_13600_13485#
+ prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_5/a_112_119# prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_13/a_376_368#
+ prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_51/a_376_368# prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_7/a_293_74#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_19/a_206_368# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_57/a_206_368#
+ prbs_generator_syn_15/sky130_fd_sc_hs__sdlclkp_2_1/a_318_74# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_29/a_437_503#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_49/a_651_503# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_25/a_27_74#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_5/a_1226_296# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_41/a_544_485#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_27/a_735_102# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_65/a_1141_508#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_65/a_735_102# prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_3/a_230_79#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_35/a_1034_424# prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_13/a_230_79#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_41/a_27_74# prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_3/a_132_392#
+ prbs_generator_syn_15/sky130_fd_sc_hs__nand2_1_49/a_117_74# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_27/a_1226_296#
+ prbs_generator_syn_15/sky130_fd_sc_hs__nand2_1_15/a_117_74# prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_41/a_376_368#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_45/a_1178_124# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_4/a_735_102#
+ prbs_generator_syn_15/sky130_fd_sc_hs__nand2_1_9/a_117_74# prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_33/a_138_385#
+ prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_17/a_132_392# prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_55/a_132_392#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_9/a_1141_508# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_19/a_437_503#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_57/a_437_503# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_4/a_1226_296#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_32/a_544_485# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_17/a_735_102#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_55/a_735_102# prbs_generator_syn_15/m3_13600_2261#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_65/a_27_74# prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_29/a_222_392#
+ prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_43/a_112_119# prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_19/X
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_25/a_1226_296# prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_31/a_376_368#
+ prbs_generator_syn_15/sky130_fd_sc_hs__or2_1_1/a_63_368# prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_17/a_230_79#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_4/a_27_74# prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_61/a_230_79#
+ prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_63/a_138_385# prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_5/a_222_392#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_8/a_1141_508# prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_41/a_293_74#
+ prbs_generator_syn_15/sky130_fd_sc_hs__nand2_1_31/a_117_74# prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_5/a_138_385#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_63/a_1141_508# prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_19/a_222_392#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_13/a_1141_508# prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_3/a_52_123#
+ prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_13/a_52_123# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_43/a_1178_124#
+ prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_61/a_376_368# prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_35/a_132_392#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_67/a_206_368# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_1/a_1226_296#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_69/a_696_458# prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_31/a_230_79#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_35/a_735_102# prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_23/a_112_119#
+ prbs_generator_syn_15/sky130_fd_sc_hs__nand2_1_35/a_117_74# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_59/a_27_74#
+ prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_13/a_293_74# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_5/a_206_368#
+ prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_50/a_376_368# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_7/a_696_458#
+ prbs_generator_syn_15/sky130_fd_sc_hs__nor2b_1_7/a_278_368# prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_17/a_52_123#
+ prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_43/a_138_385# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_7/a_1141_508#
+ prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_61/a_52_123# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_67/a_437_503#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_61/a_1141_508# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_25/a_735_102#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_59/a_696_458# prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_13/a_112_119#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_33/a_1034_424# prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_51/a_112_119#
+ prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_35/a_230_79# prbs_generator_syn_15/m3_13600_4091#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_23/a_1226_296# prbs_generator_syn_15/sky130_fd_sc_hs__nand2_1_39/a_117_74#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_29/a_27_74# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_5/a_437_503#
+ prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_17/a_293_74# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_41/a_1178_124#
+ prbs_generator_syn_15/sky130_fd_sc_hs__or2_1_1/a_152_368# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_59/a_1178_124#
+ prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_61/a_293_74# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_47/a_206_368#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_39/a_651_503# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_49/a_696_458#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_15/a_735_102# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_32/a_1034_424#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_73/a_1226_296# prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_27/a_222_392#
+ prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_41/a_112_119# prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_31/a_52_123#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_49/a_1034_424# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_29/a_1141_508#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_21/a_1226_296# prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_39/a_230_79#
+ prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_23/a_138_385# prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_51/a_230_79#
+ prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_45/a_132_392# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_37/a_206_368#
+ prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_65/a_293_74# prbs_generator_syn_15/sky130_fd_sc_hs__nand2_1_53/a_117_74#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_47/a_437_503# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_29/a_651_503#
+ prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_31/a_293_74# prbs_generator_syn_15/sky130_fd_sc_hs__nand2_1_21/a_117_74#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_69/a_544_485# prbs_generator_syn_15/sky130_fd_sc_hs__clkbuf_16_1/a_114_74#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_45/a_735_102# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_13/a_27_74#
+ prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_31/a_112_119# prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_57/a_222_392#
+ prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_35/a_52_123# prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_21/a_376_368#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_7/a_544_485# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_57/a_1178_124#
+ prbs_generator_syn_15/m3_13600_6043# prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_13/a_138_385#
+ prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_51/a_138_385# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_5/a_1141_508#
+ prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_3/a_376_368# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_27/a_206_368#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_65/a_206_368# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_37/a_437_503#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_19/a_651_503# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_57/a_651_503#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_59/a_544_485# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_71/a_1226_296#
+ prbs_generator_syn_15/sky130_fd_sc_hs__nand2_1_25/a_117_74# prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_61/a_112_119#
+ prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_47/a_222_392# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_27/a_1141_508#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_53/a_27_74# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_4/a_206_368#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_39/a_1226_296# prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_11/a_376_368#
+ prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_39/a_52_123# prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_41/a_138_385#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_4/a_1141_508# prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_25/a_132_392#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_17/a_206_368# prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_41/A
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_55/a_206_368# prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_51/a_52_123#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_27/a_437_503# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_65/a_437_503#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_49/a_544_485# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_63/a_735_102#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_47/a_1034_424# prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_50/a_112_119#
+ prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_37/a_222_392# prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_59/a_230_79#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_25/a_1141_508# prbs_generator_syn_15/sky130_fd_sc_hs__nor2b_1_4/a_27_112#
+ prbs_generator_syn_15/sky130_fd_sc_hs__sdlclkp_2_1/a_685_81# prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_1/a_132_392#
+ prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_39/a_293_74# prbs_generator_syn_15/sky130_fd_sc_hs__nand2_1_29/a_117_74#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_4/a_437_503# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_55/a_1178_124#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_21/a_27_74# prbs_generator_syn_15/m3_13600_12875#
+ prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_50/a_293_74# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_1/a_735_102#
+ prbs_generator_syn_15/sky130_fd_sc_hs__xnor2_1_31/a_138_385# prbs_generator_syn_15/sky130_fd_sc_hs__a22o_1_15/a_132_392#
+ prbs_generator_syn_15/sky130_fd_sc_hs__nand2_1_1/a_117_74# prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_17/a_437_503#
+ prbs_generator_syn_15/sky130_fd_sc_hs__dfxtp_4_55/a_437_503# prbs_generator_syn
Xprbs_generator_syn_26 prbs_generator_syn_31/clk prbs_generator_syn_27/rst prbs_generator_syn_27/cke
+ sky130_fd_sc_hs__conb_1_257/LO sky130_fd_sc_hs__conb_1_257/LO sky130_fd_sc_hs__conb_1_257/LO
+ sky130_fd_sc_hs__conb_1_257/LO sky130_fd_sc_hs__conb_1_257/LO sky130_fd_sc_hs__conb_1_257/HI
+ sky130_fd_sc_hs__conb_1_257/HI sky130_fd_sc_hs__conb_1_257/HI sky130_fd_sc_hs__conb_1_257/HI
+ sky130_fd_sc_hs__conb_1_257/HI sky130_fd_sc_hs__conb_1_257/HI prbs_generator_syn_27/cke
+ prbs_generator_syn_27/cke prbs_generator_syn_27/cke prbs_generator_syn_27/cke prbs_generator_syn_27/cke
+ prbs_generator_syn_27/eqn[31] prbs_generator_syn_27/cke prbs_generator_syn_31/eqn[9]
+ prbs_generator_syn_31/eqn[20] prbs_generator_syn_31/eqn[21] prbs_generator_syn_31/eqn[20]
+ prbs_generator_syn_31/eqn[21] sky130_fd_sc_hs__conb_1_247/HI prbs_generator_syn_31/eqn[28]
+ sky130_fd_sc_hs__conb_1_247/HI sky130_fd_sc_hs__conb_1_247/HI prbs_generator_syn_31/eqn[30]
+ prbs_generator_syn_31/eqn[30] sky130_fd_sc_hs__conb_1_259/HI sky130_fd_sc_hs__conb_1_259/HI
+ prbs_generator_syn_31/eqn[30] prbs_generator_syn_27/eqn[31] prbs_generator_syn_27/eqn[30]
+ prbs_generator_syn_27/eqn[30] prbs_generator_syn_27/eqn[28] prbs_generator_syn_27/eqn[28]
+ prbs_generator_syn_27/eqn[28] prbs_generator_syn_27/eqn[28] prbs_generator_syn_27/eqn[28]
+ prbs_generator_syn_27/eqn[28] prbs_generator_syn_27/eqn[22] prbs_generator_syn_27/eqn[22]
+ prbs_generator_syn_27/eqn[20] prbs_generator_syn_27/eqn[22] prbs_generator_syn_27/eqn[22]
+ prbs_generator_syn_27/eqn[22] prbs_generator_syn_27/eqn[22] prbs_generator_syn_27/eqn[22]
+ prbs_generator_syn_27/eqn[9] prbs_generator_syn_27/eqn[9] prbs_generator_syn_27/eqn[9]
+ prbs_generator_syn_27/eqn[9] prbs_generator_syn_27/eqn[9] prbs_generator_syn_27/eqn[9]
+ prbs_generator_syn_27/eqn[8] prbs_generator_syn_27/eqn[8] prbs_generator_syn_27/eqn[8]
+ prbs_generator_syn_27/eqn[8] prbs_generator_syn_27/eqn[8] prbs_generator_syn_27/eqn[8]
+ prbs_generator_syn_27/eqn[8] prbs_generator_syn_27/eqn[1] prbs_generator_syn_31/eqn[9]
+ prbs_generator_syn_27/inj_err prbs_generator_syn_27/eqn[31] prbs_generator_syn_27/eqn[31]
+ hr_16t4_mux_top_1/din[4] DVSS: DVDD: prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_1/a_293_74#
+ prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_15/X prbs_generator_syn_27/sky130_fd_sc_hs__nand2_1_35/B
+ prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_51/Y prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_9/A
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_9/CLK prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_47/a_27_74#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_37/a_1226_296# prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_3/B
+ prbs_generator_syn_27/sky130_fd_sc_hs__nor2b_1_7/a_27_112# prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_29/B
+ prbs_generator_syn_27/sky130_fd_sc_hs__sdlclkp_2_1/a_580_74# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_1/a_1141_508#
+ prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_5/Y prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_41/a_230_79#
+ prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_61/a_138_385# prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_43/a_132_392#
+ prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_3/a_222_392# prbs_generator_syn_27/sky130_fd_sc_hs__nor2b_1_9/a_27_112#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_61/a_27_74# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_35/a_206_368#
+ prbs_generator_syn_27/sky130_fd_sc_hs__nand2_2_3/Y prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_25/B
+ prbs_generator_syn_27/sky130_fd_sc_hs__nand2_1_11/a_117_74# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_67/a_651_503#
+ prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_45/X prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_39/a_696_458#
+ prbs_generator_syn_27/sky130_fd_sc_hs__sdlclkp_2_1/a_1198_74# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_45/a_1034_424#
+ prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_17/a_222_392# prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_55/a_222_392#
+ prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_53/Y prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_35/A
+ prbs_generator_syn_27/m3_13600_1651# prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_59/a_52_123#
+ prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_5/a_293_74# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_35/a_1226_296#
+ prbs_generator_syn_27/sky130_fd_sc_hs__nand2_1_51/B prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_5/a_651_503#
+ prbs_generator_syn_27/sky130_fd_sc_hs__nand2_1_21/B prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_8/a_27_74#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_15/a_27_74# prbs_generator_syn_27/sky130_fd_sc_hs__and2b_2_1/X
+ prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_13/X prbs_generator_syn_27/sky130_fd_sc_hs__nand2_2_3/a_27_74#
+ prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_50/a_138_385# prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_33/a_132_392#
+ prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_1/a_376_368# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_25/a_206_368#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_35/a_437_503# prbs_generator_syn_27/sky130_fd_sc_hs__sdlclkp_2_1/a_708_451#
+ prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_45/a_230_79# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_29/a_696_458#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_32/a_27_74# prbs_generator_syn_27/sky130_fd_sc_hs__nor2b_1_4/Y
+ prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_59/a_293_74# prbs_generator_syn_27/sky130_fd_sc_hs__nand2_1_47/a_117_74#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_73/a_735_102# prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_21/a_112_119#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_23/a_1141_508# prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_25/a_293_74#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_7/Q prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_3/a_112_119#
+ prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_35/B prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_51/X
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_53/a_1178_124# prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_23/a_132_392#
+ prbs_generator_syn_27/sky130_fd_sc_hs__nand2_1_3/B prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_15/a_206_368#
+ prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_63/a_132_392# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_55/a_27_74#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_25/a_437_503# prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_41/a_52_123#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_47/a_651_503# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_73/a_1141_508#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_19/a_696_458# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_57/a_696_458#
+ prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_7/X prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_43/a_1034_424#
+ prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_55/A prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_11/a_112_119#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_21/a_1141_508# prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_35/a_222_392#
+ prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_49/a_230_79# prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_67/Y
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_71/a_27_74# prbs_generator_syn_27/sky130_fd_sc_hs__nand2_1_33/B
+ prbs_generator_syn_27/sky130_fd_sc_hs__conb_1_1/LO prbs_generator_syn_27/sky130_fd_sc_hs__nand2_1_19/a_117_74#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_51/a_1178_124# prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_33/X
+ prbs_generator_syn_27/sky130_fd_sc_hs__nand2_1_29/B prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_41/Y
+ prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_53/a_132_392# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_45/a_206_368#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_15/a_437_503# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_37/a_651_503#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_39/a_544_485# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_53/a_735_102#
+ prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_45/a_52_123# prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_1/B
+ prbs_generator_syn_27/sky130_fd_sc_hs__nand2_2_3/B prbs_generator_syn_27/sky130_fd_sc_hs__clkbuf_16_1/A
+ prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_21/X prbs_generator_syn_27/sky130_fd_sc_hs__nand2_1_25/B
+ prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_39/a_376_368# prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_63/X
+ prbs_generator_syn_27/m3_13600_3481# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_69/a_1178_124#
+ prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_21/a_138_385# prbs_generator_syn_27/sky130_fd_sc_hs__nor2b_1_8/Y
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_19/a_1178_124# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_49/a_27_74#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_45/a_437_503# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_27/a_651_503#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_71/a_1141_508# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_65/a_651_503#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_29/a_544_485# prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_3/a_138_385#
+ prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_55/X prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_43/a_735_102#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_41/a_1034_424# prbs_generator_syn_27/sky130_fd_sc_hs__nand2_1_9/B
+ prbs_generator_syn_27/sky130_fd_sc_hs__nor2b_1_9/Y prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_59/a_1034_424#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_39/a_1141_508# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_33/a_1226_296#
+ prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_49/a_52_123# prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_47/Y
+ prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_43/Y prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_4/a_651_503#
+ prbs_generator_syn_27/sky130_fd_sc_hs__nand2_1_49/B prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_19/A
+ prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_11/a_138_385# prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_5/X
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_63/a_206_368# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_17/a_651_503#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_19/a_544_485# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_55/a_651_503#
+ prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_9/Y prbs_generator_syn_27/sky130_fd_sc_hs__nand2_1_17/B
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_57/a_544_485# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_67/a_696_458#
+ prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_35/X prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_19/a_27_74#
+ prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_45/a_222_392# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_32/a_1226_296#
+ prbs_generator_syn_27/sky130_fd_sc_hs__nand2_1_43/B prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_25/A
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_1/a_206_368# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_49/a_1226_296#
+ prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_1/a_112_119# prbs_generator_syn_27/sky130_fd_sc_hs__or2_1_1/X
+ prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_59/a_376_368# prbs_generator_syn_27/sky130_fd_sc_hs__nand2_1_19/B
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_5/a_696_458# prbs_generator_syn_27/sky130_fd_sc_hs__nor2b_1_1/Y
+ prbs_generator_syn_27/sky130_fd_sc_hs__nor2b_1_5/a_278_368# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_17/a_1178_124#
+ prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_39/X prbs_generator_syn_27/m3_13600_5433#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_63/a_437_503# prbs_generator_syn_27/sky130_fd_sc_hs__nand2_2_5/B
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_23/a_735_102# prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_53/A
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_61/a_735_102# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_57/a_1034_424#
+ prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_63/B prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_37/a_1141_508#
+ prbs_generator_syn_27/sky130_fd_sc_hs__nand2_1_47/B prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_29/X
+ prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_65/Y prbs_generator_syn_27/m3_13600_4701#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_1/a_437_503# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_67/a_1178_124#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_9/a_735_102# prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_13/a_132_392#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_15/a_1178_124# prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_15/A
+ prbs_generator_syn_27/sky130_fd_sc_hs__nand2_1_1/B prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_43/B
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_35/a_651_503# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_8/D
+ prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_29/A prbs_generator_syn_27/sky130_fd_sc_hs__nand2_1_7/B
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_13/a_735_102# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_47/a_696_458#
+ prbs_generator_syn_27/sky130_fd_sc_hs__nand2_1_31/B prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_51/a_735_102#
+ prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_59/X prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_35/a_1141_508#
+ prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_25/a_222_392# prbs_generator_syn_27/sky130_fd_sc_hs__sdlclkp_2_1/a_288_48#
+ prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_55/B prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_17/B
+ prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_43/A prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_7/A
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_65/a_1178_124# prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_59/Y
+ prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_41/X prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_21/a_230_79#
+ prbs_generator_syn_27/sky130_fd_sc_hs__nand2_1_57/a_117_74# prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_1/a_222_392#
+ prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_19/B prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_35/a_293_74#
+ prbs_generator_syn_27/sky130_fd_sc_hs__nand2_1_23/a_117_74# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_73/a_206_368#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_25/a_651_503# prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_1/a_138_385#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_37/a_696_458# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_67/a_544_485#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_43/a_27_74# prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_9/X
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_55/a_1034_424# prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_39/a_112_119#
+ prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_15/a_222_392# prbs_generator_syn_27/sky130_fd_sc_hs__conb_1_1/HI
+ prbs_generator_syn_27/sky130_fd_sc_hs__nand2_1_23/B prbs_generator_syn_27/sky130_fd_sc_hs__nand2_1_53/B
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_9/a_1178_124# prbs_generator_syn_27/sky130_fd_sc_hs__nor2b_1_4/A
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_47/a_1226_296# prbs_generator_syn_27/m3_13600_11045#
+ prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_17/X prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_29/a_376_368#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_5/a_544_485# prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_3/X
+ prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_31/a_132_392# prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_61/A
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_15/a_651_503# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_73/a_437_503#
+ prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_25/a_230_79# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_27/a_696_458#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_65/a_696_458# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_33/a_735_102#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_71/a_735_102# prbs_generator_syn_27/m3_13600_7263#
+ prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_43/a_222_392# prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_50/Y
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_8/a_1178_124# prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_53/B
+ prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_19/a_376_368# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_63/a_1178_124#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_4/a_696_458# prbs_generator_syn_27/sky130_fd_sc_hs__nor2b_1_4/a_278_368#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_13/a_1178_124# prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_61/a_132_392#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_53/a_206_368# prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_21/a_52_123#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_45/a_651_503# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_17/a_696_458#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_47/a_544_485# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_55/a_696_458#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_21/a_735_102# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_37/a_27_74#
+ prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_61/B prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_61/X
+ prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_59/a_112_119# prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_31/A
+ prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_33/a_222_392# prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_29/a_230_79#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_45/a_1226_296# prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_9/a_132_392#
+ prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_5/A prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_57/Y
+ prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_31/X prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_51/a_27_74#
+ prbs_generator_syn_27/sky130_fd_sc_hs__nor2b_1_8/a_27_112# prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_47/a_376_368#
+ prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_53/a_293_74# prbs_generator_syn_27/sky130_fd_sc_hs__nand2_1_43/a_117_74#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_8/a_735_102# prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_21/a_293_74#
+ prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_39/a_138_385# prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_63/Y
+ prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_51/a_132_392# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_43/a_206_368#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_53/a_437_503# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_37/a_544_485#
+ prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_57/X prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_53/a_1034_424#
+ prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_25/a_52_123# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_33/a_1141_508#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_63/Q prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_23/a_222_392#
+ prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_63/a_222_392# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_7/a_1178_124#
+ prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_53/X prbs_generator_syn_27/sky130_fd_sc_hs__nand2_2_5/Y
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_61/a_1178_124# prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_1/a_230_79#
+ prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_43/a_230_79# prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_11/a_230_79#
+ prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_41/a_132_392# prbs_generator_syn_27/sky130_fd_sc_hs__nand2_1_13/a_117_74#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_43/a_437_503# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_27/a_544_485#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_63/a_651_503# prbs_generator_syn_27/sky130_fd_sc_hs__nand2_1_7/a_117_74#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_35/a_696_458# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_65/a_544_485#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_51/a_1034_424# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_41/a_735_102#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_32/a_1141_508# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_49/a_1141_508#
+ prbs_generator_syn_27/sky130_fd_sc_hs__nand2_1_55/B prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_53/a_222_392#
+ prbs_generator_syn_27/sky130_fd_sc_hs__sdlclkp_2_1/a_114_112# prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_9/a_293_74#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_43/a_1226_296# prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_29/a_52_123#
+ prbs_generator_syn_27/sky130_fd_sc_hs__nand2_1_37/B prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_1/a_651_503#
+ prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_27/a_376_368# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_4/a_544_485#
+ prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_67/a_376_368# prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_27/X
+ prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_1/X prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_59/a_138_385#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_29/a_1178_124# prbs_generator_syn_27/m3_13600_2871#
+ prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_5/a_230_79# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_23/a_206_368#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_61/a_206_368# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_17/a_544_485#
+ prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_15/a_230_79# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_25/a_696_458#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_55/a_544_485# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_32/a_735_102#
+ prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_29/a_293_74# prbs_generator_syn_27/sky130_fd_sc_hs__nand2_1_17/a_117_74#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_69/a_1034_424# prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_29/a_112_119#
+ prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_37/X prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_31/B
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_19/a_1034_424# prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_33/A
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_9/a_206_368# prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_57/a_376_368#
+ prbs_generator_syn_27/sky130_fd_sc_hs__sdlclkp_2_1/a_706_317# prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_11/B
+ prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_1/a_52_123# prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_39/B
+ prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_21/a_132_392# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_13/a_206_368#
+ prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_43/a_52_123# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_51/a_206_368#
+ prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_47/X prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_23/a_437_503#
+ prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_11/a_52_123# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_61/a_437_503#
+ prbs_generator_syn_27/sky130_fd_sc_hs__nor2b_1_7/Y prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_51/A
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_15/a_696_458# prbs_generator_syn_27/sky130_fd_sc_hs__nor2b_1_5/Y
+ prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_9/a_230_79# prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_25/X
+ prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_19/a_112_119# prbs_generator_syn_27/sky130_fd_sc_hs__nand2_1_45/B
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_5/a_1178_124# prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_19/a_230_79#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_41/a_1226_296# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_59/a_1226_296#
+ prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_63/a_230_79# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_51/Q
+ prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_7/a_132_392# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_9/a_437_503#
+ prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_46/a_376_368# prbs_generator_syn_27/sky130_fd_sc_hs__nand2_1_33/a_117_74#
+ prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_11/a_293_74# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_27/a_1178_124#
+ prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_11/a_132_392# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_13/a_437_503#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_51/a_437_503# prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_5/a_52_123#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_35/a_544_485# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_73/a_651_503#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_45/a_696_458# prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_15/a_52_123#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_47/a_1141_508# prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_47/a_112_119#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_4/a_1178_124# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_17/a_1034_424#
+ prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_23/B prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_37/a_376_368#
+ prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_15/B prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_7/Y
+ prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_29/a_138_385# prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_33/a_230_79#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_25/a_1178_124# prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_47/a_293_74#
+ prbs_generator_syn_27/sky130_fd_sc_hs__nand2_1_37/a_117_74# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_33/a_206_368#
+ prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_15/a_293_74# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_71/a_206_368#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_25/a_544_485# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_67/a_1034_424#
+ prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_13/a_222_392# prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_9/a_52_123#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_15/a_1034_424# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_57/a_1226_296#
+ prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_19/a_52_123# prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_23/X
+ prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_63/a_52_123# prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_19/a_138_385#
+ prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_9/a_376_368# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_21/a_206_368#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_33/a_437_503# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_71/a_437_503#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_53/a_651_503# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_15/a_544_485#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_63/a_696_458# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_65/a_1034_424#
+ prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_19/a_293_74# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_45/a_1141_508#
+ prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_27/a_112_119# prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_67/a_112_119#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_1/a_1178_124# prbs_generator_syn_27/sky130_fd_sc_hs__conb_1_1/a_21_290#
+ prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_63/a_293_74# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_8/a_206_368#
+ prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_17/a_376_368# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_63/a_27_74#
+ prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_21/A prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_55/a_376_368#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_1/a_696_458# prbs_generator_syn_27/sky130_fd_sc_hs__nor2b_1_1/a_278_368#
+ prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_47/a_138_385# prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_33/a_52_123#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_9/a_1034_424# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_21/a_437_503#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_1/a_27_74# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_43/a_651_503#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_1/Q prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_45/a_544_485#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_69/a_735_102# prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_57/a_112_119#
+ prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_31/a_222_392# prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_13/A
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_55/a_1226_296# prbs_generator_syn_27/sky130_fd_sc_hs__nand2_2_5/a_27_74#
+ prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_53/a_230_79# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_8/a_437_503#
+ prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_67/a_293_74# prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_33/a_293_74#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_7/a_735_102# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_23/a_1178_124#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_41/a_206_368# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_8/a_1034_424#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_63/a_1034_424# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_59/a_735_102#
+ prbs_generator_syn_27/sky130_fd_sc_hs__nand2_1_5/B prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_43/a_1141_508#
+ prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_46/a_112_119# prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_61/a_222_392#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_13/a_1034_424# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_73/a_1178_124#
+ prbs_generator_syn_27/sky130_fd_sc_hs__nand2_1_27/B prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_13/B
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_57/a_27_74# prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_57/a_230_79#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_21/a_1178_124# prbs_generator_syn_27/sky130_fd_sc_hs__nor2b_1_1/a_27_112#
+ prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_27/a_138_385# prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_23/a_230_79#
+ prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_67/a_138_385# prbs_generator_syn_27/sky130_fd_sc_hs__nand2_1_41/B
+ prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_9/a_222_392# prbs_generator_syn_27/sky130_fd_sc_hs__nand2_1_27/a_117_74#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_32/a_206_368# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_23/a_651_503#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_41/a_437_503# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_73/a_27_74#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_61/a_651_503# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_63/a_544_485#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_49/a_735_102# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_73/a_696_458#
+ prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_37/a_112_119# prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_51/a_222_392#
+ prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_43/X prbs_generator_syn_27/sky130_fd_sc_hs__nand2_2_1/B
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_9/a_651_503# prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_53/a_52_123#
+ prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_49/X prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_25/a_376_368#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_1/a_544_485# prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_65/a_376_368#
+ prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_57/a_138_385# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_27/a_27_74#
+ prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_39/a_132_392# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_7/a_1034_424#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_13/a_651_503# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_32/a_437_503#
+ prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_27/a_230_79# prbs_generator_syn_27/m3_13600_12265#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_51/a_651_503# prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_59/B
+ prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_47/A prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_61/a_1034_424#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_41/a_1141_508# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_59/a_1141_508#
+ prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_41/a_222_392# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_53/a_1226_296#
+ prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_3/A prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_71/a_1178_124#
+ prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_9/a_112_119# prbs_generator_syn_27/sky130_fd_sc_hs__nand2_1_3/a_117_74#
+ prbs_generator_syn_27/m3_13600_8483# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_39/a_1178_124#
+ prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_57/a_52_123# prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_46/a_138_385#
+ prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_23/a_52_123# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_67/a_27_74#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_53/a_696_458# prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_17/a_112_119#
+ prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_11/A prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_55/a_112_119#
+ prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_1/A prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_51/a_1226_296#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_29/a_1034_424# prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_59/A
+ prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_23/A prbs_generator_syn_27/sky130_fd_sc_hs__nand2_1_39/B
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_5/a_27_74# prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_57/a_293_74#
+ prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_37/a_138_385# prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_59/a_132_392#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_33/a_651_503# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_71/a_651_503#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_43/a_696_458# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_73/a_544_485#
+ prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_27/a_52_123# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_57/a_1141_508#
+ prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_21/a_222_392# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_35/a_27_74#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_69/a_1226_296# prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_37/B
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_19/a_1226_296# prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_35/a_376_368#
+ prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_47/a_230_79# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_37/a_1178_124#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_5/a_1034_424# prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_49/a_132_392#
+ prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_7/a_222_392# prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_27/a_293_74#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_21/a_651_503# prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_9/a_138_385#
+ prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_11/a_222_392# prbs_generator_syn_27/m3_13600_14095#
+ prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_50/A prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_27/a_1034_424#
+ prbs_generator_syn_27/sky130_fd_sc_hs__nand2_1_13/B prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_8/a_651_503#
+ prbs_generator_syn_27/m3_13600_9703# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_35/a_1178_124#
+ prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_17/a_138_385# prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_55/a_138_385#
+ prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_7/a_230_79# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_4/a_1034_424#
+ prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_7/a_376_368# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_69/a_206_368#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_23/a_696_458# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_53/a_544_485#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_39/a_735_102# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_61/a_696_458#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_55/a_1141_508# prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_25/a_112_119#
+ prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_65/a_112_119# prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_43/a_293_74#
+ prbs_generator_syn_27/sky130_fd_sc_hs__nand2_1_57/B prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_25/a_1034_424#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_7/a_206_368# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_17/a_1226_296#
+ prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_15/a_376_368# prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_53/a_376_368#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_9/a_696_458# prbs_generator_syn_27/m3_13600_431#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_45/a_27_74# prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_47/a_52_123#
+ prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_29/a_132_392# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_59/a_206_368#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_69/a_437_503# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_41/a_651_503#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_43/a_544_485# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_13/a_696_458#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_29/a_735_102# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_51/a_696_458#
+ prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_61/Y prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_67/a_1226_296#
+ prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_5/a_132_392# prbs_generator_syn_27/sky130_fd_sc_hs__and2b_2_1/a_198_48#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_7/a_437_503# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_15/a_1226_296#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_69/a_27_74# prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_46/a_293_74#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_1/a_1034_424# prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_19/a_132_392#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_49/a_206_368# prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_7/a_52_123#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_59/a_437_503# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_32/a_651_503#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_7/a_27_74# prbs_generator_syn_27/sky130_fd_sc_hs__nand2_2_1/a_27_74#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_19/a_735_102# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_57/a_735_102#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_65/a_1226_296# prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_37/A
+ prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_33/a_376_368# prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_37/a_230_79#
+ prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_25/a_138_385# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_39/a_27_74#
+ prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_65/a_138_385# prbs_generator_syn_27/sky130_fd_sc_hs__nor2b_1_9/a_278_368#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_49/a_437_503# prbs_generator_syn_27/sky130_fd_sc_hs__and2b_2_1/a_505_74#
+ prbs_generator_syn_27/sky130_fd_sc_hs__nand2_1_51/a_117_74# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_23/a_544_485#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_33/a_696_458# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_61/a_544_485#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_9/a_1226_296# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_53/a_1141_508#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_71/a_696_458# prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_35/a_112_119#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_23/a_1034_424# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_9/a_544_485#
+ prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_63/a_376_368# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_33/a_1178_124#
+ prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_5/a_376_368# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_13/a_544_485#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_73/a_1034_424# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_21/a_696_458#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_51/a_544_485# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_8/a_1226_296#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_51/a_1141_508# prbs_generator_syn_27/sky130_fd_sc_hs__nand2_1_55/a_117_74#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_21/a_1034_424# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_63/a_1226_296#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_23/a_27_74# prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_7/a_112_119#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_13/a_1226_296# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_8/a_696_458#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_32/a_1178_124# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_49/a_1178_124#
+ prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_37/a_52_123# prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_27/a_132_392#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_71/Q prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_67/a_735_102#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_69/a_1141_508# prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_15/a_112_119#
+ prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_53/a_112_119# prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_39/a_222_392#
+ prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_55/a_230_79# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_19/a_1141_508#
+ prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_37/a_293_74# prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_43/a_376_368#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_5/a_735_102# prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_35/a_138_385#
+ prbs_generator_syn_27/sky130_fd_sc_hs__sdlclkp_2_1/a_114_424# prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_57/a_132_392#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_71/a_1034_424# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_7/a_1226_296#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_33/a_544_485# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_41/a_696_458#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_71/a_544_485# prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_21/B
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_61/a_1226_296# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_39/a_1034_424#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_17/a_27_74# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_9/a_27_74#
+ prbs_generator_syn_27/sky130_fd_sc_hs__nor2b_1_5/a_27_112# prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_47/a_132_392#
+ prbs_generator_syn_27/sky130_fd_sc_hs__nor2b_1_8/a_278_368# prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_9/B
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_39/a_206_368# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_33/a_27_74#
+ prbs_generator_syn_27/sky130_fd_sc_hs__nand2_1_41/a_117_74# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_69/a_651_503#
+ prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_51/a_293_74# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_21/a_544_485#
+ prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_7/a_138_385# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_32/a_696_458#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_47/a_735_102# prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_33/a_112_119#
+ prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_59/a_222_392# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_17/a_1141_508#
+ prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_55/a_52_123# prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_3/a_293_74#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_7/a_651_503# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_29/a_1226_296#
+ prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_23/a_376_368# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_8/a_544_485#
+ prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_47/B prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_47/a_1178_124#
+ prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_15/a_138_385# prbs_generator_syn_27/sky130_fd_sc_hs__sdlclkp_2_1/a_1195_374#
+ prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_53/a_138_385# prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_37/a_132_392#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_29/a_206_368# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_39/a_437_503#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_59/a_651_503# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_37/a_735_102#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_67/a_1141_508# prbs_generator_syn_27/sky130_fd_sc_hs__and2b_2_1/a_27_74#
+ prbs_generator_syn_27/sky130_fd_sc_hs__conb_1_1/a_165_290# prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_55/a_293_74#
+ prbs_generator_syn_27/sky130_fd_sc_hs__nand2_1_45/a_117_74# prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_63/a_112_119#
+ prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_49/a_222_392# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_37/a_1034_424#
+ prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_23/a_293_74# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_15/a_1141_508#
+ prbs_generator_syn_27/sky130_fd_sc_hs__nand2_1_5/a_117_74# prbs_generator_syn_27/m3_13600_13485#
+ prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_5/a_112_119# prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_13/a_376_368#
+ prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_51/a_376_368# prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_7/a_293_74#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_19/a_206_368# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_57/a_206_368#
+ prbs_generator_syn_27/sky130_fd_sc_hs__sdlclkp_2_1/a_318_74# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_29/a_437_503#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_49/a_651_503# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_25/a_27_74#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_5/a_1226_296# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_41/a_544_485#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_27/a_735_102# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_65/a_1141_508#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_65/a_735_102# prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_3/a_230_79#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_35/a_1034_424# prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_13/a_230_79#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_41/a_27_74# prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_3/a_132_392#
+ prbs_generator_syn_27/sky130_fd_sc_hs__nand2_1_49/a_117_74# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_27/a_1226_296#
+ prbs_generator_syn_27/sky130_fd_sc_hs__nand2_1_15/a_117_74# prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_41/a_376_368#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_45/a_1178_124# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_4/a_735_102#
+ prbs_generator_syn_27/sky130_fd_sc_hs__nand2_1_9/a_117_74# prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_33/a_138_385#
+ prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_17/a_132_392# prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_55/a_132_392#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_9/a_1141_508# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_19/a_437_503#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_57/a_437_503# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_4/a_1226_296#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_32/a_544_485# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_17/a_735_102#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_55/a_735_102# prbs_generator_syn_27/m3_13600_2261#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_65/a_27_74# prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_29/a_222_392#
+ prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_43/a_112_119# prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_19/X
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_25/a_1226_296# prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_31/a_376_368#
+ prbs_generator_syn_27/sky130_fd_sc_hs__or2_1_1/a_63_368# prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_17/a_230_79#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_4/a_27_74# prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_61/a_230_79#
+ prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_63/a_138_385# prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_5/a_222_392#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_8/a_1141_508# prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_41/a_293_74#
+ prbs_generator_syn_27/sky130_fd_sc_hs__nand2_1_31/a_117_74# prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_5/a_138_385#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_63/a_1141_508# prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_19/a_222_392#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_13/a_1141_508# prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_3/a_52_123#
+ prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_13/a_52_123# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_43/a_1178_124#
+ prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_61/a_376_368# prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_35/a_132_392#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_67/a_206_368# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_1/a_1226_296#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_69/a_696_458# prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_31/a_230_79#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_35/a_735_102# prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_23/a_112_119#
+ prbs_generator_syn_27/sky130_fd_sc_hs__nand2_1_35/a_117_74# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_59/a_27_74#
+ prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_13/a_293_74# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_5/a_206_368#
+ prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_50/a_376_368# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_7/a_696_458#
+ prbs_generator_syn_27/sky130_fd_sc_hs__nor2b_1_7/a_278_368# prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_17/a_52_123#
+ prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_43/a_138_385# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_7/a_1141_508#
+ prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_61/a_52_123# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_67/a_437_503#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_61/a_1141_508# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_25/a_735_102#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_59/a_696_458# prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_13/a_112_119#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_33/a_1034_424# prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_51/a_112_119#
+ prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_35/a_230_79# prbs_generator_syn_27/m3_13600_4091#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_23/a_1226_296# prbs_generator_syn_27/sky130_fd_sc_hs__nand2_1_39/a_117_74#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_29/a_27_74# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_5/a_437_503#
+ prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_17/a_293_74# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_41/a_1178_124#
+ prbs_generator_syn_27/sky130_fd_sc_hs__or2_1_1/a_152_368# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_59/a_1178_124#
+ prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_61/a_293_74# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_47/a_206_368#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_39/a_651_503# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_49/a_696_458#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_15/a_735_102# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_32/a_1034_424#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_73/a_1226_296# prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_27/a_222_392#
+ prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_41/a_112_119# prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_31/a_52_123#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_49/a_1034_424# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_29/a_1141_508#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_21/a_1226_296# prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_39/a_230_79#
+ prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_23/a_138_385# prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_51/a_230_79#
+ prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_45/a_132_392# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_37/a_206_368#
+ prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_65/a_293_74# prbs_generator_syn_27/sky130_fd_sc_hs__nand2_1_53/a_117_74#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_47/a_437_503# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_29/a_651_503#
+ prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_31/a_293_74# prbs_generator_syn_27/sky130_fd_sc_hs__nand2_1_21/a_117_74#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_69/a_544_485# prbs_generator_syn_27/sky130_fd_sc_hs__clkbuf_16_1/a_114_74#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_45/a_735_102# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_13/a_27_74#
+ prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_31/a_112_119# prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_57/a_222_392#
+ prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_35/a_52_123# prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_21/a_376_368#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_7/a_544_485# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_57/a_1178_124#
+ prbs_generator_syn_27/m3_13600_6043# prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_13/a_138_385#
+ prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_51/a_138_385# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_5/a_1141_508#
+ prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_3/a_376_368# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_27/a_206_368#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_65/a_206_368# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_37/a_437_503#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_19/a_651_503# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_57/a_651_503#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_59/a_544_485# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_71/a_1226_296#
+ prbs_generator_syn_27/sky130_fd_sc_hs__nand2_1_25/a_117_74# prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_61/a_112_119#
+ prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_47/a_222_392# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_27/a_1141_508#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_53/a_27_74# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_4/a_206_368#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_39/a_1226_296# prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_11/a_376_368#
+ prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_39/a_52_123# prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_41/a_138_385#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_4/a_1141_508# prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_25/a_132_392#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_17/a_206_368# prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_41/A
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_55/a_206_368# prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_51/a_52_123#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_27/a_437_503# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_65/a_437_503#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_49/a_544_485# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_63/a_735_102#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_47/a_1034_424# prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_50/a_112_119#
+ prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_37/a_222_392# prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_59/a_230_79#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_25/a_1141_508# prbs_generator_syn_27/sky130_fd_sc_hs__nor2b_1_4/a_27_112#
+ prbs_generator_syn_27/sky130_fd_sc_hs__sdlclkp_2_1/a_685_81# prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_1/a_132_392#
+ prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_39/a_293_74# prbs_generator_syn_27/sky130_fd_sc_hs__nand2_1_29/a_117_74#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_4/a_437_503# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_55/a_1178_124#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_21/a_27_74# prbs_generator_syn_27/m3_13600_12875#
+ prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_50/a_293_74# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_1/a_735_102#
+ prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_31/a_138_385# prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_15/a_132_392#
+ prbs_generator_syn_27/sky130_fd_sc_hs__nand2_1_1/a_117_74# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_17/a_437_503#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_55/a_437_503# prbs_generator_syn
Xsky130_fd_sc_hs__conb_1_6 DVSS: DVDD: DVDD: DVSS: prbs_generator_syn_3/eqn[9] sky130_fd_sc_hs__conb_1_7/HI
+ sky130_fd_sc_hs__conb_1_7/a_165_290# sky130_fd_sc_hs__conb_1_7/a_21_290# sky130_fd_sc_hs__conb_1
Xsky130_fd_sc_hs__buf_2_102 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__buf_2_103/A sky130_fd_sc_hs__buf_2_103/X
+ sky130_fd_sc_hs__buf_2_103/a_21_260# sky130_fd_sc_hs__buf_2
Xsky130_fd_sc_hs__buf_2_113 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__buf_2_113/A sky130_fd_sc_hs__buf_2_113/X
+ sky130_fd_sc_hs__buf_2_113/a_21_260# sky130_fd_sc_hs__buf_2
Xsky130_fd_sc_hs__buf_2_124 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__buf_2_125/A sky130_fd_sc_hs__buf_2_125/X
+ sky130_fd_sc_hs__buf_2_125/a_21_260# sky130_fd_sc_hs__buf_2
Xsky130_fd_sc_hs__buf_2_135 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__buf_2_135/A sky130_fd_sc_hs__buf_2_135/X
+ sky130_fd_sc_hs__buf_2_135/a_21_260# sky130_fd_sc_hs__buf_2
Xsky130_fd_sc_hs__buf_2_146 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__buf_2_147/A sky130_fd_sc_hs__buf_2_147/X
+ sky130_fd_sc_hs__buf_2_147/a_21_260# sky130_fd_sc_hs__buf_2
Xsky130_fd_sc_hs__buf_2_157 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__buf_2_157/A sky130_fd_sc_hs__buf_2_157/X
+ sky130_fd_sc_hs__buf_2_157/a_21_260# sky130_fd_sc_hs__buf_2
Xsky130_fd_sc_hs__einvp_2_14 DVSS: DVDD: DVDD: DVSS: dout_n sky130_fd_sc_hs__buf_8_1/A
+ sky130_fd_sc_hs__dlrtp_1_13/Q sky130_fd_sc_hs__einvp_2_15/a_263_323# sky130_fd_sc_hs__einvp_2_15/a_36_74#
+ sky130_fd_sc_hs__einvp_2_15/a_27_368# sky130_fd_sc_hs__einvp_2
Xsky130_fd_sc_hs__einvp_2_25 DVSS: DVDD: DVDD: DVSS: dout_n sky130_fd_sc_hs__einvp_2_9/A
+ sky130_fd_sc_hs__dlrtp_1_19/Q sky130_fd_sc_hs__einvp_2_25/a_263_323# sky130_fd_sc_hs__einvp_2_25/a_36_74#
+ sky130_fd_sc_hs__einvp_2_25/a_27_368# sky130_fd_sc_hs__einvp_2
Xsky130_fd_sc_hs__einvp_2_36 DVSS: DVDD: DVDD: DVSS: dout_n sky130_fd_sc_hs__buf_8_1/A
+ sky130_fd_sc_hs__dlrtp_1_24/Q sky130_fd_sc_hs__einvp_2_37/a_263_323# sky130_fd_sc_hs__einvp_2_37/a_36_74#
+ sky130_fd_sc_hs__einvp_2_37/a_27_368# sky130_fd_sc_hs__einvp_2
Xsky130_fd_sc_hs__einvp_2_47 DVSS: DVDD: DVDD: DVSS: dout_n sky130_fd_sc_hs__buf_8_1/A
+ sky130_fd_sc_hs__dlrtp_1_33/Q sky130_fd_sc_hs__einvp_2_47/a_263_323# sky130_fd_sc_hs__einvp_2_47/a_36_74#
+ sky130_fd_sc_hs__einvp_2_47/a_27_368# sky130_fd_sc_hs__einvp_2
Xsky130_fd_sc_hs__einvp_2_58 DVSS: DVDD: DVDD: DVSS: dout_p sky130_fd_sc_hs__einvp_2_99/A
+ sky130_fd_sc_hs__dlrtp_1_43/Q sky130_fd_sc_hs__einvp_2_59/a_263_323# sky130_fd_sc_hs__einvp_2_59/a_36_74#
+ sky130_fd_sc_hs__einvp_2_59/a_27_368# sky130_fd_sc_hs__einvp_2
Xsky130_fd_sc_hs__einvp_2_69 DVSS: DVDD: DVDD: DVSS: dout_p sky130_fd_sc_hs__einvp_2_97/A
+ sky130_fd_sc_hs__dlrtp_1_59/Q sky130_fd_sc_hs__einvp_2_69/a_263_323# sky130_fd_sc_hs__einvp_2_69/a_36_74#
+ sky130_fd_sc_hs__einvp_2_69/a_27_368# sky130_fd_sc_hs__einvp_2
Xsky130_fd_sc_hs__conb_1_13 DVSS: DVDD: DVDD: DVSS: prbs_generator_syn_9/eqn[9] sky130_fd_sc_hs__conb_1_13/HI
+ sky130_fd_sc_hs__conb_1_13/a_165_290# sky130_fd_sc_hs__conb_1_13/a_21_290# sky130_fd_sc_hs__conb_1
Xsky130_fd_sc_hs__conb_1_24 DVSS: DVDD: DVDD: DVSS: prbs_generator_syn_1/eqn[31] prbs_generator_syn_1/cke
+ sky130_fd_sc_hs__conb_1_25/a_165_290# sky130_fd_sc_hs__conb_1_25/a_21_290# sky130_fd_sc_hs__conb_1
Xsky130_fd_sc_hs__conb_1_35 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__conb_1_35/LO
+ sky130_fd_sc_hs__conb_1_35/HI sky130_fd_sc_hs__conb_1_35/a_165_290# sky130_fd_sc_hs__conb_1_35/a_21_290#
+ sky130_fd_sc_hs__conb_1
Xsky130_fd_sc_hs__conb_1_46 DVSS: DVDD: DVDD: DVSS: prbs_generator_syn_3/eqn[31] prbs_generator_syn_3/cke
+ sky130_fd_sc_hs__conb_1_47/a_165_290# sky130_fd_sc_hs__conb_1_47/a_21_290# sky130_fd_sc_hs__conb_1
Xsky130_fd_sc_hs__conb_1_57 DVSS: DVDD: DVDD: DVSS: prbs_generator_syn_9/eqn[31] prbs_generator_syn_9/cke
+ sky130_fd_sc_hs__conb_1_57/a_165_290# sky130_fd_sc_hs__conb_1_57/a_21_290# sky130_fd_sc_hs__conb_1
Xsky130_fd_sc_hs__conb_1_68 DVSS: DVDD: DVDD: DVSS: prbs_generator_syn_7/eqn[28] sky130_fd_sc_hs__conb_1_69/HI
+ sky130_fd_sc_hs__conb_1_69/a_165_290# sky130_fd_sc_hs__conb_1_69/a_21_290# sky130_fd_sc_hs__conb_1
Xsky130_fd_sc_hs__inv_4_20 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__inv_4_21/Y sky130_fd_sc_hs__inv_4_21/A
+ sky130_fd_sc_hs__inv_4
Xsky130_fd_sc_hs__inv_4_31 DVSS: DVDD: DVDD: DVSS: osc_core_1/pi1_r[3] osc_core_1/pi1_l[3]
+ sky130_fd_sc_hs__inv_4
Xsky130_fd_sc_hs__conb_1_79 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__conb_1_79/LO
+ sky130_fd_sc_hs__conb_1_79/HI sky130_fd_sc_hs__conb_1_79/a_165_290# sky130_fd_sc_hs__conb_1_79/a_21_290#
+ sky130_fd_sc_hs__conb_1
Xsky130_fd_sc_hs__inv_4_42 DVSS: DVDD: DVDD: DVSS: osc_core_1/pi2_r[1] osc_core_1/pi2_l[1]
+ sky130_fd_sc_hs__inv_4
Xsky130_fd_sc_hs__inv_4_53 DVSS: DVDD: DVDD: DVSS: osc_core_1/pi4_r[3] osc_core_1/pi4_l[3]
+ sky130_fd_sc_hs__inv_4
Xsky130_fd_sc_hs__inv_4_64 DVSS: DVDD: DVDD: DVSS: osc_core_1/pi3_r[1] osc_core_1/pi3_l[1]
+ sky130_fd_sc_hs__inv_4
Xsky130_fd_sc_hs__inv_4_75 DVSS: DVDD: DVDD: DVSS: osc_core_1/pi5_r[1] osc_core_1/pi5_l[1]
+ sky130_fd_sc_hs__inv_4
Xsky130_fd_sc_hs__inv_4_86 DVSS: DVDD: DVDD: DVSS: hr_16t4_mux_top_3/din[2] hr_16t4_mux_top_1/din[2]
+ sky130_fd_sc_hs__inv_4
Xsky130_fd_sc_hs__dlrtp_1_15 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__dlrtp_1_15/Q
+ sky130_fd_sc_hs__clkbuf_2_3/X sky130_fd_sc_hs__conb_1_119/HI sky130_fd_sc_hs__buf_2_103/X
+ sky130_fd_sc_hs__dlrtp_1_15/a_216_424# sky130_fd_sc_hs__dlrtp_1_15/a_759_508# sky130_fd_sc_hs__dlrtp_1_15/a_565_74#
+ sky130_fd_sc_hs__dlrtp_1_15/a_27_424# sky130_fd_sc_hs__dlrtp_1_15/a_1045_74# sky130_fd_sc_hs__dlrtp_1_15/a_643_74#
+ sky130_fd_sc_hs__dlrtp_1_15/a_817_48# sky130_fd_sc_hs__dlrtp_1_15/a_568_392# sky130_fd_sc_hs__dlrtp_1_15/a_363_74#
+ sky130_fd_sc_hs__dlrtp_1_15/a_769_74# sky130_fd_sc_hs__dlrtp_1
Xsky130_fd_sc_hs__dlrtp_1_26 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__dlrtp_1_27/Q
+ sky130_fd_sc_hs__clkbuf_2_3/A sky130_fd_sc_hs__conb_1_119/HI sky130_fd_sc_hs__dlrtp_1_27/D
+ sky130_fd_sc_hs__dlrtp_1_27/a_216_424# sky130_fd_sc_hs__dlrtp_1_27/a_759_508# sky130_fd_sc_hs__dlrtp_1_27/a_565_74#
+ sky130_fd_sc_hs__dlrtp_1_27/a_27_424# sky130_fd_sc_hs__dlrtp_1_27/a_1045_74# sky130_fd_sc_hs__dlrtp_1_27/a_643_74#
+ sky130_fd_sc_hs__dlrtp_1_27/a_817_48# sky130_fd_sc_hs__dlrtp_1_27/a_568_392# sky130_fd_sc_hs__dlrtp_1_27/a_363_74#
+ sky130_fd_sc_hs__dlrtp_1_27/a_769_74# sky130_fd_sc_hs__dlrtp_1
Xsky130_fd_sc_hs__dlrtp_1_37 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__dlrtp_1_37/Q
+ sky130_fd_sc_hs__clkbuf_2_3/A sky130_fd_sc_hs__conb_1_121/HI sky130_fd_sc_hs__buf_2_135/X
+ sky130_fd_sc_hs__dlrtp_1_37/a_216_424# sky130_fd_sc_hs__dlrtp_1_37/a_759_508# sky130_fd_sc_hs__dlrtp_1_37/a_565_74#
+ sky130_fd_sc_hs__dlrtp_1_37/a_27_424# sky130_fd_sc_hs__dlrtp_1_37/a_1045_74# sky130_fd_sc_hs__dlrtp_1_37/a_643_74#
+ sky130_fd_sc_hs__dlrtp_1_37/a_817_48# sky130_fd_sc_hs__dlrtp_1_37/a_568_392# sky130_fd_sc_hs__dlrtp_1_37/a_363_74#
+ sky130_fd_sc_hs__dlrtp_1_37/a_769_74# sky130_fd_sc_hs__dlrtp_1
Xsky130_fd_sc_hs__dlrtp_1_48 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__dlrtp_1_49/Q
+ sky130_fd_sc_hs__clkbuf_16_53/A sky130_fd_sc_hs__conb_1_123/HI sky130_fd_sc_hs__buf_2_29/X
+ sky130_fd_sc_hs__dlrtp_1_49/a_216_424# sky130_fd_sc_hs__dlrtp_1_49/a_759_508# sky130_fd_sc_hs__dlrtp_1_49/a_565_74#
+ sky130_fd_sc_hs__dlrtp_1_49/a_27_424# sky130_fd_sc_hs__dlrtp_1_49/a_1045_74# sky130_fd_sc_hs__dlrtp_1_49/a_643_74#
+ sky130_fd_sc_hs__dlrtp_1_49/a_817_48# sky130_fd_sc_hs__dlrtp_1_49/a_568_392# sky130_fd_sc_hs__dlrtp_1_49/a_363_74#
+ sky130_fd_sc_hs__dlrtp_1_49/a_769_74# sky130_fd_sc_hs__dlrtp_1
Xsky130_fd_sc_hs__dlrtp_1_59 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__dlrtp_1_59/Q
+ sky130_fd_sc_hs__clkbuf_16_53/A sky130_fd_sc_hs__conb_1_125/HI sky130_fd_sc_hs__buf_2_55/X
+ sky130_fd_sc_hs__dlrtp_1_59/a_216_424# sky130_fd_sc_hs__dlrtp_1_59/a_759_508# sky130_fd_sc_hs__dlrtp_1_59/a_565_74#
+ sky130_fd_sc_hs__dlrtp_1_59/a_27_424# sky130_fd_sc_hs__dlrtp_1_59/a_1045_74# sky130_fd_sc_hs__dlrtp_1_59/a_643_74#
+ sky130_fd_sc_hs__dlrtp_1_59/a_817_48# sky130_fd_sc_hs__dlrtp_1_59/a_568_392# sky130_fd_sc_hs__dlrtp_1_59/a_363_74#
+ sky130_fd_sc_hs__dlrtp_1_59/a_769_74# sky130_fd_sc_hs__dlrtp_1
Xsky130_fd_sc_hs__einvp_2_8 DVSS: DVDD: DVDD: DVSS: dout_n sky130_fd_sc_hs__einvp_2_9/A
+ sky130_fd_sc_hs__dlrtp_1_9/Q sky130_fd_sc_hs__einvp_2_9/a_263_323# sky130_fd_sc_hs__einvp_2_9/a_36_74#
+ sky130_fd_sc_hs__einvp_2_9/a_27_368# sky130_fd_sc_hs__einvp_2
Xsky130_fd_sc_hs__clkbuf_16_80 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__or2b_2_1/A
+ sky130_fd_sc_hs__clkbuf_8_75/X sky130_fd_sc_hs__clkbuf_16_81/a_114_74# sky130_fd_sc_hs__clkbuf_16
Xsky130_fd_sc_hs__clkbuf_16_91 DVSS: DVDD: DVDD: DVSS: prbs_generator_syn_19/inj_err
+ prbs_generator_syn_31/inj_err sky130_fd_sc_hs__clkbuf_16_91/a_114_74# sky130_fd_sc_hs__clkbuf_16
Xsky130_fd_sc_hs__buf_2_18 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__buf_2_33/A sky130_fd_sc_hs__buf_2_19/X
+ sky130_fd_sc_hs__buf_2_19/a_21_260# sky130_fd_sc_hs__buf_2
Xsky130_fd_sc_hs__buf_2_29 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__buf_2_39/X sky130_fd_sc_hs__buf_2_29/X
+ sky130_fd_sc_hs__buf_2_29/a_21_260# sky130_fd_sc_hs__buf_2
Xsky130_fd_sc_hs__nand2_2_10 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__inv_4_17/A sky130_fd_sc_hs__nand2_2_11/B
+ sky130_fd_sc_hs__inv_4_15/Y sky130_fd_sc_hs__nand2_2_11/a_27_74# sky130_fd_sc_hs__nand2_2
Xsky130_fd_sc_hs__nand2_2_21 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__inv_4_25/A sky130_fd_sc_hs__nand2_2_21/B
+ sky130_fd_sc_hs__nand2_2_27/B sky130_fd_sc_hs__nand2_2_21/a_27_74# sky130_fd_sc_hs__nand2_2
Xsky130_fd_sc_hs__nand2_2_32 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__nand2_2_33/Y
+ sky130_fd_sc_hs__or4_2_1/B sky130_fd_sc_hs__or4_2_1/A sky130_fd_sc_hs__nand2_2_33/a_27_74#
+ sky130_fd_sc_hs__nand2_2
Xsky130_fd_sc_hs__conb_1_207 DVSS: DVDD: DVDD: DVSS: prbs_generator_syn_19/eqn[31]
+ prbs_generator_syn_19/cke sky130_fd_sc_hs__conb_1_207/a_165_290# sky130_fd_sc_hs__conb_1_207/a_21_290#
+ sky130_fd_sc_hs__conb_1
Xsky130_fd_sc_hs__conb_1_218 DVSS: DVDD: DVDD: DVSS: prbs_generator_syn_25/eqn[30]
+ sky130_fd_sc_hs__conb_1_219/HI sky130_fd_sc_hs__conb_1_219/a_165_290# sky130_fd_sc_hs__conb_1_219/a_21_290#
+ sky130_fd_sc_hs__conb_1
Xsky130_fd_sc_hs__conb_1_229 DVSS: DVDD: DVDD: DVSS: prbs_generator_syn_23/eqn[31]
+ prbs_generator_syn_23/cke sky130_fd_sc_hs__conb_1_229/a_165_290# sky130_fd_sc_hs__conb_1_229/a_21_290#
+ sky130_fd_sc_hs__conb_1
Xsky130_fd_sc_hs__o21bai_2_6 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__nand2_2_7/A
+ sky130_fd_sc_hs__inv_8_1/Y sky130_fd_sc_hs__dlrtp_1_71/D sky130_fd_sc_hs__buf_2_59/A
+ sky130_fd_sc_hs__o21bai_2_7/a_27_74# sky130_fd_sc_hs__o21bai_2_7/a_225_74# sky130_fd_sc_hs__o21bai_2_7/a_507_368#
+ sky130_fd_sc_hs__o21bai_2
Xsky130_fd_sc_hs__o21ai_2_11 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__inv_4_11/Y sky130_fd_sc_hs__nand2_2_3/B
+ sky130_fd_sc_hs__o21ai_2_55/A1 sky130_fd_sc_hs__o21ai_2_11/Y sky130_fd_sc_hs__o21ai_2_11/a_116_368#
+ sky130_fd_sc_hs__o21ai_2_11/a_27_74# sky130_fd_sc_hs__o21ai_2
Xsky130_fd_sc_hs__o21ai_2_22 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__inv_4_15/Y sky130_fd_sc_hs__o21ai_2_23/A2
+ sky130_fd_sc_hs__buf_2_77/X sky130_fd_sc_hs__o21ai_2_23/Y sky130_fd_sc_hs__o21ai_2_23/a_116_368#
+ sky130_fd_sc_hs__o21ai_2_23/a_27_74# sky130_fd_sc_hs__o21ai_2
Xsky130_fd_sc_hs__o21ai_2_33 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__inv_4_19/Y sky130_fd_sc_hs__clkinv_4_7/Y
+ sky130_fd_sc_hs__o21ai_4_1/A1 sky130_fd_sc_hs__buf_2_89/A sky130_fd_sc_hs__o21ai_2_33/a_116_368#
+ sky130_fd_sc_hs__o21ai_2_33/a_27_74# sky130_fd_sc_hs__o21ai_2
Xsky130_fd_sc_hs__o21ai_2_44 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__nand2_2_27/B
+ sky130_fd_sc_hs__nand2_2_21/B sky130_fd_sc_hs__or2b_4_1/A sky130_fd_sc_hs__o21ai_2_45/Y
+ sky130_fd_sc_hs__o21ai_2_45/a_116_368# sky130_fd_sc_hs__o21ai_2_45/a_27_74# sky130_fd_sc_hs__o21ai_2
Xsky130_fd_sc_hs__o21ai_2_55 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__inv_4_29/A sky130_fd_sc_hs__nand2_2_5/B
+ sky130_fd_sc_hs__o21ai_2_55/A1 sky130_fd_sc_hs__buf_2_149/A sky130_fd_sc_hs__o21ai_2_55/a_116_368#
+ sky130_fd_sc_hs__o21ai_2_55/a_27_74# sky130_fd_sc_hs__o21ai_2
Xsky130_fd_sc_hs__clkinv_4_14 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__o21ai_2_55/A1
+ sky130_fd_sc_hs__or4_2_1/B sky130_fd_sc_hs__clkinv_4
Xprbs_generator_syn_16 prbs_generator_syn_19/clk prbs_generator_syn_19/rst prbs_generator_syn_17/cke
+ sky130_fd_sc_hs__conb_1_161/LO sky130_fd_sc_hs__conb_1_161/LO sky130_fd_sc_hs__conb_1_161/LO
+ sky130_fd_sc_hs__conb_1_161/HI sky130_fd_sc_hs__conb_1_161/HI sky130_fd_sc_hs__conb_1_161/HI
+ sky130_fd_sc_hs__conb_1_161/HI sky130_fd_sc_hs__conb_1_161/HI sky130_fd_sc_hs__conb_1_161/LO
+ sky130_fd_sc_hs__conb_1_161/LO sky130_fd_sc_hs__conb_1_161/LO prbs_generator_syn_17/eqn[31]
+ prbs_generator_syn_19/eqn[13] prbs_generator_syn_19/eqn[13] sky130_fd_sc_hs__conb_1_193/HI
+ prbs_generator_syn_19/eqn[13] sky130_fd_sc_hs__conb_1_193/HI prbs_generator_syn_19/eqn[13]
+ prbs_generator_syn_17/eqn[1] prbs_generator_syn_17/eqn[2] prbs_generator_syn_17/eqn[1]
+ prbs_generator_syn_17/eqn[2] prbs_generator_syn_17/eqn[1] prbs_generator_syn_17/eqn[2]
+ sky130_fd_sc_hs__conb_1_165/LO sky130_fd_sc_hs__conb_1_165/HI sky130_fd_sc_hs__conb_1_165/HI
+ sky130_fd_sc_hs__conb_1_165/LO sky130_fd_sc_hs__conb_1_165/LO sky130_fd_sc_hs__conb_1_165/LO
+ sky130_fd_sc_hs__conb_1_165/LO sky130_fd_sc_hs__conb_1_165/LO prbs_generator_syn_17/eqn[31]
+ prbs_generator_syn_17/eqn[30] prbs_generator_syn_17/eqn[30] prbs_generator_syn_17/eqn[30]
+ prbs_generator_syn_17/eqn[30] prbs_generator_syn_17/eqn[30] prbs_generator_syn_17/eqn[30]
+ prbs_generator_syn_17/eqn[30] prbs_generator_syn_17/eqn[30] prbs_generator_syn_17/eqn[22]
+ prbs_generator_syn_17/eqn[22] prbs_generator_syn_17/eqn[20] prbs_generator_syn_17/eqn[22]
+ prbs_generator_syn_17/eqn[22] prbs_generator_syn_17/eqn[22] prbs_generator_syn_17/eqn[22]
+ prbs_generator_syn_17/eqn[22] prbs_generator_syn_17/eqn[22] prbs_generator_syn_17/eqn[13]
+ prbs_generator_syn_17/eqn[13] prbs_generator_syn_17/eqn[13] prbs_generator_syn_17/eqn[9]
+ prbs_generator_syn_17/eqn[9] prbs_generator_syn_17/eqn[9] prbs_generator_syn_17/eqn[9]
+ prbs_generator_syn_17/eqn[9] prbs_generator_syn_17/eqn[9] prbs_generator_syn_17/eqn[9]
+ prbs_generator_syn_17/eqn[9] prbs_generator_syn_17/eqn[2] prbs_generator_syn_17/eqn[1]
+ prbs_generator_syn_17/eqn[2] prbs_generator_syn_19/inj_err prbs_generator_syn_17/eqn[31]
+ prbs_generator_syn_17/eqn[31] prbs_generator_syn_17/out DVSS: DVDD: prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_1/a_293_74#
+ prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_15/X prbs_generator_syn_17/sky130_fd_sc_hs__nand2_1_35/B
+ prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_51/Y prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_9/A
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_9/CLK prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_47/a_27_74#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_37/a_1226_296# prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_3/B
+ prbs_generator_syn_17/sky130_fd_sc_hs__nor2b_1_7/a_27_112# prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_29/B
+ prbs_generator_syn_17/sky130_fd_sc_hs__sdlclkp_2_1/a_580_74# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_1/a_1141_508#
+ prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_5/Y prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_41/a_230_79#
+ prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_61/a_138_385# prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_43/a_132_392#
+ prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_3/a_222_392# prbs_generator_syn_17/sky130_fd_sc_hs__nor2b_1_9/a_27_112#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_61/a_27_74# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_35/a_206_368#
+ prbs_generator_syn_17/sky130_fd_sc_hs__nand2_2_3/Y prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_25/B
+ prbs_generator_syn_17/sky130_fd_sc_hs__nand2_1_11/a_117_74# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_67/a_651_503#
+ prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_45/X prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_39/a_696_458#
+ prbs_generator_syn_17/sky130_fd_sc_hs__sdlclkp_2_1/a_1198_74# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_45/a_1034_424#
+ prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_17/a_222_392# prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_55/a_222_392#
+ prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_53/Y prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_35/A
+ prbs_generator_syn_17/m3_13600_1651# prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_59/a_52_123#
+ prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_5/a_293_74# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_35/a_1226_296#
+ prbs_generator_syn_17/sky130_fd_sc_hs__nand2_1_51/B prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_5/a_651_503#
+ prbs_generator_syn_17/sky130_fd_sc_hs__nand2_1_21/B prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_8/a_27_74#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_15/a_27_74# prbs_generator_syn_17/sky130_fd_sc_hs__and2b_2_1/X
+ prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_13/X prbs_generator_syn_17/sky130_fd_sc_hs__nand2_2_3/a_27_74#
+ prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_50/a_138_385# prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_33/a_132_392#
+ prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_1/a_376_368# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_25/a_206_368#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_35/a_437_503# prbs_generator_syn_17/sky130_fd_sc_hs__sdlclkp_2_1/a_708_451#
+ prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_45/a_230_79# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_29/a_696_458#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_32/a_27_74# prbs_generator_syn_17/sky130_fd_sc_hs__nor2b_1_4/Y
+ prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_59/a_293_74# prbs_generator_syn_17/sky130_fd_sc_hs__nand2_1_47/a_117_74#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_73/a_735_102# prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_21/a_112_119#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_23/a_1141_508# prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_25/a_293_74#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_7/Q prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_3/a_112_119#
+ prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_35/B prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_51/X
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_53/a_1178_124# prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_23/a_132_392#
+ prbs_generator_syn_17/sky130_fd_sc_hs__nand2_1_3/B prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_15/a_206_368#
+ prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_63/a_132_392# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_55/a_27_74#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_25/a_437_503# prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_41/a_52_123#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_47/a_651_503# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_73/a_1141_508#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_19/a_696_458# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_57/a_696_458#
+ prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_7/X prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_43/a_1034_424#
+ prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_55/A prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_11/a_112_119#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_21/a_1141_508# prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_35/a_222_392#
+ prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_49/a_230_79# prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_67/Y
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_71/a_27_74# prbs_generator_syn_17/sky130_fd_sc_hs__nand2_1_33/B
+ prbs_generator_syn_17/sky130_fd_sc_hs__conb_1_1/LO prbs_generator_syn_17/sky130_fd_sc_hs__nand2_1_19/a_117_74#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_51/a_1178_124# prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_33/X
+ prbs_generator_syn_17/sky130_fd_sc_hs__nand2_1_29/B prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_41/Y
+ prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_53/a_132_392# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_45/a_206_368#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_15/a_437_503# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_37/a_651_503#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_39/a_544_485# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_53/a_735_102#
+ prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_45/a_52_123# prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_1/B
+ prbs_generator_syn_17/sky130_fd_sc_hs__nand2_2_3/B prbs_generator_syn_17/sky130_fd_sc_hs__clkbuf_16_1/A
+ prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_21/X prbs_generator_syn_17/sky130_fd_sc_hs__nand2_1_25/B
+ prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_39/a_376_368# prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_63/X
+ prbs_generator_syn_17/m3_13600_3481# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_69/a_1178_124#
+ prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_21/a_138_385# prbs_generator_syn_17/sky130_fd_sc_hs__nor2b_1_8/Y
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_19/a_1178_124# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_49/a_27_74#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_45/a_437_503# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_27/a_651_503#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_71/a_1141_508# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_65/a_651_503#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_29/a_544_485# prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_3/a_138_385#
+ prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_55/X prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_43/a_735_102#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_41/a_1034_424# prbs_generator_syn_17/sky130_fd_sc_hs__nand2_1_9/B
+ prbs_generator_syn_17/sky130_fd_sc_hs__nor2b_1_9/Y prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_59/a_1034_424#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_39/a_1141_508# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_33/a_1226_296#
+ prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_49/a_52_123# prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_47/Y
+ prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_43/Y prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_4/a_651_503#
+ prbs_generator_syn_17/sky130_fd_sc_hs__nand2_1_49/B prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_19/A
+ prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_11/a_138_385# prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_5/X
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_63/a_206_368# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_17/a_651_503#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_19/a_544_485# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_55/a_651_503#
+ prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_9/Y prbs_generator_syn_17/sky130_fd_sc_hs__nand2_1_17/B
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_57/a_544_485# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_67/a_696_458#
+ prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_35/X prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_19/a_27_74#
+ prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_45/a_222_392# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_32/a_1226_296#
+ prbs_generator_syn_17/sky130_fd_sc_hs__nand2_1_43/B prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_25/A
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_1/a_206_368# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_49/a_1226_296#
+ prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_1/a_112_119# prbs_generator_syn_17/sky130_fd_sc_hs__or2_1_1/X
+ prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_59/a_376_368# prbs_generator_syn_17/sky130_fd_sc_hs__nand2_1_19/B
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_5/a_696_458# prbs_generator_syn_17/sky130_fd_sc_hs__nor2b_1_1/Y
+ prbs_generator_syn_17/sky130_fd_sc_hs__nor2b_1_5/a_278_368# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_17/a_1178_124#
+ prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_39/X prbs_generator_syn_17/m3_13600_5433#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_63/a_437_503# prbs_generator_syn_17/sky130_fd_sc_hs__nand2_2_5/B
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_23/a_735_102# prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_53/A
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_61/a_735_102# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_57/a_1034_424#
+ prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_63/B prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_37/a_1141_508#
+ prbs_generator_syn_17/sky130_fd_sc_hs__nand2_1_47/B prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_29/X
+ prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_65/Y prbs_generator_syn_17/m3_13600_4701#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_1/a_437_503# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_67/a_1178_124#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_9/a_735_102# prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_13/a_132_392#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_15/a_1178_124# prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_15/A
+ prbs_generator_syn_17/sky130_fd_sc_hs__nand2_1_1/B prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_43/B
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_35/a_651_503# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_8/D
+ prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_29/A prbs_generator_syn_17/sky130_fd_sc_hs__nand2_1_7/B
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_13/a_735_102# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_47/a_696_458#
+ prbs_generator_syn_17/sky130_fd_sc_hs__nand2_1_31/B prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_51/a_735_102#
+ prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_59/X prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_35/a_1141_508#
+ prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_25/a_222_392# prbs_generator_syn_17/sky130_fd_sc_hs__sdlclkp_2_1/a_288_48#
+ prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_55/B prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_17/B
+ prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_43/A prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_7/A
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_65/a_1178_124# prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_59/Y
+ prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_41/X prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_21/a_230_79#
+ prbs_generator_syn_17/sky130_fd_sc_hs__nand2_1_57/a_117_74# prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_1/a_222_392#
+ prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_19/B prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_35/a_293_74#
+ prbs_generator_syn_17/sky130_fd_sc_hs__nand2_1_23/a_117_74# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_73/a_206_368#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_25/a_651_503# prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_1/a_138_385#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_37/a_696_458# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_67/a_544_485#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_43/a_27_74# prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_9/X
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_55/a_1034_424# prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_39/a_112_119#
+ prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_15/a_222_392# prbs_generator_syn_17/sky130_fd_sc_hs__conb_1_1/HI
+ prbs_generator_syn_17/sky130_fd_sc_hs__nand2_1_23/B prbs_generator_syn_17/sky130_fd_sc_hs__nand2_1_53/B
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_9/a_1178_124# prbs_generator_syn_17/sky130_fd_sc_hs__nor2b_1_4/A
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_47/a_1226_296# prbs_generator_syn_17/m3_13600_11045#
+ prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_17/X prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_29/a_376_368#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_5/a_544_485# prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_3/X
+ prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_31/a_132_392# prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_61/A
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_15/a_651_503# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_73/a_437_503#
+ prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_25/a_230_79# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_27/a_696_458#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_65/a_696_458# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_33/a_735_102#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_71/a_735_102# prbs_generator_syn_17/m3_13600_7263#
+ prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_43/a_222_392# prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_50/Y
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_8/a_1178_124# prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_53/B
+ prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_19/a_376_368# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_63/a_1178_124#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_4/a_696_458# prbs_generator_syn_17/sky130_fd_sc_hs__nor2b_1_4/a_278_368#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_13/a_1178_124# prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_61/a_132_392#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_53/a_206_368# prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_21/a_52_123#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_45/a_651_503# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_17/a_696_458#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_47/a_544_485# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_55/a_696_458#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_21/a_735_102# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_37/a_27_74#
+ prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_61/B prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_61/X
+ prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_59/a_112_119# prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_31/A
+ prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_33/a_222_392# prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_29/a_230_79#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_45/a_1226_296# prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_9/a_132_392#
+ prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_5/A prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_57/Y
+ prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_31/X prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_51/a_27_74#
+ prbs_generator_syn_17/sky130_fd_sc_hs__nor2b_1_8/a_27_112# prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_47/a_376_368#
+ prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_53/a_293_74# prbs_generator_syn_17/sky130_fd_sc_hs__nand2_1_43/a_117_74#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_8/a_735_102# prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_21/a_293_74#
+ prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_39/a_138_385# prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_63/Y
+ prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_51/a_132_392# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_43/a_206_368#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_53/a_437_503# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_37/a_544_485#
+ prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_57/X prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_53/a_1034_424#
+ prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_25/a_52_123# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_33/a_1141_508#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_63/Q prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_23/a_222_392#
+ prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_63/a_222_392# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_7/a_1178_124#
+ prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_53/X prbs_generator_syn_17/sky130_fd_sc_hs__nand2_2_5/Y
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_61/a_1178_124# prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_1/a_230_79#
+ prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_43/a_230_79# prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_11/a_230_79#
+ prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_41/a_132_392# prbs_generator_syn_17/sky130_fd_sc_hs__nand2_1_13/a_117_74#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_43/a_437_503# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_27/a_544_485#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_63/a_651_503# prbs_generator_syn_17/sky130_fd_sc_hs__nand2_1_7/a_117_74#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_35/a_696_458# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_65/a_544_485#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_51/a_1034_424# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_41/a_735_102#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_32/a_1141_508# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_49/a_1141_508#
+ prbs_generator_syn_17/sky130_fd_sc_hs__nand2_1_55/B prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_53/a_222_392#
+ prbs_generator_syn_17/sky130_fd_sc_hs__sdlclkp_2_1/a_114_112# prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_9/a_293_74#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_43/a_1226_296# prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_29/a_52_123#
+ prbs_generator_syn_17/sky130_fd_sc_hs__nand2_1_37/B prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_1/a_651_503#
+ prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_27/a_376_368# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_4/a_544_485#
+ prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_67/a_376_368# prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_27/X
+ prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_1/X prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_59/a_138_385#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_29/a_1178_124# prbs_generator_syn_17/m3_13600_2871#
+ prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_5/a_230_79# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_23/a_206_368#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_61/a_206_368# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_17/a_544_485#
+ prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_15/a_230_79# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_25/a_696_458#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_55/a_544_485# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_32/a_735_102#
+ prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_29/a_293_74# prbs_generator_syn_17/sky130_fd_sc_hs__nand2_1_17/a_117_74#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_69/a_1034_424# prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_29/a_112_119#
+ prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_37/X prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_31/B
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_19/a_1034_424# prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_33/A
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_9/a_206_368# prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_57/a_376_368#
+ prbs_generator_syn_17/sky130_fd_sc_hs__sdlclkp_2_1/a_706_317# prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_11/B
+ prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_1/a_52_123# prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_39/B
+ prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_21/a_132_392# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_13/a_206_368#
+ prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_43/a_52_123# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_51/a_206_368#
+ prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_47/X prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_23/a_437_503#
+ prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_11/a_52_123# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_61/a_437_503#
+ prbs_generator_syn_17/sky130_fd_sc_hs__nor2b_1_7/Y prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_51/A
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_15/a_696_458# prbs_generator_syn_17/sky130_fd_sc_hs__nor2b_1_5/Y
+ prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_9/a_230_79# prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_25/X
+ prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_19/a_112_119# prbs_generator_syn_17/sky130_fd_sc_hs__nand2_1_45/B
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_5/a_1178_124# prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_19/a_230_79#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_41/a_1226_296# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_59/a_1226_296#
+ prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_63/a_230_79# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_51/Q
+ prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_7/a_132_392# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_9/a_437_503#
+ prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_46/a_376_368# prbs_generator_syn_17/sky130_fd_sc_hs__nand2_1_33/a_117_74#
+ prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_11/a_293_74# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_27/a_1178_124#
+ prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_11/a_132_392# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_13/a_437_503#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_51/a_437_503# prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_5/a_52_123#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_35/a_544_485# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_73/a_651_503#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_45/a_696_458# prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_15/a_52_123#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_47/a_1141_508# prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_47/a_112_119#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_4/a_1178_124# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_17/a_1034_424#
+ prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_23/B prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_37/a_376_368#
+ prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_15/B prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_7/Y
+ prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_29/a_138_385# prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_33/a_230_79#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_25/a_1178_124# prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_47/a_293_74#
+ prbs_generator_syn_17/sky130_fd_sc_hs__nand2_1_37/a_117_74# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_33/a_206_368#
+ prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_15/a_293_74# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_71/a_206_368#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_25/a_544_485# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_67/a_1034_424#
+ prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_13/a_222_392# prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_9/a_52_123#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_15/a_1034_424# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_57/a_1226_296#
+ prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_19/a_52_123# prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_23/X
+ prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_63/a_52_123# prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_19/a_138_385#
+ prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_9/a_376_368# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_21/a_206_368#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_33/a_437_503# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_71/a_437_503#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_53/a_651_503# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_15/a_544_485#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_63/a_696_458# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_65/a_1034_424#
+ prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_19/a_293_74# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_45/a_1141_508#
+ prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_27/a_112_119# prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_67/a_112_119#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_1/a_1178_124# prbs_generator_syn_17/sky130_fd_sc_hs__conb_1_1/a_21_290#
+ prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_63/a_293_74# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_8/a_206_368#
+ prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_17/a_376_368# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_63/a_27_74#
+ prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_21/A prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_55/a_376_368#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_1/a_696_458# prbs_generator_syn_17/sky130_fd_sc_hs__nor2b_1_1/a_278_368#
+ prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_47/a_138_385# prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_33/a_52_123#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_9/a_1034_424# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_21/a_437_503#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_1/a_27_74# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_43/a_651_503#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_1/Q prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_45/a_544_485#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_69/a_735_102# prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_57/a_112_119#
+ prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_31/a_222_392# prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_13/A
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_55/a_1226_296# prbs_generator_syn_17/sky130_fd_sc_hs__nand2_2_5/a_27_74#
+ prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_53/a_230_79# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_8/a_437_503#
+ prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_67/a_293_74# prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_33/a_293_74#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_7/a_735_102# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_23/a_1178_124#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_41/a_206_368# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_8/a_1034_424#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_63/a_1034_424# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_59/a_735_102#
+ prbs_generator_syn_17/sky130_fd_sc_hs__nand2_1_5/B prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_43/a_1141_508#
+ prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_46/a_112_119# prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_61/a_222_392#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_13/a_1034_424# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_73/a_1178_124#
+ prbs_generator_syn_17/sky130_fd_sc_hs__nand2_1_27/B prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_13/B
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_57/a_27_74# prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_57/a_230_79#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_21/a_1178_124# prbs_generator_syn_17/sky130_fd_sc_hs__nor2b_1_1/a_27_112#
+ prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_27/a_138_385# prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_23/a_230_79#
+ prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_67/a_138_385# prbs_generator_syn_17/sky130_fd_sc_hs__nand2_1_41/B
+ prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_9/a_222_392# prbs_generator_syn_17/sky130_fd_sc_hs__nand2_1_27/a_117_74#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_32/a_206_368# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_23/a_651_503#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_41/a_437_503# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_73/a_27_74#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_61/a_651_503# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_63/a_544_485#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_49/a_735_102# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_73/a_696_458#
+ prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_37/a_112_119# prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_51/a_222_392#
+ prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_43/X prbs_generator_syn_17/sky130_fd_sc_hs__nand2_2_1/B
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_9/a_651_503# prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_53/a_52_123#
+ prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_49/X prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_25/a_376_368#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_1/a_544_485# prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_65/a_376_368#
+ prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_57/a_138_385# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_27/a_27_74#
+ prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_39/a_132_392# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_7/a_1034_424#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_13/a_651_503# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_32/a_437_503#
+ prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_27/a_230_79# prbs_generator_syn_17/m3_13600_12265#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_51/a_651_503# prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_59/B
+ prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_47/A prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_61/a_1034_424#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_41/a_1141_508# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_59/a_1141_508#
+ prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_41/a_222_392# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_53/a_1226_296#
+ prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_3/A prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_71/a_1178_124#
+ prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_9/a_112_119# prbs_generator_syn_17/sky130_fd_sc_hs__nand2_1_3/a_117_74#
+ prbs_generator_syn_17/m3_13600_8483# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_39/a_1178_124#
+ prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_57/a_52_123# prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_46/a_138_385#
+ prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_23/a_52_123# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_67/a_27_74#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_53/a_696_458# prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_17/a_112_119#
+ prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_11/A prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_55/a_112_119#
+ prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_1/A prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_51/a_1226_296#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_29/a_1034_424# prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_59/A
+ prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_23/A prbs_generator_syn_17/sky130_fd_sc_hs__nand2_1_39/B
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_5/a_27_74# prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_57/a_293_74#
+ prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_37/a_138_385# prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_59/a_132_392#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_33/a_651_503# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_71/a_651_503#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_43/a_696_458# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_73/a_544_485#
+ prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_27/a_52_123# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_57/a_1141_508#
+ prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_21/a_222_392# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_35/a_27_74#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_69/a_1226_296# prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_37/B
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_19/a_1226_296# prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_35/a_376_368#
+ prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_47/a_230_79# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_37/a_1178_124#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_5/a_1034_424# prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_49/a_132_392#
+ prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_7/a_222_392# prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_27/a_293_74#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_21/a_651_503# prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_9/a_138_385#
+ prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_11/a_222_392# prbs_generator_syn_17/m3_13600_14095#
+ prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_50/A prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_27/a_1034_424#
+ prbs_generator_syn_17/sky130_fd_sc_hs__nand2_1_13/B prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_8/a_651_503#
+ prbs_generator_syn_17/m3_13600_9703# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_35/a_1178_124#
+ prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_17/a_138_385# prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_55/a_138_385#
+ prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_7/a_230_79# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_4/a_1034_424#
+ prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_7/a_376_368# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_69/a_206_368#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_23/a_696_458# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_53/a_544_485#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_39/a_735_102# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_61/a_696_458#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_55/a_1141_508# prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_25/a_112_119#
+ prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_65/a_112_119# prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_43/a_293_74#
+ prbs_generator_syn_17/sky130_fd_sc_hs__nand2_1_57/B prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_25/a_1034_424#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_7/a_206_368# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_17/a_1226_296#
+ prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_15/a_376_368# prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_53/a_376_368#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_9/a_696_458# prbs_generator_syn_17/m3_13600_431#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_45/a_27_74# prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_47/a_52_123#
+ prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_29/a_132_392# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_59/a_206_368#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_69/a_437_503# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_41/a_651_503#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_43/a_544_485# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_13/a_696_458#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_29/a_735_102# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_51/a_696_458#
+ prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_61/Y prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_67/a_1226_296#
+ prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_5/a_132_392# prbs_generator_syn_17/sky130_fd_sc_hs__and2b_2_1/a_198_48#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_7/a_437_503# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_15/a_1226_296#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_69/a_27_74# prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_46/a_293_74#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_1/a_1034_424# prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_19/a_132_392#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_49/a_206_368# prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_7/a_52_123#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_59/a_437_503# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_32/a_651_503#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_7/a_27_74# prbs_generator_syn_17/sky130_fd_sc_hs__nand2_2_1/a_27_74#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_19/a_735_102# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_57/a_735_102#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_65/a_1226_296# prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_37/A
+ prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_33/a_376_368# prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_37/a_230_79#
+ prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_25/a_138_385# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_39/a_27_74#
+ prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_65/a_138_385# prbs_generator_syn_17/sky130_fd_sc_hs__nor2b_1_9/a_278_368#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_49/a_437_503# prbs_generator_syn_17/sky130_fd_sc_hs__and2b_2_1/a_505_74#
+ prbs_generator_syn_17/sky130_fd_sc_hs__nand2_1_51/a_117_74# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_23/a_544_485#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_33/a_696_458# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_61/a_544_485#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_9/a_1226_296# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_53/a_1141_508#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_71/a_696_458# prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_35/a_112_119#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_23/a_1034_424# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_9/a_544_485#
+ prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_63/a_376_368# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_33/a_1178_124#
+ prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_5/a_376_368# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_13/a_544_485#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_73/a_1034_424# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_21/a_696_458#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_51/a_544_485# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_8/a_1226_296#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_51/a_1141_508# prbs_generator_syn_17/sky130_fd_sc_hs__nand2_1_55/a_117_74#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_21/a_1034_424# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_63/a_1226_296#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_23/a_27_74# prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_7/a_112_119#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_13/a_1226_296# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_8/a_696_458#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_32/a_1178_124# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_49/a_1178_124#
+ prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_37/a_52_123# prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_27/a_132_392#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_71/Q prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_67/a_735_102#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_69/a_1141_508# prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_15/a_112_119#
+ prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_53/a_112_119# prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_39/a_222_392#
+ prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_55/a_230_79# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_19/a_1141_508#
+ prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_37/a_293_74# prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_43/a_376_368#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_5/a_735_102# prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_35/a_138_385#
+ prbs_generator_syn_17/sky130_fd_sc_hs__sdlclkp_2_1/a_114_424# prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_57/a_132_392#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_71/a_1034_424# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_7/a_1226_296#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_33/a_544_485# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_41/a_696_458#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_71/a_544_485# prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_21/B
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_61/a_1226_296# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_39/a_1034_424#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_17/a_27_74# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_9/a_27_74#
+ prbs_generator_syn_17/sky130_fd_sc_hs__nor2b_1_5/a_27_112# prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_47/a_132_392#
+ prbs_generator_syn_17/sky130_fd_sc_hs__nor2b_1_8/a_278_368# prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_9/B
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_39/a_206_368# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_33/a_27_74#
+ prbs_generator_syn_17/sky130_fd_sc_hs__nand2_1_41/a_117_74# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_69/a_651_503#
+ prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_51/a_293_74# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_21/a_544_485#
+ prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_7/a_138_385# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_32/a_696_458#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_47/a_735_102# prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_33/a_112_119#
+ prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_59/a_222_392# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_17/a_1141_508#
+ prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_55/a_52_123# prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_3/a_293_74#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_7/a_651_503# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_29/a_1226_296#
+ prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_23/a_376_368# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_8/a_544_485#
+ prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_47/B prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_47/a_1178_124#
+ prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_15/a_138_385# prbs_generator_syn_17/sky130_fd_sc_hs__sdlclkp_2_1/a_1195_374#
+ prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_53/a_138_385# prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_37/a_132_392#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_29/a_206_368# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_39/a_437_503#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_59/a_651_503# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_37/a_735_102#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_67/a_1141_508# prbs_generator_syn_17/sky130_fd_sc_hs__and2b_2_1/a_27_74#
+ prbs_generator_syn_17/sky130_fd_sc_hs__conb_1_1/a_165_290# prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_55/a_293_74#
+ prbs_generator_syn_17/sky130_fd_sc_hs__nand2_1_45/a_117_74# prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_63/a_112_119#
+ prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_49/a_222_392# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_37/a_1034_424#
+ prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_23/a_293_74# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_15/a_1141_508#
+ prbs_generator_syn_17/sky130_fd_sc_hs__nand2_1_5/a_117_74# prbs_generator_syn_17/m3_13600_13485#
+ prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_5/a_112_119# prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_13/a_376_368#
+ prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_51/a_376_368# prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_7/a_293_74#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_19/a_206_368# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_57/a_206_368#
+ prbs_generator_syn_17/sky130_fd_sc_hs__sdlclkp_2_1/a_318_74# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_29/a_437_503#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_49/a_651_503# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_25/a_27_74#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_5/a_1226_296# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_41/a_544_485#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_27/a_735_102# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_65/a_1141_508#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_65/a_735_102# prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_3/a_230_79#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_35/a_1034_424# prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_13/a_230_79#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_41/a_27_74# prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_3/a_132_392#
+ prbs_generator_syn_17/sky130_fd_sc_hs__nand2_1_49/a_117_74# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_27/a_1226_296#
+ prbs_generator_syn_17/sky130_fd_sc_hs__nand2_1_15/a_117_74# prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_41/a_376_368#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_45/a_1178_124# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_4/a_735_102#
+ prbs_generator_syn_17/sky130_fd_sc_hs__nand2_1_9/a_117_74# prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_33/a_138_385#
+ prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_17/a_132_392# prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_55/a_132_392#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_9/a_1141_508# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_19/a_437_503#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_57/a_437_503# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_4/a_1226_296#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_32/a_544_485# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_17/a_735_102#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_55/a_735_102# prbs_generator_syn_17/m3_13600_2261#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_65/a_27_74# prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_29/a_222_392#
+ prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_43/a_112_119# prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_19/X
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_25/a_1226_296# prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_31/a_376_368#
+ prbs_generator_syn_17/sky130_fd_sc_hs__or2_1_1/a_63_368# prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_17/a_230_79#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_4/a_27_74# prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_61/a_230_79#
+ prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_63/a_138_385# prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_5/a_222_392#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_8/a_1141_508# prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_41/a_293_74#
+ prbs_generator_syn_17/sky130_fd_sc_hs__nand2_1_31/a_117_74# prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_5/a_138_385#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_63/a_1141_508# prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_19/a_222_392#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_13/a_1141_508# prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_3/a_52_123#
+ prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_13/a_52_123# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_43/a_1178_124#
+ prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_61/a_376_368# prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_35/a_132_392#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_67/a_206_368# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_1/a_1226_296#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_69/a_696_458# prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_31/a_230_79#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_35/a_735_102# prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_23/a_112_119#
+ prbs_generator_syn_17/sky130_fd_sc_hs__nand2_1_35/a_117_74# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_59/a_27_74#
+ prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_13/a_293_74# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_5/a_206_368#
+ prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_50/a_376_368# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_7/a_696_458#
+ prbs_generator_syn_17/sky130_fd_sc_hs__nor2b_1_7/a_278_368# prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_17/a_52_123#
+ prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_43/a_138_385# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_7/a_1141_508#
+ prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_61/a_52_123# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_67/a_437_503#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_61/a_1141_508# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_25/a_735_102#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_59/a_696_458# prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_13/a_112_119#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_33/a_1034_424# prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_51/a_112_119#
+ prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_35/a_230_79# prbs_generator_syn_17/m3_13600_4091#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_23/a_1226_296# prbs_generator_syn_17/sky130_fd_sc_hs__nand2_1_39/a_117_74#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_29/a_27_74# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_5/a_437_503#
+ prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_17/a_293_74# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_41/a_1178_124#
+ prbs_generator_syn_17/sky130_fd_sc_hs__or2_1_1/a_152_368# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_59/a_1178_124#
+ prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_61/a_293_74# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_47/a_206_368#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_39/a_651_503# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_49/a_696_458#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_15/a_735_102# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_32/a_1034_424#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_73/a_1226_296# prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_27/a_222_392#
+ prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_41/a_112_119# prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_31/a_52_123#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_49/a_1034_424# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_29/a_1141_508#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_21/a_1226_296# prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_39/a_230_79#
+ prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_23/a_138_385# prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_51/a_230_79#
+ prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_45/a_132_392# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_37/a_206_368#
+ prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_65/a_293_74# prbs_generator_syn_17/sky130_fd_sc_hs__nand2_1_53/a_117_74#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_47/a_437_503# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_29/a_651_503#
+ prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_31/a_293_74# prbs_generator_syn_17/sky130_fd_sc_hs__nand2_1_21/a_117_74#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_69/a_544_485# prbs_generator_syn_17/sky130_fd_sc_hs__clkbuf_16_1/a_114_74#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_45/a_735_102# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_13/a_27_74#
+ prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_31/a_112_119# prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_57/a_222_392#
+ prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_35/a_52_123# prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_21/a_376_368#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_7/a_544_485# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_57/a_1178_124#
+ prbs_generator_syn_17/m3_13600_6043# prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_13/a_138_385#
+ prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_51/a_138_385# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_5/a_1141_508#
+ prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_3/a_376_368# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_27/a_206_368#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_65/a_206_368# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_37/a_437_503#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_19/a_651_503# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_57/a_651_503#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_59/a_544_485# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_71/a_1226_296#
+ prbs_generator_syn_17/sky130_fd_sc_hs__nand2_1_25/a_117_74# prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_61/a_112_119#
+ prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_47/a_222_392# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_27/a_1141_508#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_53/a_27_74# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_4/a_206_368#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_39/a_1226_296# prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_11/a_376_368#
+ prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_39/a_52_123# prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_41/a_138_385#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_4/a_1141_508# prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_25/a_132_392#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_17/a_206_368# prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_41/A
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_55/a_206_368# prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_51/a_52_123#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_27/a_437_503# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_65/a_437_503#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_49/a_544_485# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_63/a_735_102#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_47/a_1034_424# prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_50/a_112_119#
+ prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_37/a_222_392# prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_59/a_230_79#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_25/a_1141_508# prbs_generator_syn_17/sky130_fd_sc_hs__nor2b_1_4/a_27_112#
+ prbs_generator_syn_17/sky130_fd_sc_hs__sdlclkp_2_1/a_685_81# prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_1/a_132_392#
+ prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_39/a_293_74# prbs_generator_syn_17/sky130_fd_sc_hs__nand2_1_29/a_117_74#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_4/a_437_503# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_55/a_1178_124#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_21/a_27_74# prbs_generator_syn_17/m3_13600_12875#
+ prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_50/a_293_74# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_1/a_735_102#
+ prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_31/a_138_385# prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_15/a_132_392#
+ prbs_generator_syn_17/sky130_fd_sc_hs__nand2_1_1/a_117_74# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_17/a_437_503#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_55/a_437_503# prbs_generator_syn
Xprbs_generator_syn_27 prbs_generator_syn_31/clk prbs_generator_syn_27/rst prbs_generator_syn_27/cke
+ sky130_fd_sc_hs__conb_1_257/LO sky130_fd_sc_hs__conb_1_257/LO sky130_fd_sc_hs__conb_1_257/LO
+ sky130_fd_sc_hs__conb_1_257/LO sky130_fd_sc_hs__conb_1_257/LO sky130_fd_sc_hs__conb_1_257/HI
+ sky130_fd_sc_hs__conb_1_257/HI sky130_fd_sc_hs__conb_1_257/HI sky130_fd_sc_hs__conb_1_257/HI
+ sky130_fd_sc_hs__conb_1_257/HI sky130_fd_sc_hs__conb_1_257/HI prbs_generator_syn_27/cke
+ prbs_generator_syn_27/cke prbs_generator_syn_27/cke prbs_generator_syn_27/cke prbs_generator_syn_27/cke
+ prbs_generator_syn_27/eqn[31] prbs_generator_syn_27/cke prbs_generator_syn_31/eqn[9]
+ prbs_generator_syn_31/eqn[20] prbs_generator_syn_31/eqn[21] prbs_generator_syn_31/eqn[20]
+ prbs_generator_syn_31/eqn[21] sky130_fd_sc_hs__conb_1_247/HI prbs_generator_syn_31/eqn[28]
+ sky130_fd_sc_hs__conb_1_247/HI sky130_fd_sc_hs__conb_1_247/HI prbs_generator_syn_31/eqn[30]
+ prbs_generator_syn_31/eqn[30] sky130_fd_sc_hs__conb_1_259/HI sky130_fd_sc_hs__conb_1_259/HI
+ prbs_generator_syn_31/eqn[30] prbs_generator_syn_27/eqn[31] prbs_generator_syn_27/eqn[30]
+ prbs_generator_syn_27/eqn[30] prbs_generator_syn_27/eqn[28] prbs_generator_syn_27/eqn[28]
+ prbs_generator_syn_27/eqn[28] prbs_generator_syn_27/eqn[28] prbs_generator_syn_27/eqn[28]
+ prbs_generator_syn_27/eqn[28] prbs_generator_syn_27/eqn[22] prbs_generator_syn_27/eqn[22]
+ prbs_generator_syn_27/eqn[20] prbs_generator_syn_27/eqn[22] prbs_generator_syn_27/eqn[22]
+ prbs_generator_syn_27/eqn[22] prbs_generator_syn_27/eqn[22] prbs_generator_syn_27/eqn[22]
+ prbs_generator_syn_27/eqn[9] prbs_generator_syn_27/eqn[9] prbs_generator_syn_27/eqn[9]
+ prbs_generator_syn_27/eqn[9] prbs_generator_syn_27/eqn[9] prbs_generator_syn_27/eqn[9]
+ prbs_generator_syn_27/eqn[8] prbs_generator_syn_27/eqn[8] prbs_generator_syn_27/eqn[8]
+ prbs_generator_syn_27/eqn[8] prbs_generator_syn_27/eqn[8] prbs_generator_syn_27/eqn[8]
+ prbs_generator_syn_27/eqn[8] prbs_generator_syn_27/eqn[1] prbs_generator_syn_31/eqn[9]
+ prbs_generator_syn_27/inj_err prbs_generator_syn_27/eqn[31] prbs_generator_syn_27/eqn[31]
+ hr_16t4_mux_top_1/din[4] DVSS: DVDD: prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_1/a_293_74#
+ prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_15/X prbs_generator_syn_27/sky130_fd_sc_hs__nand2_1_35/B
+ prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_51/Y prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_9/A
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_9/CLK prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_47/a_27_74#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_37/a_1226_296# prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_3/B
+ prbs_generator_syn_27/sky130_fd_sc_hs__nor2b_1_7/a_27_112# prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_29/B
+ prbs_generator_syn_27/sky130_fd_sc_hs__sdlclkp_2_1/a_580_74# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_1/a_1141_508#
+ prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_5/Y prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_41/a_230_79#
+ prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_61/a_138_385# prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_43/a_132_392#
+ prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_3/a_222_392# prbs_generator_syn_27/sky130_fd_sc_hs__nor2b_1_9/a_27_112#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_61/a_27_74# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_35/a_206_368#
+ prbs_generator_syn_27/sky130_fd_sc_hs__nand2_2_3/Y prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_25/B
+ prbs_generator_syn_27/sky130_fd_sc_hs__nand2_1_11/a_117_74# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_67/a_651_503#
+ prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_45/X prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_39/a_696_458#
+ prbs_generator_syn_27/sky130_fd_sc_hs__sdlclkp_2_1/a_1198_74# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_45/a_1034_424#
+ prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_17/a_222_392# prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_55/a_222_392#
+ prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_53/Y prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_35/A
+ prbs_generator_syn_27/m3_13600_1651# prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_59/a_52_123#
+ prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_5/a_293_74# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_35/a_1226_296#
+ prbs_generator_syn_27/sky130_fd_sc_hs__nand2_1_51/B prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_5/a_651_503#
+ prbs_generator_syn_27/sky130_fd_sc_hs__nand2_1_21/B prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_8/a_27_74#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_15/a_27_74# prbs_generator_syn_27/sky130_fd_sc_hs__and2b_2_1/X
+ prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_13/X prbs_generator_syn_27/sky130_fd_sc_hs__nand2_2_3/a_27_74#
+ prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_50/a_138_385# prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_33/a_132_392#
+ prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_1/a_376_368# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_25/a_206_368#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_35/a_437_503# prbs_generator_syn_27/sky130_fd_sc_hs__sdlclkp_2_1/a_708_451#
+ prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_45/a_230_79# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_29/a_696_458#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_32/a_27_74# prbs_generator_syn_27/sky130_fd_sc_hs__nor2b_1_4/Y
+ prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_59/a_293_74# prbs_generator_syn_27/sky130_fd_sc_hs__nand2_1_47/a_117_74#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_73/a_735_102# prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_21/a_112_119#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_23/a_1141_508# prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_25/a_293_74#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_7/Q prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_3/a_112_119#
+ prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_35/B prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_51/X
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_53/a_1178_124# prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_23/a_132_392#
+ prbs_generator_syn_27/sky130_fd_sc_hs__nand2_1_3/B prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_15/a_206_368#
+ prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_63/a_132_392# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_55/a_27_74#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_25/a_437_503# prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_41/a_52_123#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_47/a_651_503# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_73/a_1141_508#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_19/a_696_458# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_57/a_696_458#
+ prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_7/X prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_43/a_1034_424#
+ prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_55/A prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_11/a_112_119#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_21/a_1141_508# prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_35/a_222_392#
+ prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_49/a_230_79# prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_67/Y
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_71/a_27_74# prbs_generator_syn_27/sky130_fd_sc_hs__nand2_1_33/B
+ prbs_generator_syn_27/sky130_fd_sc_hs__conb_1_1/LO prbs_generator_syn_27/sky130_fd_sc_hs__nand2_1_19/a_117_74#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_51/a_1178_124# prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_33/X
+ prbs_generator_syn_27/sky130_fd_sc_hs__nand2_1_29/B prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_41/Y
+ prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_53/a_132_392# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_45/a_206_368#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_15/a_437_503# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_37/a_651_503#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_39/a_544_485# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_53/a_735_102#
+ prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_45/a_52_123# prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_1/B
+ prbs_generator_syn_27/sky130_fd_sc_hs__nand2_2_3/B prbs_generator_syn_27/sky130_fd_sc_hs__clkbuf_16_1/A
+ prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_21/X prbs_generator_syn_27/sky130_fd_sc_hs__nand2_1_25/B
+ prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_39/a_376_368# prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_63/X
+ prbs_generator_syn_27/m3_13600_3481# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_69/a_1178_124#
+ prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_21/a_138_385# prbs_generator_syn_27/sky130_fd_sc_hs__nor2b_1_8/Y
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_19/a_1178_124# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_49/a_27_74#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_45/a_437_503# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_27/a_651_503#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_71/a_1141_508# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_65/a_651_503#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_29/a_544_485# prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_3/a_138_385#
+ prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_55/X prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_43/a_735_102#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_41/a_1034_424# prbs_generator_syn_27/sky130_fd_sc_hs__nand2_1_9/B
+ prbs_generator_syn_27/sky130_fd_sc_hs__nor2b_1_9/Y prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_59/a_1034_424#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_39/a_1141_508# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_33/a_1226_296#
+ prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_49/a_52_123# prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_47/Y
+ prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_43/Y prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_4/a_651_503#
+ prbs_generator_syn_27/sky130_fd_sc_hs__nand2_1_49/B prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_19/A
+ prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_11/a_138_385# prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_5/X
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_63/a_206_368# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_17/a_651_503#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_19/a_544_485# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_55/a_651_503#
+ prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_9/Y prbs_generator_syn_27/sky130_fd_sc_hs__nand2_1_17/B
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_57/a_544_485# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_67/a_696_458#
+ prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_35/X prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_19/a_27_74#
+ prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_45/a_222_392# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_32/a_1226_296#
+ prbs_generator_syn_27/sky130_fd_sc_hs__nand2_1_43/B prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_25/A
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_1/a_206_368# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_49/a_1226_296#
+ prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_1/a_112_119# prbs_generator_syn_27/sky130_fd_sc_hs__or2_1_1/X
+ prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_59/a_376_368# prbs_generator_syn_27/sky130_fd_sc_hs__nand2_1_19/B
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_5/a_696_458# prbs_generator_syn_27/sky130_fd_sc_hs__nor2b_1_1/Y
+ prbs_generator_syn_27/sky130_fd_sc_hs__nor2b_1_5/a_278_368# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_17/a_1178_124#
+ prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_39/X prbs_generator_syn_27/m3_13600_5433#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_63/a_437_503# prbs_generator_syn_27/sky130_fd_sc_hs__nand2_2_5/B
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_23/a_735_102# prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_53/A
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_61/a_735_102# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_57/a_1034_424#
+ prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_63/B prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_37/a_1141_508#
+ prbs_generator_syn_27/sky130_fd_sc_hs__nand2_1_47/B prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_29/X
+ prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_65/Y prbs_generator_syn_27/m3_13600_4701#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_1/a_437_503# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_67/a_1178_124#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_9/a_735_102# prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_13/a_132_392#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_15/a_1178_124# prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_15/A
+ prbs_generator_syn_27/sky130_fd_sc_hs__nand2_1_1/B prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_43/B
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_35/a_651_503# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_8/D
+ prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_29/A prbs_generator_syn_27/sky130_fd_sc_hs__nand2_1_7/B
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_13/a_735_102# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_47/a_696_458#
+ prbs_generator_syn_27/sky130_fd_sc_hs__nand2_1_31/B prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_51/a_735_102#
+ prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_59/X prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_35/a_1141_508#
+ prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_25/a_222_392# prbs_generator_syn_27/sky130_fd_sc_hs__sdlclkp_2_1/a_288_48#
+ prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_55/B prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_17/B
+ prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_43/A prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_7/A
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_65/a_1178_124# prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_59/Y
+ prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_41/X prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_21/a_230_79#
+ prbs_generator_syn_27/sky130_fd_sc_hs__nand2_1_57/a_117_74# prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_1/a_222_392#
+ prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_19/B prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_35/a_293_74#
+ prbs_generator_syn_27/sky130_fd_sc_hs__nand2_1_23/a_117_74# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_73/a_206_368#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_25/a_651_503# prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_1/a_138_385#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_37/a_696_458# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_67/a_544_485#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_43/a_27_74# prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_9/X
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_55/a_1034_424# prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_39/a_112_119#
+ prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_15/a_222_392# prbs_generator_syn_27/sky130_fd_sc_hs__conb_1_1/HI
+ prbs_generator_syn_27/sky130_fd_sc_hs__nand2_1_23/B prbs_generator_syn_27/sky130_fd_sc_hs__nand2_1_53/B
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_9/a_1178_124# prbs_generator_syn_27/sky130_fd_sc_hs__nor2b_1_4/A
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_47/a_1226_296# prbs_generator_syn_27/m3_13600_11045#
+ prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_17/X prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_29/a_376_368#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_5/a_544_485# prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_3/X
+ prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_31/a_132_392# prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_61/A
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_15/a_651_503# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_73/a_437_503#
+ prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_25/a_230_79# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_27/a_696_458#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_65/a_696_458# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_33/a_735_102#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_71/a_735_102# prbs_generator_syn_27/m3_13600_7263#
+ prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_43/a_222_392# prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_50/Y
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_8/a_1178_124# prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_53/B
+ prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_19/a_376_368# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_63/a_1178_124#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_4/a_696_458# prbs_generator_syn_27/sky130_fd_sc_hs__nor2b_1_4/a_278_368#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_13/a_1178_124# prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_61/a_132_392#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_53/a_206_368# prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_21/a_52_123#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_45/a_651_503# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_17/a_696_458#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_47/a_544_485# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_55/a_696_458#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_21/a_735_102# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_37/a_27_74#
+ prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_61/B prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_61/X
+ prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_59/a_112_119# prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_31/A
+ prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_33/a_222_392# prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_29/a_230_79#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_45/a_1226_296# prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_9/a_132_392#
+ prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_5/A prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_57/Y
+ prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_31/X prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_51/a_27_74#
+ prbs_generator_syn_27/sky130_fd_sc_hs__nor2b_1_8/a_27_112# prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_47/a_376_368#
+ prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_53/a_293_74# prbs_generator_syn_27/sky130_fd_sc_hs__nand2_1_43/a_117_74#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_8/a_735_102# prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_21/a_293_74#
+ prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_39/a_138_385# prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_63/Y
+ prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_51/a_132_392# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_43/a_206_368#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_53/a_437_503# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_37/a_544_485#
+ prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_57/X prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_53/a_1034_424#
+ prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_25/a_52_123# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_33/a_1141_508#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_63/Q prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_23/a_222_392#
+ prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_63/a_222_392# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_7/a_1178_124#
+ prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_53/X prbs_generator_syn_27/sky130_fd_sc_hs__nand2_2_5/Y
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_61/a_1178_124# prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_1/a_230_79#
+ prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_43/a_230_79# prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_11/a_230_79#
+ prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_41/a_132_392# prbs_generator_syn_27/sky130_fd_sc_hs__nand2_1_13/a_117_74#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_43/a_437_503# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_27/a_544_485#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_63/a_651_503# prbs_generator_syn_27/sky130_fd_sc_hs__nand2_1_7/a_117_74#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_35/a_696_458# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_65/a_544_485#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_51/a_1034_424# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_41/a_735_102#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_32/a_1141_508# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_49/a_1141_508#
+ prbs_generator_syn_27/sky130_fd_sc_hs__nand2_1_55/B prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_53/a_222_392#
+ prbs_generator_syn_27/sky130_fd_sc_hs__sdlclkp_2_1/a_114_112# prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_9/a_293_74#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_43/a_1226_296# prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_29/a_52_123#
+ prbs_generator_syn_27/sky130_fd_sc_hs__nand2_1_37/B prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_1/a_651_503#
+ prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_27/a_376_368# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_4/a_544_485#
+ prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_67/a_376_368# prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_27/X
+ prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_1/X prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_59/a_138_385#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_29/a_1178_124# prbs_generator_syn_27/m3_13600_2871#
+ prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_5/a_230_79# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_23/a_206_368#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_61/a_206_368# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_17/a_544_485#
+ prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_15/a_230_79# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_25/a_696_458#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_55/a_544_485# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_32/a_735_102#
+ prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_29/a_293_74# prbs_generator_syn_27/sky130_fd_sc_hs__nand2_1_17/a_117_74#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_69/a_1034_424# prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_29/a_112_119#
+ prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_37/X prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_31/B
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_19/a_1034_424# prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_33/A
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_9/a_206_368# prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_57/a_376_368#
+ prbs_generator_syn_27/sky130_fd_sc_hs__sdlclkp_2_1/a_706_317# prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_11/B
+ prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_1/a_52_123# prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_39/B
+ prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_21/a_132_392# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_13/a_206_368#
+ prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_43/a_52_123# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_51/a_206_368#
+ prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_47/X prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_23/a_437_503#
+ prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_11/a_52_123# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_61/a_437_503#
+ prbs_generator_syn_27/sky130_fd_sc_hs__nor2b_1_7/Y prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_51/A
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_15/a_696_458# prbs_generator_syn_27/sky130_fd_sc_hs__nor2b_1_5/Y
+ prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_9/a_230_79# prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_25/X
+ prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_19/a_112_119# prbs_generator_syn_27/sky130_fd_sc_hs__nand2_1_45/B
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_5/a_1178_124# prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_19/a_230_79#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_41/a_1226_296# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_59/a_1226_296#
+ prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_63/a_230_79# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_51/Q
+ prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_7/a_132_392# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_9/a_437_503#
+ prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_46/a_376_368# prbs_generator_syn_27/sky130_fd_sc_hs__nand2_1_33/a_117_74#
+ prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_11/a_293_74# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_27/a_1178_124#
+ prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_11/a_132_392# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_13/a_437_503#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_51/a_437_503# prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_5/a_52_123#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_35/a_544_485# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_73/a_651_503#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_45/a_696_458# prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_15/a_52_123#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_47/a_1141_508# prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_47/a_112_119#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_4/a_1178_124# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_17/a_1034_424#
+ prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_23/B prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_37/a_376_368#
+ prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_15/B prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_7/Y
+ prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_29/a_138_385# prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_33/a_230_79#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_25/a_1178_124# prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_47/a_293_74#
+ prbs_generator_syn_27/sky130_fd_sc_hs__nand2_1_37/a_117_74# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_33/a_206_368#
+ prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_15/a_293_74# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_71/a_206_368#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_25/a_544_485# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_67/a_1034_424#
+ prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_13/a_222_392# prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_9/a_52_123#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_15/a_1034_424# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_57/a_1226_296#
+ prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_19/a_52_123# prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_23/X
+ prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_63/a_52_123# prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_19/a_138_385#
+ prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_9/a_376_368# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_21/a_206_368#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_33/a_437_503# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_71/a_437_503#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_53/a_651_503# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_15/a_544_485#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_63/a_696_458# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_65/a_1034_424#
+ prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_19/a_293_74# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_45/a_1141_508#
+ prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_27/a_112_119# prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_67/a_112_119#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_1/a_1178_124# prbs_generator_syn_27/sky130_fd_sc_hs__conb_1_1/a_21_290#
+ prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_63/a_293_74# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_8/a_206_368#
+ prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_17/a_376_368# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_63/a_27_74#
+ prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_21/A prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_55/a_376_368#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_1/a_696_458# prbs_generator_syn_27/sky130_fd_sc_hs__nor2b_1_1/a_278_368#
+ prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_47/a_138_385# prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_33/a_52_123#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_9/a_1034_424# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_21/a_437_503#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_1/a_27_74# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_43/a_651_503#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_1/Q prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_45/a_544_485#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_69/a_735_102# prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_57/a_112_119#
+ prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_31/a_222_392# prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_13/A
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_55/a_1226_296# prbs_generator_syn_27/sky130_fd_sc_hs__nand2_2_5/a_27_74#
+ prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_53/a_230_79# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_8/a_437_503#
+ prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_67/a_293_74# prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_33/a_293_74#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_7/a_735_102# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_23/a_1178_124#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_41/a_206_368# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_8/a_1034_424#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_63/a_1034_424# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_59/a_735_102#
+ prbs_generator_syn_27/sky130_fd_sc_hs__nand2_1_5/B prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_43/a_1141_508#
+ prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_46/a_112_119# prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_61/a_222_392#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_13/a_1034_424# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_73/a_1178_124#
+ prbs_generator_syn_27/sky130_fd_sc_hs__nand2_1_27/B prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_13/B
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_57/a_27_74# prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_57/a_230_79#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_21/a_1178_124# prbs_generator_syn_27/sky130_fd_sc_hs__nor2b_1_1/a_27_112#
+ prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_27/a_138_385# prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_23/a_230_79#
+ prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_67/a_138_385# prbs_generator_syn_27/sky130_fd_sc_hs__nand2_1_41/B
+ prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_9/a_222_392# prbs_generator_syn_27/sky130_fd_sc_hs__nand2_1_27/a_117_74#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_32/a_206_368# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_23/a_651_503#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_41/a_437_503# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_73/a_27_74#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_61/a_651_503# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_63/a_544_485#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_49/a_735_102# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_73/a_696_458#
+ prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_37/a_112_119# prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_51/a_222_392#
+ prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_43/X prbs_generator_syn_27/sky130_fd_sc_hs__nand2_2_1/B
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_9/a_651_503# prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_53/a_52_123#
+ prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_49/X prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_25/a_376_368#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_1/a_544_485# prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_65/a_376_368#
+ prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_57/a_138_385# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_27/a_27_74#
+ prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_39/a_132_392# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_7/a_1034_424#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_13/a_651_503# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_32/a_437_503#
+ prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_27/a_230_79# prbs_generator_syn_27/m3_13600_12265#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_51/a_651_503# prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_59/B
+ prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_47/A prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_61/a_1034_424#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_41/a_1141_508# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_59/a_1141_508#
+ prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_41/a_222_392# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_53/a_1226_296#
+ prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_3/A prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_71/a_1178_124#
+ prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_9/a_112_119# prbs_generator_syn_27/sky130_fd_sc_hs__nand2_1_3/a_117_74#
+ prbs_generator_syn_27/m3_13600_8483# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_39/a_1178_124#
+ prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_57/a_52_123# prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_46/a_138_385#
+ prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_23/a_52_123# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_67/a_27_74#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_53/a_696_458# prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_17/a_112_119#
+ prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_11/A prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_55/a_112_119#
+ prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_1/A prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_51/a_1226_296#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_29/a_1034_424# prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_59/A
+ prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_23/A prbs_generator_syn_27/sky130_fd_sc_hs__nand2_1_39/B
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_5/a_27_74# prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_57/a_293_74#
+ prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_37/a_138_385# prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_59/a_132_392#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_33/a_651_503# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_71/a_651_503#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_43/a_696_458# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_73/a_544_485#
+ prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_27/a_52_123# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_57/a_1141_508#
+ prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_21/a_222_392# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_35/a_27_74#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_69/a_1226_296# prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_37/B
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_19/a_1226_296# prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_35/a_376_368#
+ prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_47/a_230_79# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_37/a_1178_124#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_5/a_1034_424# prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_49/a_132_392#
+ prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_7/a_222_392# prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_27/a_293_74#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_21/a_651_503# prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_9/a_138_385#
+ prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_11/a_222_392# prbs_generator_syn_27/m3_13600_14095#
+ prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_50/A prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_27/a_1034_424#
+ prbs_generator_syn_27/sky130_fd_sc_hs__nand2_1_13/B prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_8/a_651_503#
+ prbs_generator_syn_27/m3_13600_9703# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_35/a_1178_124#
+ prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_17/a_138_385# prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_55/a_138_385#
+ prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_7/a_230_79# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_4/a_1034_424#
+ prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_7/a_376_368# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_69/a_206_368#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_23/a_696_458# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_53/a_544_485#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_39/a_735_102# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_61/a_696_458#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_55/a_1141_508# prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_25/a_112_119#
+ prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_65/a_112_119# prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_43/a_293_74#
+ prbs_generator_syn_27/sky130_fd_sc_hs__nand2_1_57/B prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_25/a_1034_424#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_7/a_206_368# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_17/a_1226_296#
+ prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_15/a_376_368# prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_53/a_376_368#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_9/a_696_458# prbs_generator_syn_27/m3_13600_431#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_45/a_27_74# prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_47/a_52_123#
+ prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_29/a_132_392# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_59/a_206_368#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_69/a_437_503# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_41/a_651_503#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_43/a_544_485# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_13/a_696_458#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_29/a_735_102# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_51/a_696_458#
+ prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_61/Y prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_67/a_1226_296#
+ prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_5/a_132_392# prbs_generator_syn_27/sky130_fd_sc_hs__and2b_2_1/a_198_48#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_7/a_437_503# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_15/a_1226_296#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_69/a_27_74# prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_46/a_293_74#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_1/a_1034_424# prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_19/a_132_392#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_49/a_206_368# prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_7/a_52_123#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_59/a_437_503# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_32/a_651_503#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_7/a_27_74# prbs_generator_syn_27/sky130_fd_sc_hs__nand2_2_1/a_27_74#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_19/a_735_102# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_57/a_735_102#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_65/a_1226_296# prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_37/A
+ prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_33/a_376_368# prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_37/a_230_79#
+ prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_25/a_138_385# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_39/a_27_74#
+ prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_65/a_138_385# prbs_generator_syn_27/sky130_fd_sc_hs__nor2b_1_9/a_278_368#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_49/a_437_503# prbs_generator_syn_27/sky130_fd_sc_hs__and2b_2_1/a_505_74#
+ prbs_generator_syn_27/sky130_fd_sc_hs__nand2_1_51/a_117_74# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_23/a_544_485#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_33/a_696_458# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_61/a_544_485#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_9/a_1226_296# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_53/a_1141_508#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_71/a_696_458# prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_35/a_112_119#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_23/a_1034_424# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_9/a_544_485#
+ prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_63/a_376_368# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_33/a_1178_124#
+ prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_5/a_376_368# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_13/a_544_485#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_73/a_1034_424# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_21/a_696_458#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_51/a_544_485# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_8/a_1226_296#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_51/a_1141_508# prbs_generator_syn_27/sky130_fd_sc_hs__nand2_1_55/a_117_74#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_21/a_1034_424# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_63/a_1226_296#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_23/a_27_74# prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_7/a_112_119#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_13/a_1226_296# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_8/a_696_458#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_32/a_1178_124# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_49/a_1178_124#
+ prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_37/a_52_123# prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_27/a_132_392#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_71/Q prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_67/a_735_102#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_69/a_1141_508# prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_15/a_112_119#
+ prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_53/a_112_119# prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_39/a_222_392#
+ prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_55/a_230_79# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_19/a_1141_508#
+ prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_37/a_293_74# prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_43/a_376_368#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_5/a_735_102# prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_35/a_138_385#
+ prbs_generator_syn_27/sky130_fd_sc_hs__sdlclkp_2_1/a_114_424# prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_57/a_132_392#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_71/a_1034_424# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_7/a_1226_296#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_33/a_544_485# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_41/a_696_458#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_71/a_544_485# prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_21/B
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_61/a_1226_296# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_39/a_1034_424#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_17/a_27_74# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_9/a_27_74#
+ prbs_generator_syn_27/sky130_fd_sc_hs__nor2b_1_5/a_27_112# prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_47/a_132_392#
+ prbs_generator_syn_27/sky130_fd_sc_hs__nor2b_1_8/a_278_368# prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_9/B
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_39/a_206_368# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_33/a_27_74#
+ prbs_generator_syn_27/sky130_fd_sc_hs__nand2_1_41/a_117_74# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_69/a_651_503#
+ prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_51/a_293_74# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_21/a_544_485#
+ prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_7/a_138_385# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_32/a_696_458#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_47/a_735_102# prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_33/a_112_119#
+ prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_59/a_222_392# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_17/a_1141_508#
+ prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_55/a_52_123# prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_3/a_293_74#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_7/a_651_503# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_29/a_1226_296#
+ prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_23/a_376_368# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_8/a_544_485#
+ prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_47/B prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_47/a_1178_124#
+ prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_15/a_138_385# prbs_generator_syn_27/sky130_fd_sc_hs__sdlclkp_2_1/a_1195_374#
+ prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_53/a_138_385# prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_37/a_132_392#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_29/a_206_368# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_39/a_437_503#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_59/a_651_503# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_37/a_735_102#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_67/a_1141_508# prbs_generator_syn_27/sky130_fd_sc_hs__and2b_2_1/a_27_74#
+ prbs_generator_syn_27/sky130_fd_sc_hs__conb_1_1/a_165_290# prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_55/a_293_74#
+ prbs_generator_syn_27/sky130_fd_sc_hs__nand2_1_45/a_117_74# prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_63/a_112_119#
+ prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_49/a_222_392# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_37/a_1034_424#
+ prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_23/a_293_74# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_15/a_1141_508#
+ prbs_generator_syn_27/sky130_fd_sc_hs__nand2_1_5/a_117_74# prbs_generator_syn_27/m3_13600_13485#
+ prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_5/a_112_119# prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_13/a_376_368#
+ prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_51/a_376_368# prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_7/a_293_74#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_19/a_206_368# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_57/a_206_368#
+ prbs_generator_syn_27/sky130_fd_sc_hs__sdlclkp_2_1/a_318_74# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_29/a_437_503#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_49/a_651_503# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_25/a_27_74#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_5/a_1226_296# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_41/a_544_485#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_27/a_735_102# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_65/a_1141_508#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_65/a_735_102# prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_3/a_230_79#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_35/a_1034_424# prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_13/a_230_79#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_41/a_27_74# prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_3/a_132_392#
+ prbs_generator_syn_27/sky130_fd_sc_hs__nand2_1_49/a_117_74# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_27/a_1226_296#
+ prbs_generator_syn_27/sky130_fd_sc_hs__nand2_1_15/a_117_74# prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_41/a_376_368#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_45/a_1178_124# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_4/a_735_102#
+ prbs_generator_syn_27/sky130_fd_sc_hs__nand2_1_9/a_117_74# prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_33/a_138_385#
+ prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_17/a_132_392# prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_55/a_132_392#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_9/a_1141_508# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_19/a_437_503#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_57/a_437_503# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_4/a_1226_296#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_32/a_544_485# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_17/a_735_102#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_55/a_735_102# prbs_generator_syn_27/m3_13600_2261#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_65/a_27_74# prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_29/a_222_392#
+ prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_43/a_112_119# prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_19/X
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_25/a_1226_296# prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_31/a_376_368#
+ prbs_generator_syn_27/sky130_fd_sc_hs__or2_1_1/a_63_368# prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_17/a_230_79#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_4/a_27_74# prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_61/a_230_79#
+ prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_63/a_138_385# prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_5/a_222_392#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_8/a_1141_508# prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_41/a_293_74#
+ prbs_generator_syn_27/sky130_fd_sc_hs__nand2_1_31/a_117_74# prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_5/a_138_385#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_63/a_1141_508# prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_19/a_222_392#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_13/a_1141_508# prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_3/a_52_123#
+ prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_13/a_52_123# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_43/a_1178_124#
+ prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_61/a_376_368# prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_35/a_132_392#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_67/a_206_368# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_1/a_1226_296#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_69/a_696_458# prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_31/a_230_79#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_35/a_735_102# prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_23/a_112_119#
+ prbs_generator_syn_27/sky130_fd_sc_hs__nand2_1_35/a_117_74# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_59/a_27_74#
+ prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_13/a_293_74# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_5/a_206_368#
+ prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_50/a_376_368# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_7/a_696_458#
+ prbs_generator_syn_27/sky130_fd_sc_hs__nor2b_1_7/a_278_368# prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_17/a_52_123#
+ prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_43/a_138_385# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_7/a_1141_508#
+ prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_61/a_52_123# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_67/a_437_503#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_61/a_1141_508# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_25/a_735_102#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_59/a_696_458# prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_13/a_112_119#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_33/a_1034_424# prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_51/a_112_119#
+ prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_35/a_230_79# prbs_generator_syn_27/m3_13600_4091#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_23/a_1226_296# prbs_generator_syn_27/sky130_fd_sc_hs__nand2_1_39/a_117_74#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_29/a_27_74# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_5/a_437_503#
+ prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_17/a_293_74# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_41/a_1178_124#
+ prbs_generator_syn_27/sky130_fd_sc_hs__or2_1_1/a_152_368# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_59/a_1178_124#
+ prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_61/a_293_74# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_47/a_206_368#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_39/a_651_503# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_49/a_696_458#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_15/a_735_102# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_32/a_1034_424#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_73/a_1226_296# prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_27/a_222_392#
+ prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_41/a_112_119# prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_31/a_52_123#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_49/a_1034_424# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_29/a_1141_508#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_21/a_1226_296# prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_39/a_230_79#
+ prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_23/a_138_385# prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_51/a_230_79#
+ prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_45/a_132_392# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_37/a_206_368#
+ prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_65/a_293_74# prbs_generator_syn_27/sky130_fd_sc_hs__nand2_1_53/a_117_74#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_47/a_437_503# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_29/a_651_503#
+ prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_31/a_293_74# prbs_generator_syn_27/sky130_fd_sc_hs__nand2_1_21/a_117_74#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_69/a_544_485# prbs_generator_syn_27/sky130_fd_sc_hs__clkbuf_16_1/a_114_74#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_45/a_735_102# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_13/a_27_74#
+ prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_31/a_112_119# prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_57/a_222_392#
+ prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_35/a_52_123# prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_21/a_376_368#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_7/a_544_485# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_57/a_1178_124#
+ prbs_generator_syn_27/m3_13600_6043# prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_13/a_138_385#
+ prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_51/a_138_385# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_5/a_1141_508#
+ prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_3/a_376_368# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_27/a_206_368#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_65/a_206_368# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_37/a_437_503#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_19/a_651_503# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_57/a_651_503#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_59/a_544_485# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_71/a_1226_296#
+ prbs_generator_syn_27/sky130_fd_sc_hs__nand2_1_25/a_117_74# prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_61/a_112_119#
+ prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_47/a_222_392# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_27/a_1141_508#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_53/a_27_74# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_4/a_206_368#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_39/a_1226_296# prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_11/a_376_368#
+ prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_39/a_52_123# prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_41/a_138_385#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_4/a_1141_508# prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_25/a_132_392#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_17/a_206_368# prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_41/A
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_55/a_206_368# prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_51/a_52_123#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_27/a_437_503# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_65/a_437_503#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_49/a_544_485# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_63/a_735_102#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_47/a_1034_424# prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_50/a_112_119#
+ prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_37/a_222_392# prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_59/a_230_79#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_25/a_1141_508# prbs_generator_syn_27/sky130_fd_sc_hs__nor2b_1_4/a_27_112#
+ prbs_generator_syn_27/sky130_fd_sc_hs__sdlclkp_2_1/a_685_81# prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_1/a_132_392#
+ prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_39/a_293_74# prbs_generator_syn_27/sky130_fd_sc_hs__nand2_1_29/a_117_74#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_4/a_437_503# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_55/a_1178_124#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_21/a_27_74# prbs_generator_syn_27/m3_13600_12875#
+ prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_50/a_293_74# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_1/a_735_102#
+ prbs_generator_syn_27/sky130_fd_sc_hs__xnor2_1_31/a_138_385# prbs_generator_syn_27/sky130_fd_sc_hs__a22o_1_15/a_132_392#
+ prbs_generator_syn_27/sky130_fd_sc_hs__nand2_1_1/a_117_74# prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_17/a_437_503#
+ prbs_generator_syn_27/sky130_fd_sc_hs__dfxtp_4_55/a_437_503# prbs_generator_syn
Xsky130_fd_sc_hs__conb_1_7 DVSS: DVDD: DVDD: DVSS: prbs_generator_syn_3/eqn[9] sky130_fd_sc_hs__conb_1_7/HI
+ sky130_fd_sc_hs__conb_1_7/a_165_290# sky130_fd_sc_hs__conb_1_7/a_21_290# sky130_fd_sc_hs__conb_1
Xsky130_fd_sc_hs__buf_2_103 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__buf_2_103/A sky130_fd_sc_hs__buf_2_103/X
+ sky130_fd_sc_hs__buf_2_103/a_21_260# sky130_fd_sc_hs__buf_2
Xsky130_fd_sc_hs__buf_2_114 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__buf_2_115/A sky130_fd_sc_hs__buf_2_115/X
+ sky130_fd_sc_hs__buf_2_115/a_21_260# sky130_fd_sc_hs__buf_2
Xsky130_fd_sc_hs__buf_2_125 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__buf_2_125/A sky130_fd_sc_hs__buf_2_125/X
+ sky130_fd_sc_hs__buf_2_125/a_21_260# sky130_fd_sc_hs__buf_2
Xsky130_fd_sc_hs__buf_2_136 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__buf_2_137/A sky130_fd_sc_hs__buf_2_137/X
+ sky130_fd_sc_hs__buf_2_137/a_21_260# sky130_fd_sc_hs__buf_2
Xsky130_fd_sc_hs__buf_2_147 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__buf_2_147/A sky130_fd_sc_hs__buf_2_147/X
+ sky130_fd_sc_hs__buf_2_147/a_21_260# sky130_fd_sc_hs__buf_2
Xsky130_fd_sc_hs__buf_2_158 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__buf_2_159/A sky130_fd_sc_hs__buf_2_159/X
+ sky130_fd_sc_hs__buf_2_159/a_21_260# sky130_fd_sc_hs__buf_2
Xsky130_fd_sc_hs__einvp_2_15 DVSS: DVDD: DVDD: DVSS: dout_n sky130_fd_sc_hs__buf_8_1/A
+ sky130_fd_sc_hs__dlrtp_1_13/Q sky130_fd_sc_hs__einvp_2_15/a_263_323# sky130_fd_sc_hs__einvp_2_15/a_36_74#
+ sky130_fd_sc_hs__einvp_2_15/a_27_368# sky130_fd_sc_hs__einvp_2
Xsky130_fd_sc_hs__einvp_2_26 DVSS: DVDD: DVDD: DVSS: dout_n sky130_fd_sc_hs__einvp_2_9/A
+ sky130_fd_sc_hs__einvp_2_27/TE sky130_fd_sc_hs__einvp_2_27/a_263_323# sky130_fd_sc_hs__einvp_2_27/a_36_74#
+ sky130_fd_sc_hs__einvp_2_27/a_27_368# sky130_fd_sc_hs__einvp_2
Xsky130_fd_sc_hs__einvp_2_37 DVSS: DVDD: DVDD: DVSS: dout_n sky130_fd_sc_hs__buf_8_1/A
+ sky130_fd_sc_hs__dlrtp_1_24/Q sky130_fd_sc_hs__einvp_2_37/a_263_323# sky130_fd_sc_hs__einvp_2_37/a_36_74#
+ sky130_fd_sc_hs__einvp_2_37/a_27_368# sky130_fd_sc_hs__einvp_2
Xsky130_fd_sc_hs__einvp_2_48 DVSS: DVDD: DVDD: DVSS: dout_n sky130_fd_sc_hs__buf_8_1/A
+ sky130_fd_sc_hs__einvp_2_49/TE sky130_fd_sc_hs__einvp_2_49/a_263_323# sky130_fd_sc_hs__einvp_2_49/a_36_74#
+ sky130_fd_sc_hs__einvp_2_49/a_27_368# sky130_fd_sc_hs__einvp_2
Xsky130_fd_sc_hs__einvp_2_59 DVSS: DVDD: DVDD: DVSS: dout_p sky130_fd_sc_hs__einvp_2_99/A
+ sky130_fd_sc_hs__dlrtp_1_43/Q sky130_fd_sc_hs__einvp_2_59/a_263_323# sky130_fd_sc_hs__einvp_2_59/a_36_74#
+ sky130_fd_sc_hs__einvp_2_59/a_27_368# sky130_fd_sc_hs__einvp_2
Xsky130_fd_sc_hs__conb_1_14 DVSS: DVDD: DVDD: DVSS: prbs_generator_syn_9/eqn[16] sky130_fd_sc_hs__conb_1_15/HI
+ sky130_fd_sc_hs__conb_1_15/a_165_290# sky130_fd_sc_hs__conb_1_15/a_21_290# sky130_fd_sc_hs__conb_1
Xsky130_fd_sc_hs__conb_1_25 DVSS: DVDD: DVDD: DVSS: prbs_generator_syn_1/eqn[31] prbs_generator_syn_1/cke
+ sky130_fd_sc_hs__conb_1_25/a_165_290# sky130_fd_sc_hs__conb_1_25/a_21_290# sky130_fd_sc_hs__conb_1
Xsky130_fd_sc_hs__conb_1_36 DVSS: DVDD: DVDD: DVSS: prbs_generator_syn_3/eqn[28] sky130_fd_sc_hs__conb_1_37/HI
+ sky130_fd_sc_hs__conb_1_37/a_165_290# sky130_fd_sc_hs__conb_1_37/a_21_290# sky130_fd_sc_hs__conb_1
Xsky130_fd_sc_hs__conb_1_47 DVSS: DVDD: DVDD: DVSS: prbs_generator_syn_3/eqn[31] prbs_generator_syn_3/cke
+ sky130_fd_sc_hs__conb_1_47/a_165_290# sky130_fd_sc_hs__conb_1_47/a_21_290# sky130_fd_sc_hs__conb_1
Xsky130_fd_sc_hs__conb_1_58 DVSS: DVDD: DVDD: DVSS: prbs_generator_syn_11/eqn[9] sky130_fd_sc_hs__conb_1_59/HI
+ sky130_fd_sc_hs__conb_1_59/a_165_290# sky130_fd_sc_hs__conb_1_59/a_21_290# sky130_fd_sc_hs__conb_1
Xsky130_fd_sc_hs__inv_4_10 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__inv_4_11/Y sky130_fd_sc_hs__inv_4_11/A
+ sky130_fd_sc_hs__inv_4
Xsky130_fd_sc_hs__conb_1_69 DVSS: DVDD: DVDD: DVSS: prbs_generator_syn_7/eqn[28] sky130_fd_sc_hs__conb_1_69/HI
+ sky130_fd_sc_hs__conb_1_69/a_165_290# sky130_fd_sc_hs__conb_1_69/a_21_290# sky130_fd_sc_hs__conb_1
Xsky130_fd_sc_hs__inv_4_21 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__inv_4_21/Y sky130_fd_sc_hs__inv_4_21/A
+ sky130_fd_sc_hs__inv_4
Xsky130_fd_sc_hs__inv_4_32 DVSS: DVDD: DVDD: DVSS: osc_core_1/pi1_r[1] osc_core_1/pi1_l[1]
+ sky130_fd_sc_hs__inv_4
Xsky130_fd_sc_hs__inv_4_43 DVSS: DVDD: DVDD: DVSS: osc_core_1/pi2_r[1] osc_core_1/pi2_l[1]
+ sky130_fd_sc_hs__inv_4
Xsky130_fd_sc_hs__inv_4_54 DVSS: DVDD: DVDD: DVSS: osc_core_1/pi4_r[0] osc_core_1/pi4_l[0]
+ sky130_fd_sc_hs__inv_4
Xsky130_fd_sc_hs__inv_4_65 DVSS: DVDD: DVDD: DVSS: osc_core_1/pi3_r[1] osc_core_1/pi3_l[1]
+ sky130_fd_sc_hs__inv_4
Xsky130_fd_sc_hs__inv_4_76 DVSS: DVDD: DVDD: DVSS: hr_16t4_mux_top_3/din[10] prbs_generator_syn_19/out
+ sky130_fd_sc_hs__inv_4
Xsky130_fd_sc_hs__inv_4_87 DVSS: DVDD: DVDD: DVSS: hr_16t4_mux_top_3/din[2] hr_16t4_mux_top_1/din[2]
+ sky130_fd_sc_hs__inv_4
Xsky130_fd_sc_hs__dlrtp_1_16 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__dlrtp_1_17/Q
+ sky130_fd_sc_hs__dlrtp_1_9/GATE sky130_fd_sc_hs__conb_1_119/HI sky130_fd_sc_hs__dlrtp_1_17/D
+ sky130_fd_sc_hs__dlrtp_1_17/a_216_424# sky130_fd_sc_hs__dlrtp_1_17/a_759_508# sky130_fd_sc_hs__dlrtp_1_17/a_565_74#
+ sky130_fd_sc_hs__dlrtp_1_17/a_27_424# sky130_fd_sc_hs__dlrtp_1_17/a_1045_74# sky130_fd_sc_hs__dlrtp_1_17/a_643_74#
+ sky130_fd_sc_hs__dlrtp_1_17/a_817_48# sky130_fd_sc_hs__dlrtp_1_17/a_568_392# sky130_fd_sc_hs__dlrtp_1_17/a_363_74#
+ sky130_fd_sc_hs__dlrtp_1_17/a_769_74# sky130_fd_sc_hs__dlrtp_1
Xsky130_fd_sc_hs__dlrtp_1_27 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__dlrtp_1_27/Q
+ sky130_fd_sc_hs__clkbuf_2_3/A sky130_fd_sc_hs__conb_1_119/HI sky130_fd_sc_hs__dlrtp_1_27/D
+ sky130_fd_sc_hs__dlrtp_1_27/a_216_424# sky130_fd_sc_hs__dlrtp_1_27/a_759_508# sky130_fd_sc_hs__dlrtp_1_27/a_565_74#
+ sky130_fd_sc_hs__dlrtp_1_27/a_27_424# sky130_fd_sc_hs__dlrtp_1_27/a_1045_74# sky130_fd_sc_hs__dlrtp_1_27/a_643_74#
+ sky130_fd_sc_hs__dlrtp_1_27/a_817_48# sky130_fd_sc_hs__dlrtp_1_27/a_568_392# sky130_fd_sc_hs__dlrtp_1_27/a_363_74#
+ sky130_fd_sc_hs__dlrtp_1_27/a_769_74# sky130_fd_sc_hs__dlrtp_1
Xsky130_fd_sc_hs__dlrtp_1_38 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__dlrtp_1_39/Q
+ sky130_fd_sc_hs__clkbuf_16_53/A sky130_fd_sc_hs__conb_1_123/HI sky130_fd_sc_hs__buf_2_30/X
+ sky130_fd_sc_hs__dlrtp_1_39/a_216_424# sky130_fd_sc_hs__dlrtp_1_39/a_759_508# sky130_fd_sc_hs__dlrtp_1_39/a_565_74#
+ sky130_fd_sc_hs__dlrtp_1_39/a_27_424# sky130_fd_sc_hs__dlrtp_1_39/a_1045_74# sky130_fd_sc_hs__dlrtp_1_39/a_643_74#
+ sky130_fd_sc_hs__dlrtp_1_39/a_817_48# sky130_fd_sc_hs__dlrtp_1_39/a_568_392# sky130_fd_sc_hs__dlrtp_1_39/a_363_74#
+ sky130_fd_sc_hs__dlrtp_1_39/a_769_74# sky130_fd_sc_hs__dlrtp_1
Xsky130_fd_sc_hs__dlrtp_1_49 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__dlrtp_1_49/Q
+ sky130_fd_sc_hs__clkbuf_16_53/A sky130_fd_sc_hs__conb_1_123/HI sky130_fd_sc_hs__buf_2_29/X
+ sky130_fd_sc_hs__dlrtp_1_49/a_216_424# sky130_fd_sc_hs__dlrtp_1_49/a_759_508# sky130_fd_sc_hs__dlrtp_1_49/a_565_74#
+ sky130_fd_sc_hs__dlrtp_1_49/a_27_424# sky130_fd_sc_hs__dlrtp_1_49/a_1045_74# sky130_fd_sc_hs__dlrtp_1_49/a_643_74#
+ sky130_fd_sc_hs__dlrtp_1_49/a_817_48# sky130_fd_sc_hs__dlrtp_1_49/a_568_392# sky130_fd_sc_hs__dlrtp_1_49/a_363_74#
+ sky130_fd_sc_hs__dlrtp_1_49/a_769_74# sky130_fd_sc_hs__dlrtp_1
Xsky130_fd_sc_hs__einvp_2_9 DVSS: DVDD: DVDD: DVSS: dout_n sky130_fd_sc_hs__einvp_2_9/A
+ sky130_fd_sc_hs__dlrtp_1_9/Q sky130_fd_sc_hs__einvp_2_9/a_263_323# sky130_fd_sc_hs__einvp_2_9/a_36_74#
+ sky130_fd_sc_hs__einvp_2_9/a_27_368# sky130_fd_sc_hs__einvp_2
Xsky130_fd_sc_hs__clkbuf_16_70 DVSS: DVDD: DVDD: DVSS: prbs_generator_syn_13/rst prbs_generator_syn_19/rst
+ sky130_fd_sc_hs__clkbuf_16_71/a_114_74# sky130_fd_sc_hs__clkbuf_16
Xsky130_fd_sc_hs__clkbuf_16_81 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__or2b_2_1/A
+ sky130_fd_sc_hs__clkbuf_8_75/X sky130_fd_sc_hs__clkbuf_16_81/a_114_74# sky130_fd_sc_hs__clkbuf_16
Xsky130_fd_sc_hs__clkbuf_16_92 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__clkbuf_16_93/X
+ sky130_fd_sc_hs__clkbuf_4_115/X sky130_fd_sc_hs__clkbuf_16_93/a_114_74# sky130_fd_sc_hs__clkbuf_16
Xsky130_fd_sc_hs__clkbuf_8_100 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__clkinv_8_19/A
+ rst sky130_fd_sc_hs__clkbuf_8_101/a_125_368# sky130_fd_sc_hs__clkbuf_8
Xsky130_fd_sc_hs__buf_2_19 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__buf_2_33/A sky130_fd_sc_hs__buf_2_19/X
+ sky130_fd_sc_hs__buf_2_19/a_21_260# sky130_fd_sc_hs__buf_2
Xsky130_fd_sc_hs__nand2_2_11 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__inv_4_17/A sky130_fd_sc_hs__nand2_2_11/B
+ sky130_fd_sc_hs__inv_4_15/Y sky130_fd_sc_hs__nand2_2_11/a_27_74# sky130_fd_sc_hs__nand2_2
Xsky130_fd_sc_hs__nand2_2_22 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__nand2_2_23/Y
+ sky130_fd_sc_hs__nor4_2_1/C sky130_fd_sc_hs__nor4_2_1/B sky130_fd_sc_hs__nand2_2_23/a_27_74#
+ sky130_fd_sc_hs__nand2_2
Xsky130_fd_sc_hs__nand2_2_33 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__nand2_2_33/Y
+ sky130_fd_sc_hs__or4_2_1/B sky130_fd_sc_hs__or4_2_1/A sky130_fd_sc_hs__nand2_2_33/a_27_74#
+ sky130_fd_sc_hs__nand2_2
Xsky130_fd_sc_hs__conb_1_208 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__conb_1_209/LO
+ sky130_fd_sc_hs__conb_1_209/HI sky130_fd_sc_hs__conb_1_209/a_165_290# sky130_fd_sc_hs__conb_1_209/a_21_290#
+ sky130_fd_sc_hs__conb_1
Xsky130_fd_sc_hs__conb_1_219 DVSS: DVDD: DVDD: DVSS: prbs_generator_syn_25/eqn[30]
+ sky130_fd_sc_hs__conb_1_219/HI sky130_fd_sc_hs__conb_1_219/a_165_290# sky130_fd_sc_hs__conb_1_219/a_21_290#
+ sky130_fd_sc_hs__conb_1
Xprbs_generator_syn_0 prbs_generator_syn_9/clk prbs_generator_syn_9/rst prbs_generator_syn_1/cke
+ sky130_fd_sc_hs__conb_1_41/LO prbs_generator_syn_5/eqn[5] prbs_generator_syn_5/eqn[1]
+ prbs_generator_syn_5/eqn[1] prbs_generator_syn_5/eqn[1] prbs_generator_syn_5/eqn[1]
+ sky130_fd_sc_hs__conb_1_41/HI sky130_fd_sc_hs__conb_1_41/LO sky130_fd_sc_hs__conb_1_41/LO
+ sky130_fd_sc_hs__conb_1_41/LO sky130_fd_sc_hs__conb_1_41/LO prbs_generator_syn_1/eqn[31]
+ prbs_generator_syn_5/eqn[13] sky130_fd_sc_hs__conb_1_27/HI prbs_generator_syn_5/eqn[13]
+ sky130_fd_sc_hs__conb_1_27/HI prbs_generator_syn_5/eqn[13] sky130_fd_sc_hs__conb_1_27/HI
+ prbs_generator_syn_3/eqn[9] prbs_generator_syn_3/eqn[20] prbs_generator_syn_3/eqn[20]
+ prbs_generator_syn_3/eqn[20] prbs_generator_syn_3/eqn[20] prbs_generator_syn_3/eqn[28]
+ prbs_generator_syn_3/eqn[28] sky130_fd_sc_hs__conb_1_37/HI sky130_fd_sc_hs__conb_1_37/HI
+ prbs_generator_syn_3/eqn[30] sky130_fd_sc_hs__conb_1_45/HI prbs_generator_syn_3/eqn[30]
+ sky130_fd_sc_hs__conb_1_45/HI prbs_generator_syn_3/eqn[30] prbs_generator_syn_1/eqn[31]
+ prbs_generator_syn_1/eqn[30] prbs_generator_syn_1/eqn[30] prbs_generator_syn_1/eqn[30]
+ prbs_generator_syn_1/eqn[30] prbs_generator_syn_1/eqn[30] prbs_generator_syn_1/eqn[30]
+ prbs_generator_syn_1/eqn[30] prbs_generator_syn_1/eqn[30] sky130_fd_sc_hs__conb_1_3/LO
+ sky130_fd_sc_hs__conb_1_3/LO sky130_fd_sc_hs__conb_1_3/HI sky130_fd_sc_hs__conb_1_3/LO
+ sky130_fd_sc_hs__conb_1_3/LO sky130_fd_sc_hs__conb_1_3/LO sky130_fd_sc_hs__conb_1_3/LO
+ sky130_fd_sc_hs__conb_1_3/LO sky130_fd_sc_hs__conb_1_3/LO prbs_generator_syn_1/eqn[9]
+ prbs_generator_syn_1/eqn[9] prbs_generator_syn_1/eqn[9] prbs_generator_syn_1/eqn[9]
+ prbs_generator_syn_1/eqn[9] prbs_generator_syn_1/eqn[8] prbs_generator_syn_1/eqn[8]
+ prbs_generator_syn_1/eqn[8] prbs_generator_syn_1/eqn[8] prbs_generator_syn_1/eqn[8]
+ prbs_generator_syn_1/eqn[8] prbs_generator_syn_1/eqn[8] prbs_generator_syn_1/eqn[1]
+ prbs_generator_syn_3/eqn[9] prbs_generator_syn_9/inj_err prbs_generator_syn_1/eqn[31]
+ prbs_generator_syn_1/eqn[31] prbs_generator_syn_1/out DVSS: DVDD: prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_1/a_293_74#
+ prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_15/X prbs_generator_syn_1/sky130_fd_sc_hs__nand2_1_35/B
+ prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_51/Y prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_9/A
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_9/CLK prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_47/a_27_74#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_37/a_1226_296# prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_3/B
+ prbs_generator_syn_1/sky130_fd_sc_hs__nor2b_1_7/a_27_112# prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_29/B
+ prbs_generator_syn_1/sky130_fd_sc_hs__sdlclkp_2_1/a_580_74# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_1/a_1141_508#
+ prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_5/Y prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_41/a_230_79#
+ prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_61/a_138_385# prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_43/a_132_392#
+ prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_3/a_222_392# prbs_generator_syn_1/sky130_fd_sc_hs__nor2b_1_9/a_27_112#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_61/a_27_74# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_35/a_206_368#
+ prbs_generator_syn_1/sky130_fd_sc_hs__nand2_2_3/Y prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_25/B
+ prbs_generator_syn_1/sky130_fd_sc_hs__nand2_1_11/a_117_74# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_67/a_651_503#
+ prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_45/X prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_39/a_696_458#
+ prbs_generator_syn_1/sky130_fd_sc_hs__sdlclkp_2_1/a_1198_74# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_45/a_1034_424#
+ prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_17/a_222_392# prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_55/a_222_392#
+ prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_53/Y prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_35/A
+ prbs_generator_syn_1/m3_13600_1651# prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_59/a_52_123#
+ prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_5/a_293_74# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_35/a_1226_296#
+ prbs_generator_syn_1/sky130_fd_sc_hs__nand2_1_51/B prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_5/a_651_503#
+ prbs_generator_syn_1/sky130_fd_sc_hs__nand2_1_21/B prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_8/a_27_74#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_15/a_27_74# prbs_generator_syn_1/sky130_fd_sc_hs__and2b_2_1/X
+ prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_13/X prbs_generator_syn_1/sky130_fd_sc_hs__nand2_2_3/a_27_74#
+ prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_50/a_138_385# prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_33/a_132_392#
+ prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_1/a_376_368# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_25/a_206_368#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_35/a_437_503# prbs_generator_syn_1/sky130_fd_sc_hs__sdlclkp_2_1/a_708_451#
+ prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_45/a_230_79# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_29/a_696_458#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_32/a_27_74# prbs_generator_syn_1/sky130_fd_sc_hs__nor2b_1_4/Y
+ prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_59/a_293_74# prbs_generator_syn_1/sky130_fd_sc_hs__nand2_1_47/a_117_74#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_73/a_735_102# prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_21/a_112_119#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_23/a_1141_508# prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_25/a_293_74#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_7/Q prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_3/a_112_119#
+ prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_35/B prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_51/X
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_53/a_1178_124# prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_23/a_132_392#
+ prbs_generator_syn_1/sky130_fd_sc_hs__nand2_1_3/B prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_15/a_206_368#
+ prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_63/a_132_392# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_55/a_27_74#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_25/a_437_503# prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_41/a_52_123#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_47/a_651_503# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_73/a_1141_508#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_19/a_696_458# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_57/a_696_458#
+ prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_7/X prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_43/a_1034_424#
+ prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_55/A prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_11/a_112_119#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_21/a_1141_508# prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_35/a_222_392#
+ prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_49/a_230_79# prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_67/Y
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_71/a_27_74# prbs_generator_syn_1/sky130_fd_sc_hs__nand2_1_33/B
+ prbs_generator_syn_1/sky130_fd_sc_hs__conb_1_1/LO prbs_generator_syn_1/sky130_fd_sc_hs__nand2_1_19/a_117_74#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_51/a_1178_124# prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_33/X
+ prbs_generator_syn_1/sky130_fd_sc_hs__nand2_1_29/B prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_41/Y
+ prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_53/a_132_392# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_45/a_206_368#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_15/a_437_503# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_37/a_651_503#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_39/a_544_485# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_53/a_735_102#
+ prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_45/a_52_123# prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_1/B
+ prbs_generator_syn_1/sky130_fd_sc_hs__nand2_2_3/B prbs_generator_syn_1/sky130_fd_sc_hs__clkbuf_16_1/A
+ prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_21/X prbs_generator_syn_1/sky130_fd_sc_hs__nand2_1_25/B
+ prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_39/a_376_368# prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_63/X
+ prbs_generator_syn_1/m3_13600_3481# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_69/a_1178_124#
+ prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_21/a_138_385# prbs_generator_syn_1/sky130_fd_sc_hs__nor2b_1_8/Y
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_19/a_1178_124# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_49/a_27_74#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_45/a_437_503# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_27/a_651_503#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_71/a_1141_508# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_65/a_651_503#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_29/a_544_485# prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_3/a_138_385#
+ prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_55/X prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_43/a_735_102#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_41/a_1034_424# prbs_generator_syn_1/sky130_fd_sc_hs__nand2_1_9/B
+ prbs_generator_syn_1/sky130_fd_sc_hs__nor2b_1_9/Y prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_59/a_1034_424#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_39/a_1141_508# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_33/a_1226_296#
+ prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_49/a_52_123# prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_47/Y
+ prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_43/Y prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_4/a_651_503#
+ prbs_generator_syn_1/sky130_fd_sc_hs__nand2_1_49/B prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_19/A
+ prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_11/a_138_385# prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_5/X
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_63/a_206_368# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_17/a_651_503#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_19/a_544_485# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_55/a_651_503#
+ prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_9/Y prbs_generator_syn_1/sky130_fd_sc_hs__nand2_1_17/B
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_57/a_544_485# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_67/a_696_458#
+ prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_35/X prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_19/a_27_74#
+ prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_45/a_222_392# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_32/a_1226_296#
+ prbs_generator_syn_1/sky130_fd_sc_hs__nand2_1_43/B prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_25/A
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_1/a_206_368# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_49/a_1226_296#
+ prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_1/a_112_119# prbs_generator_syn_1/sky130_fd_sc_hs__or2_1_1/X
+ prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_59/a_376_368# prbs_generator_syn_1/sky130_fd_sc_hs__nand2_1_19/B
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_5/a_696_458# prbs_generator_syn_1/sky130_fd_sc_hs__nor2b_1_1/Y
+ prbs_generator_syn_1/sky130_fd_sc_hs__nor2b_1_5/a_278_368# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_17/a_1178_124#
+ prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_39/X prbs_generator_syn_1/m3_13600_5433#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_63/a_437_503# prbs_generator_syn_1/sky130_fd_sc_hs__nand2_2_5/B
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_23/a_735_102# prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_53/A
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_61/a_735_102# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_57/a_1034_424#
+ prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_63/B prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_37/a_1141_508#
+ prbs_generator_syn_1/sky130_fd_sc_hs__nand2_1_47/B prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_29/X
+ prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_65/Y prbs_generator_syn_1/m3_13600_4701#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_1/a_437_503# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_67/a_1178_124#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_9/a_735_102# prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_13/a_132_392#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_15/a_1178_124# prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_15/A
+ prbs_generator_syn_1/sky130_fd_sc_hs__nand2_1_1/B prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_43/B
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_35/a_651_503# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_8/D
+ prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_29/A prbs_generator_syn_1/sky130_fd_sc_hs__nand2_1_7/B
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_13/a_735_102# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_47/a_696_458#
+ prbs_generator_syn_1/sky130_fd_sc_hs__nand2_1_31/B prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_51/a_735_102#
+ prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_59/X prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_35/a_1141_508#
+ prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_25/a_222_392# prbs_generator_syn_1/sky130_fd_sc_hs__sdlclkp_2_1/a_288_48#
+ prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_55/B prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_17/B
+ prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_43/A prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_7/A
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_65/a_1178_124# prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_59/Y
+ prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_41/X prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_21/a_230_79#
+ prbs_generator_syn_1/sky130_fd_sc_hs__nand2_1_57/a_117_74# prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_1/a_222_392#
+ prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_19/B prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_35/a_293_74#
+ prbs_generator_syn_1/sky130_fd_sc_hs__nand2_1_23/a_117_74# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_73/a_206_368#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_25/a_651_503# prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_1/a_138_385#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_37/a_696_458# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_67/a_544_485#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_43/a_27_74# prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_9/X
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_55/a_1034_424# prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_39/a_112_119#
+ prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_15/a_222_392# prbs_generator_syn_1/sky130_fd_sc_hs__conb_1_1/HI
+ prbs_generator_syn_1/sky130_fd_sc_hs__nand2_1_23/B prbs_generator_syn_1/sky130_fd_sc_hs__nand2_1_53/B
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_9/a_1178_124# prbs_generator_syn_1/sky130_fd_sc_hs__nor2b_1_4/A
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_47/a_1226_296# prbs_generator_syn_1/m3_13600_11045#
+ prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_17/X prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_29/a_376_368#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_5/a_544_485# prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_3/X
+ prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_31/a_132_392# prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_61/A
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_15/a_651_503# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_73/a_437_503#
+ prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_25/a_230_79# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_27/a_696_458#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_65/a_696_458# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_33/a_735_102#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_71/a_735_102# prbs_generator_syn_1/m3_13600_7263#
+ prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_43/a_222_392# prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_50/Y
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_8/a_1178_124# prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_53/B
+ prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_19/a_376_368# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_63/a_1178_124#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_4/a_696_458# prbs_generator_syn_1/sky130_fd_sc_hs__nor2b_1_4/a_278_368#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_13/a_1178_124# prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_61/a_132_392#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_53/a_206_368# prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_21/a_52_123#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_45/a_651_503# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_17/a_696_458#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_47/a_544_485# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_55/a_696_458#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_21/a_735_102# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_37/a_27_74#
+ prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_61/B prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_61/X
+ prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_59/a_112_119# prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_31/A
+ prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_33/a_222_392# prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_29/a_230_79#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_45/a_1226_296# prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_9/a_132_392#
+ prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_5/A prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_57/Y
+ prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_31/X prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_51/a_27_74#
+ prbs_generator_syn_1/sky130_fd_sc_hs__nor2b_1_8/a_27_112# prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_47/a_376_368#
+ prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_53/a_293_74# prbs_generator_syn_1/sky130_fd_sc_hs__nand2_1_43/a_117_74#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_8/a_735_102# prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_21/a_293_74#
+ prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_39/a_138_385# prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_63/Y
+ prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_51/a_132_392# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_43/a_206_368#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_53/a_437_503# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_37/a_544_485#
+ prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_57/X prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_53/a_1034_424#
+ prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_25/a_52_123# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_33/a_1141_508#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_63/Q prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_23/a_222_392#
+ prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_63/a_222_392# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_7/a_1178_124#
+ prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_53/X prbs_generator_syn_1/sky130_fd_sc_hs__nand2_2_5/Y
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_61/a_1178_124# prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_1/a_230_79#
+ prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_43/a_230_79# prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_11/a_230_79#
+ prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_41/a_132_392# prbs_generator_syn_1/sky130_fd_sc_hs__nand2_1_13/a_117_74#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_43/a_437_503# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_27/a_544_485#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_63/a_651_503# prbs_generator_syn_1/sky130_fd_sc_hs__nand2_1_7/a_117_74#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_35/a_696_458# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_65/a_544_485#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_51/a_1034_424# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_41/a_735_102#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_32/a_1141_508# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_49/a_1141_508#
+ prbs_generator_syn_1/sky130_fd_sc_hs__nand2_1_55/B prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_53/a_222_392#
+ prbs_generator_syn_1/sky130_fd_sc_hs__sdlclkp_2_1/a_114_112# prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_9/a_293_74#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_43/a_1226_296# prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_29/a_52_123#
+ prbs_generator_syn_1/sky130_fd_sc_hs__nand2_1_37/B prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_1/a_651_503#
+ prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_27/a_376_368# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_4/a_544_485#
+ prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_67/a_376_368# prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_27/X
+ prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_1/X prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_59/a_138_385#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_29/a_1178_124# prbs_generator_syn_1/m3_13600_2871#
+ prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_5/a_230_79# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_23/a_206_368#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_61/a_206_368# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_17/a_544_485#
+ prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_15/a_230_79# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_25/a_696_458#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_55/a_544_485# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_32/a_735_102#
+ prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_29/a_293_74# prbs_generator_syn_1/sky130_fd_sc_hs__nand2_1_17/a_117_74#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_69/a_1034_424# prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_29/a_112_119#
+ prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_37/X prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_31/B
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_19/a_1034_424# prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_33/A
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_9/a_206_368# prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_57/a_376_368#
+ prbs_generator_syn_1/sky130_fd_sc_hs__sdlclkp_2_1/a_706_317# prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_11/B
+ prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_1/a_52_123# prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_39/B
+ prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_21/a_132_392# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_13/a_206_368#
+ prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_43/a_52_123# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_51/a_206_368#
+ prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_47/X prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_23/a_437_503#
+ prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_11/a_52_123# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_61/a_437_503#
+ prbs_generator_syn_1/sky130_fd_sc_hs__nor2b_1_7/Y prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_51/A
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_15/a_696_458# prbs_generator_syn_1/sky130_fd_sc_hs__nor2b_1_5/Y
+ prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_9/a_230_79# prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_25/X
+ prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_19/a_112_119# prbs_generator_syn_1/sky130_fd_sc_hs__nand2_1_45/B
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_5/a_1178_124# prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_19/a_230_79#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_41/a_1226_296# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_59/a_1226_296#
+ prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_63/a_230_79# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_51/Q
+ prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_7/a_132_392# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_9/a_437_503#
+ prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_46/a_376_368# prbs_generator_syn_1/sky130_fd_sc_hs__nand2_1_33/a_117_74#
+ prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_11/a_293_74# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_27/a_1178_124#
+ prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_11/a_132_392# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_13/a_437_503#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_51/a_437_503# prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_5/a_52_123#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_35/a_544_485# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_73/a_651_503#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_45/a_696_458# prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_15/a_52_123#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_47/a_1141_508# prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_47/a_112_119#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_4/a_1178_124# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_17/a_1034_424#
+ prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_23/B prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_37/a_376_368#
+ prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_15/B prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_7/Y
+ prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_29/a_138_385# prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_33/a_230_79#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_25/a_1178_124# prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_47/a_293_74#
+ prbs_generator_syn_1/sky130_fd_sc_hs__nand2_1_37/a_117_74# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_33/a_206_368#
+ prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_15/a_293_74# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_71/a_206_368#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_25/a_544_485# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_67/a_1034_424#
+ prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_13/a_222_392# prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_9/a_52_123#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_15/a_1034_424# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_57/a_1226_296#
+ prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_19/a_52_123# prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_23/X
+ prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_63/a_52_123# prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_19/a_138_385#
+ prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_9/a_376_368# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_21/a_206_368#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_33/a_437_503# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_71/a_437_503#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_53/a_651_503# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_15/a_544_485#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_63/a_696_458# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_65/a_1034_424#
+ prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_19/a_293_74# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_45/a_1141_508#
+ prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_27/a_112_119# prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_67/a_112_119#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_1/a_1178_124# prbs_generator_syn_1/sky130_fd_sc_hs__conb_1_1/a_21_290#
+ prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_63/a_293_74# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_8/a_206_368#
+ prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_17/a_376_368# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_63/a_27_74#
+ prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_21/A prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_55/a_376_368#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_1/a_696_458# prbs_generator_syn_1/sky130_fd_sc_hs__nor2b_1_1/a_278_368#
+ prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_47/a_138_385# prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_33/a_52_123#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_9/a_1034_424# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_21/a_437_503#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_1/a_27_74# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_43/a_651_503#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_1/Q prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_45/a_544_485#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_69/a_735_102# prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_57/a_112_119#
+ prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_31/a_222_392# prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_13/A
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_55/a_1226_296# prbs_generator_syn_1/sky130_fd_sc_hs__nand2_2_5/a_27_74#
+ prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_53/a_230_79# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_8/a_437_503#
+ prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_67/a_293_74# prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_33/a_293_74#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_7/a_735_102# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_23/a_1178_124#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_41/a_206_368# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_8/a_1034_424#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_63/a_1034_424# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_59/a_735_102#
+ prbs_generator_syn_1/sky130_fd_sc_hs__nand2_1_5/B prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_43/a_1141_508#
+ prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_46/a_112_119# prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_61/a_222_392#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_13/a_1034_424# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_73/a_1178_124#
+ prbs_generator_syn_1/sky130_fd_sc_hs__nand2_1_27/B prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_13/B
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_57/a_27_74# prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_57/a_230_79#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_21/a_1178_124# prbs_generator_syn_1/sky130_fd_sc_hs__nor2b_1_1/a_27_112#
+ prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_27/a_138_385# prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_23/a_230_79#
+ prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_67/a_138_385# prbs_generator_syn_1/sky130_fd_sc_hs__nand2_1_41/B
+ prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_9/a_222_392# prbs_generator_syn_1/sky130_fd_sc_hs__nand2_1_27/a_117_74#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_32/a_206_368# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_23/a_651_503#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_41/a_437_503# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_73/a_27_74#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_61/a_651_503# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_63/a_544_485#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_49/a_735_102# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_73/a_696_458#
+ prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_37/a_112_119# prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_51/a_222_392#
+ prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_43/X prbs_generator_syn_1/sky130_fd_sc_hs__nand2_2_1/B
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_9/a_651_503# prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_53/a_52_123#
+ prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_49/X prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_25/a_376_368#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_1/a_544_485# prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_65/a_376_368#
+ prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_57/a_138_385# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_27/a_27_74#
+ prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_39/a_132_392# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_7/a_1034_424#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_13/a_651_503# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_32/a_437_503#
+ prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_27/a_230_79# prbs_generator_syn_1/m3_13600_12265#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_51/a_651_503# prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_59/B
+ prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_47/A prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_61/a_1034_424#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_41/a_1141_508# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_59/a_1141_508#
+ prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_41/a_222_392# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_53/a_1226_296#
+ prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_3/A prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_71/a_1178_124#
+ prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_9/a_112_119# prbs_generator_syn_1/sky130_fd_sc_hs__nand2_1_3/a_117_74#
+ prbs_generator_syn_1/m3_13600_8483# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_39/a_1178_124#
+ prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_57/a_52_123# prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_46/a_138_385#
+ prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_23/a_52_123# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_67/a_27_74#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_53/a_696_458# prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_17/a_112_119#
+ prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_11/A prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_55/a_112_119#
+ prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_1/A prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_51/a_1226_296#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_29/a_1034_424# prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_59/A
+ prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_23/A prbs_generator_syn_1/sky130_fd_sc_hs__nand2_1_39/B
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_5/a_27_74# prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_57/a_293_74#
+ prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_37/a_138_385# prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_59/a_132_392#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_33/a_651_503# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_71/a_651_503#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_43/a_696_458# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_73/a_544_485#
+ prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_27/a_52_123# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_57/a_1141_508#
+ prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_21/a_222_392# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_35/a_27_74#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_69/a_1226_296# prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_37/B
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_19/a_1226_296# prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_35/a_376_368#
+ prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_47/a_230_79# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_37/a_1178_124#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_5/a_1034_424# prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_49/a_132_392#
+ prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_7/a_222_392# prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_27/a_293_74#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_21/a_651_503# prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_9/a_138_385#
+ prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_11/a_222_392# prbs_generator_syn_1/m3_13600_14095#
+ prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_50/A prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_27/a_1034_424#
+ prbs_generator_syn_1/sky130_fd_sc_hs__nand2_1_13/B prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_8/a_651_503#
+ prbs_generator_syn_1/m3_13600_9703# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_35/a_1178_124#
+ prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_17/a_138_385# prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_55/a_138_385#
+ prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_7/a_230_79# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_4/a_1034_424#
+ prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_7/a_376_368# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_69/a_206_368#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_23/a_696_458# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_53/a_544_485#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_39/a_735_102# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_61/a_696_458#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_55/a_1141_508# prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_25/a_112_119#
+ prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_65/a_112_119# prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_43/a_293_74#
+ prbs_generator_syn_1/sky130_fd_sc_hs__nand2_1_57/B prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_25/a_1034_424#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_7/a_206_368# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_17/a_1226_296#
+ prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_15/a_376_368# prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_53/a_376_368#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_9/a_696_458# prbs_generator_syn_1/m3_13600_431#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_45/a_27_74# prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_47/a_52_123#
+ prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_29/a_132_392# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_59/a_206_368#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_69/a_437_503# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_41/a_651_503#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_43/a_544_485# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_13/a_696_458#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_29/a_735_102# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_51/a_696_458#
+ prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_61/Y prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_67/a_1226_296#
+ prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_5/a_132_392# prbs_generator_syn_1/sky130_fd_sc_hs__and2b_2_1/a_198_48#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_7/a_437_503# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_15/a_1226_296#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_69/a_27_74# prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_46/a_293_74#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_1/a_1034_424# prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_19/a_132_392#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_49/a_206_368# prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_7/a_52_123#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_59/a_437_503# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_32/a_651_503#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_7/a_27_74# prbs_generator_syn_1/sky130_fd_sc_hs__nand2_2_1/a_27_74#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_19/a_735_102# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_57/a_735_102#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_65/a_1226_296# prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_37/A
+ prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_33/a_376_368# prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_37/a_230_79#
+ prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_25/a_138_385# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_39/a_27_74#
+ prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_65/a_138_385# prbs_generator_syn_1/sky130_fd_sc_hs__nor2b_1_9/a_278_368#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_49/a_437_503# prbs_generator_syn_1/sky130_fd_sc_hs__and2b_2_1/a_505_74#
+ prbs_generator_syn_1/sky130_fd_sc_hs__nand2_1_51/a_117_74# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_23/a_544_485#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_33/a_696_458# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_61/a_544_485#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_9/a_1226_296# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_53/a_1141_508#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_71/a_696_458# prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_35/a_112_119#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_23/a_1034_424# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_9/a_544_485#
+ prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_63/a_376_368# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_33/a_1178_124#
+ prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_5/a_376_368# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_13/a_544_485#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_73/a_1034_424# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_21/a_696_458#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_51/a_544_485# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_8/a_1226_296#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_51/a_1141_508# prbs_generator_syn_1/sky130_fd_sc_hs__nand2_1_55/a_117_74#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_21/a_1034_424# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_63/a_1226_296#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_23/a_27_74# prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_7/a_112_119#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_13/a_1226_296# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_8/a_696_458#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_32/a_1178_124# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_49/a_1178_124#
+ prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_37/a_52_123# prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_27/a_132_392#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_71/Q prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_67/a_735_102#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_69/a_1141_508# prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_15/a_112_119#
+ prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_53/a_112_119# prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_39/a_222_392#
+ prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_55/a_230_79# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_19/a_1141_508#
+ prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_37/a_293_74# prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_43/a_376_368#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_5/a_735_102# prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_35/a_138_385#
+ prbs_generator_syn_1/sky130_fd_sc_hs__sdlclkp_2_1/a_114_424# prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_57/a_132_392#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_71/a_1034_424# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_7/a_1226_296#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_33/a_544_485# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_41/a_696_458#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_71/a_544_485# prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_21/B
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_61/a_1226_296# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_39/a_1034_424#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_17/a_27_74# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_9/a_27_74#
+ prbs_generator_syn_1/sky130_fd_sc_hs__nor2b_1_5/a_27_112# prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_47/a_132_392#
+ prbs_generator_syn_1/sky130_fd_sc_hs__nor2b_1_8/a_278_368# prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_9/B
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_39/a_206_368# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_33/a_27_74#
+ prbs_generator_syn_1/sky130_fd_sc_hs__nand2_1_41/a_117_74# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_69/a_651_503#
+ prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_51/a_293_74# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_21/a_544_485#
+ prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_7/a_138_385# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_32/a_696_458#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_47/a_735_102# prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_33/a_112_119#
+ prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_59/a_222_392# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_17/a_1141_508#
+ prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_55/a_52_123# prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_3/a_293_74#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_7/a_651_503# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_29/a_1226_296#
+ prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_23/a_376_368# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_8/a_544_485#
+ prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_47/B prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_47/a_1178_124#
+ prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_15/a_138_385# prbs_generator_syn_1/sky130_fd_sc_hs__sdlclkp_2_1/a_1195_374#
+ prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_53/a_138_385# prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_37/a_132_392#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_29/a_206_368# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_39/a_437_503#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_59/a_651_503# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_37/a_735_102#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_67/a_1141_508# prbs_generator_syn_1/sky130_fd_sc_hs__and2b_2_1/a_27_74#
+ prbs_generator_syn_1/sky130_fd_sc_hs__conb_1_1/a_165_290# prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_55/a_293_74#
+ prbs_generator_syn_1/sky130_fd_sc_hs__nand2_1_45/a_117_74# prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_63/a_112_119#
+ prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_49/a_222_392# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_37/a_1034_424#
+ prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_23/a_293_74# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_15/a_1141_508#
+ prbs_generator_syn_1/sky130_fd_sc_hs__nand2_1_5/a_117_74# prbs_generator_syn_1/m3_13600_13485#
+ prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_5/a_112_119# prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_13/a_376_368#
+ prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_51/a_376_368# prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_7/a_293_74#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_19/a_206_368# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_57/a_206_368#
+ prbs_generator_syn_1/sky130_fd_sc_hs__sdlclkp_2_1/a_318_74# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_29/a_437_503#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_49/a_651_503# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_25/a_27_74#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_5/a_1226_296# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_41/a_544_485#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_27/a_735_102# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_65/a_1141_508#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_65/a_735_102# prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_3/a_230_79#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_35/a_1034_424# prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_13/a_230_79#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_41/a_27_74# prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_3/a_132_392#
+ prbs_generator_syn_1/sky130_fd_sc_hs__nand2_1_49/a_117_74# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_27/a_1226_296#
+ prbs_generator_syn_1/sky130_fd_sc_hs__nand2_1_15/a_117_74# prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_41/a_376_368#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_45/a_1178_124# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_4/a_735_102#
+ prbs_generator_syn_1/sky130_fd_sc_hs__nand2_1_9/a_117_74# prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_33/a_138_385#
+ prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_17/a_132_392# prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_55/a_132_392#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_9/a_1141_508# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_19/a_437_503#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_57/a_437_503# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_4/a_1226_296#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_32/a_544_485# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_17/a_735_102#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_55/a_735_102# prbs_generator_syn_1/m3_13600_2261#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_65/a_27_74# prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_29/a_222_392#
+ prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_43/a_112_119# prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_19/X
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_25/a_1226_296# prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_31/a_376_368#
+ prbs_generator_syn_1/sky130_fd_sc_hs__or2_1_1/a_63_368# prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_17/a_230_79#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_4/a_27_74# prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_61/a_230_79#
+ prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_63/a_138_385# prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_5/a_222_392#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_8/a_1141_508# prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_41/a_293_74#
+ prbs_generator_syn_1/sky130_fd_sc_hs__nand2_1_31/a_117_74# prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_5/a_138_385#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_63/a_1141_508# prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_19/a_222_392#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_13/a_1141_508# prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_3/a_52_123#
+ prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_13/a_52_123# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_43/a_1178_124#
+ prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_61/a_376_368# prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_35/a_132_392#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_67/a_206_368# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_1/a_1226_296#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_69/a_696_458# prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_31/a_230_79#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_35/a_735_102# prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_23/a_112_119#
+ prbs_generator_syn_1/sky130_fd_sc_hs__nand2_1_35/a_117_74# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_59/a_27_74#
+ prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_13/a_293_74# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_5/a_206_368#
+ prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_50/a_376_368# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_7/a_696_458#
+ prbs_generator_syn_1/sky130_fd_sc_hs__nor2b_1_7/a_278_368# prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_17/a_52_123#
+ prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_43/a_138_385# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_7/a_1141_508#
+ prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_61/a_52_123# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_67/a_437_503#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_61/a_1141_508# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_25/a_735_102#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_59/a_696_458# prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_13/a_112_119#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_33/a_1034_424# prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_51/a_112_119#
+ prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_35/a_230_79# prbs_generator_syn_1/m3_13600_4091#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_23/a_1226_296# prbs_generator_syn_1/sky130_fd_sc_hs__nand2_1_39/a_117_74#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_29/a_27_74# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_5/a_437_503#
+ prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_17/a_293_74# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_41/a_1178_124#
+ prbs_generator_syn_1/sky130_fd_sc_hs__or2_1_1/a_152_368# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_59/a_1178_124#
+ prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_61/a_293_74# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_47/a_206_368#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_39/a_651_503# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_49/a_696_458#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_15/a_735_102# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_32/a_1034_424#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_73/a_1226_296# prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_27/a_222_392#
+ prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_41/a_112_119# prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_31/a_52_123#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_49/a_1034_424# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_29/a_1141_508#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_21/a_1226_296# prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_39/a_230_79#
+ prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_23/a_138_385# prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_51/a_230_79#
+ prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_45/a_132_392# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_37/a_206_368#
+ prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_65/a_293_74# prbs_generator_syn_1/sky130_fd_sc_hs__nand2_1_53/a_117_74#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_47/a_437_503# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_29/a_651_503#
+ prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_31/a_293_74# prbs_generator_syn_1/sky130_fd_sc_hs__nand2_1_21/a_117_74#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_69/a_544_485# prbs_generator_syn_1/sky130_fd_sc_hs__clkbuf_16_1/a_114_74#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_45/a_735_102# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_13/a_27_74#
+ prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_31/a_112_119# prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_57/a_222_392#
+ prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_35/a_52_123# prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_21/a_376_368#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_7/a_544_485# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_57/a_1178_124#
+ prbs_generator_syn_1/m3_13600_6043# prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_13/a_138_385#
+ prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_51/a_138_385# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_5/a_1141_508#
+ prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_3/a_376_368# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_27/a_206_368#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_65/a_206_368# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_37/a_437_503#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_19/a_651_503# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_57/a_651_503#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_59/a_544_485# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_71/a_1226_296#
+ prbs_generator_syn_1/sky130_fd_sc_hs__nand2_1_25/a_117_74# prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_61/a_112_119#
+ prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_47/a_222_392# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_27/a_1141_508#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_53/a_27_74# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_4/a_206_368#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_39/a_1226_296# prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_11/a_376_368#
+ prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_39/a_52_123# prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_41/a_138_385#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_4/a_1141_508# prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_25/a_132_392#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_17/a_206_368# prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_41/A
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_55/a_206_368# prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_51/a_52_123#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_27/a_437_503# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_65/a_437_503#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_49/a_544_485# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_63/a_735_102#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_47/a_1034_424# prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_50/a_112_119#
+ prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_37/a_222_392# prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_59/a_230_79#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_25/a_1141_508# prbs_generator_syn_1/sky130_fd_sc_hs__nor2b_1_4/a_27_112#
+ prbs_generator_syn_1/sky130_fd_sc_hs__sdlclkp_2_1/a_685_81# prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_1/a_132_392#
+ prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_39/a_293_74# prbs_generator_syn_1/sky130_fd_sc_hs__nand2_1_29/a_117_74#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_4/a_437_503# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_55/a_1178_124#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_21/a_27_74# prbs_generator_syn_1/m3_13600_12875#
+ prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_50/a_293_74# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_1/a_735_102#
+ prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_31/a_138_385# prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_15/a_132_392#
+ prbs_generator_syn_1/sky130_fd_sc_hs__nand2_1_1/a_117_74# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_17/a_437_503#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_55/a_437_503# prbs_generator_syn
Xsky130_fd_sc_hs__o21bai_2_7 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__nand2_2_7/A
+ sky130_fd_sc_hs__inv_8_1/Y sky130_fd_sc_hs__dlrtp_1_71/D sky130_fd_sc_hs__buf_2_59/A
+ sky130_fd_sc_hs__o21bai_2_7/a_27_74# sky130_fd_sc_hs__o21bai_2_7/a_225_74# sky130_fd_sc_hs__o21bai_2_7/a_507_368#
+ sky130_fd_sc_hs__o21bai_2
Xsky130_fd_sc_hs__o21ai_2_12 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__inv_4_13/Y sky130_fd_sc_hs__nand2_2_9/B
+ sky130_fd_sc_hs__o21ai_2_55/A1 sky130_fd_sc_hs__buf_2_47/A sky130_fd_sc_hs__o21ai_2_13/a_116_368#
+ sky130_fd_sc_hs__o21ai_2_13/a_27_74# sky130_fd_sc_hs__o21ai_2
Xsky130_fd_sc_hs__o21ai_2_23 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__inv_4_15/Y sky130_fd_sc_hs__o21ai_2_23/A2
+ sky130_fd_sc_hs__buf_2_77/X sky130_fd_sc_hs__o21ai_2_23/Y sky130_fd_sc_hs__o21ai_2_23/a_116_368#
+ sky130_fd_sc_hs__o21ai_2_23/a_27_74# sky130_fd_sc_hs__o21ai_2
Xsky130_fd_sc_hs__o21ai_2_34 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__inv_4_21/Y sky130_fd_sc_hs__buf_8_3/X
+ sky130_fd_sc_hs__clkinv_4_7/Y sky130_fd_sc_hs__buf_2_91/A sky130_fd_sc_hs__o21ai_2_35/a_116_368#
+ sky130_fd_sc_hs__o21ai_2_35/a_27_74# sky130_fd_sc_hs__o21ai_2
Xsky130_fd_sc_hs__o21ai_2_45 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__nand2_2_27/B
+ sky130_fd_sc_hs__nand2_2_21/B sky130_fd_sc_hs__or2b_4_1/A sky130_fd_sc_hs__o21ai_2_45/Y
+ sky130_fd_sc_hs__o21ai_2_45/a_116_368# sky130_fd_sc_hs__o21ai_2_45/a_27_74# sky130_fd_sc_hs__o21ai_2
Xsky130_fd_sc_hs__o21ai_2_56 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__inv_4_29/A sky130_fd_sc_hs__o21ai_2_3/A2
+ sky130_fd_sc_hs__or2b_4_3/X sky130_fd_sc_hs__buf_2_157/A sky130_fd_sc_hs__o21ai_2_57/a_116_368#
+ sky130_fd_sc_hs__o21ai_2_57/a_27_74# sky130_fd_sc_hs__o21ai_2
Xsky130_fd_sc_hs__clkinv_4_15 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__o21ai_2_55/A1
+ sky130_fd_sc_hs__or4_2_1/B sky130_fd_sc_hs__clkinv_4
Xprbs_generator_syn_17 prbs_generator_syn_19/clk prbs_generator_syn_19/rst prbs_generator_syn_17/cke
+ sky130_fd_sc_hs__conb_1_161/LO sky130_fd_sc_hs__conb_1_161/LO sky130_fd_sc_hs__conb_1_161/LO
+ sky130_fd_sc_hs__conb_1_161/HI sky130_fd_sc_hs__conb_1_161/HI sky130_fd_sc_hs__conb_1_161/HI
+ sky130_fd_sc_hs__conb_1_161/HI sky130_fd_sc_hs__conb_1_161/HI sky130_fd_sc_hs__conb_1_161/LO
+ sky130_fd_sc_hs__conb_1_161/LO sky130_fd_sc_hs__conb_1_161/LO prbs_generator_syn_17/eqn[31]
+ prbs_generator_syn_19/eqn[13] prbs_generator_syn_19/eqn[13] sky130_fd_sc_hs__conb_1_193/HI
+ prbs_generator_syn_19/eqn[13] sky130_fd_sc_hs__conb_1_193/HI prbs_generator_syn_19/eqn[13]
+ prbs_generator_syn_17/eqn[1] prbs_generator_syn_17/eqn[2] prbs_generator_syn_17/eqn[1]
+ prbs_generator_syn_17/eqn[2] prbs_generator_syn_17/eqn[1] prbs_generator_syn_17/eqn[2]
+ sky130_fd_sc_hs__conb_1_165/LO sky130_fd_sc_hs__conb_1_165/HI sky130_fd_sc_hs__conb_1_165/HI
+ sky130_fd_sc_hs__conb_1_165/LO sky130_fd_sc_hs__conb_1_165/LO sky130_fd_sc_hs__conb_1_165/LO
+ sky130_fd_sc_hs__conb_1_165/LO sky130_fd_sc_hs__conb_1_165/LO prbs_generator_syn_17/eqn[31]
+ prbs_generator_syn_17/eqn[30] prbs_generator_syn_17/eqn[30] prbs_generator_syn_17/eqn[30]
+ prbs_generator_syn_17/eqn[30] prbs_generator_syn_17/eqn[30] prbs_generator_syn_17/eqn[30]
+ prbs_generator_syn_17/eqn[30] prbs_generator_syn_17/eqn[30] prbs_generator_syn_17/eqn[22]
+ prbs_generator_syn_17/eqn[22] prbs_generator_syn_17/eqn[20] prbs_generator_syn_17/eqn[22]
+ prbs_generator_syn_17/eqn[22] prbs_generator_syn_17/eqn[22] prbs_generator_syn_17/eqn[22]
+ prbs_generator_syn_17/eqn[22] prbs_generator_syn_17/eqn[22] prbs_generator_syn_17/eqn[13]
+ prbs_generator_syn_17/eqn[13] prbs_generator_syn_17/eqn[13] prbs_generator_syn_17/eqn[9]
+ prbs_generator_syn_17/eqn[9] prbs_generator_syn_17/eqn[9] prbs_generator_syn_17/eqn[9]
+ prbs_generator_syn_17/eqn[9] prbs_generator_syn_17/eqn[9] prbs_generator_syn_17/eqn[9]
+ prbs_generator_syn_17/eqn[9] prbs_generator_syn_17/eqn[2] prbs_generator_syn_17/eqn[1]
+ prbs_generator_syn_17/eqn[2] prbs_generator_syn_19/inj_err prbs_generator_syn_17/eqn[31]
+ prbs_generator_syn_17/eqn[31] prbs_generator_syn_17/out DVSS: DVDD: prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_1/a_293_74#
+ prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_15/X prbs_generator_syn_17/sky130_fd_sc_hs__nand2_1_35/B
+ prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_51/Y prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_9/A
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_9/CLK prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_47/a_27_74#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_37/a_1226_296# prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_3/B
+ prbs_generator_syn_17/sky130_fd_sc_hs__nor2b_1_7/a_27_112# prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_29/B
+ prbs_generator_syn_17/sky130_fd_sc_hs__sdlclkp_2_1/a_580_74# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_1/a_1141_508#
+ prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_5/Y prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_41/a_230_79#
+ prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_61/a_138_385# prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_43/a_132_392#
+ prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_3/a_222_392# prbs_generator_syn_17/sky130_fd_sc_hs__nor2b_1_9/a_27_112#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_61/a_27_74# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_35/a_206_368#
+ prbs_generator_syn_17/sky130_fd_sc_hs__nand2_2_3/Y prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_25/B
+ prbs_generator_syn_17/sky130_fd_sc_hs__nand2_1_11/a_117_74# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_67/a_651_503#
+ prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_45/X prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_39/a_696_458#
+ prbs_generator_syn_17/sky130_fd_sc_hs__sdlclkp_2_1/a_1198_74# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_45/a_1034_424#
+ prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_17/a_222_392# prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_55/a_222_392#
+ prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_53/Y prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_35/A
+ prbs_generator_syn_17/m3_13600_1651# prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_59/a_52_123#
+ prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_5/a_293_74# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_35/a_1226_296#
+ prbs_generator_syn_17/sky130_fd_sc_hs__nand2_1_51/B prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_5/a_651_503#
+ prbs_generator_syn_17/sky130_fd_sc_hs__nand2_1_21/B prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_8/a_27_74#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_15/a_27_74# prbs_generator_syn_17/sky130_fd_sc_hs__and2b_2_1/X
+ prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_13/X prbs_generator_syn_17/sky130_fd_sc_hs__nand2_2_3/a_27_74#
+ prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_50/a_138_385# prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_33/a_132_392#
+ prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_1/a_376_368# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_25/a_206_368#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_35/a_437_503# prbs_generator_syn_17/sky130_fd_sc_hs__sdlclkp_2_1/a_708_451#
+ prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_45/a_230_79# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_29/a_696_458#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_32/a_27_74# prbs_generator_syn_17/sky130_fd_sc_hs__nor2b_1_4/Y
+ prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_59/a_293_74# prbs_generator_syn_17/sky130_fd_sc_hs__nand2_1_47/a_117_74#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_73/a_735_102# prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_21/a_112_119#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_23/a_1141_508# prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_25/a_293_74#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_7/Q prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_3/a_112_119#
+ prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_35/B prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_51/X
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_53/a_1178_124# prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_23/a_132_392#
+ prbs_generator_syn_17/sky130_fd_sc_hs__nand2_1_3/B prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_15/a_206_368#
+ prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_63/a_132_392# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_55/a_27_74#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_25/a_437_503# prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_41/a_52_123#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_47/a_651_503# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_73/a_1141_508#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_19/a_696_458# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_57/a_696_458#
+ prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_7/X prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_43/a_1034_424#
+ prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_55/A prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_11/a_112_119#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_21/a_1141_508# prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_35/a_222_392#
+ prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_49/a_230_79# prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_67/Y
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_71/a_27_74# prbs_generator_syn_17/sky130_fd_sc_hs__nand2_1_33/B
+ prbs_generator_syn_17/sky130_fd_sc_hs__conb_1_1/LO prbs_generator_syn_17/sky130_fd_sc_hs__nand2_1_19/a_117_74#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_51/a_1178_124# prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_33/X
+ prbs_generator_syn_17/sky130_fd_sc_hs__nand2_1_29/B prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_41/Y
+ prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_53/a_132_392# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_45/a_206_368#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_15/a_437_503# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_37/a_651_503#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_39/a_544_485# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_53/a_735_102#
+ prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_45/a_52_123# prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_1/B
+ prbs_generator_syn_17/sky130_fd_sc_hs__nand2_2_3/B prbs_generator_syn_17/sky130_fd_sc_hs__clkbuf_16_1/A
+ prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_21/X prbs_generator_syn_17/sky130_fd_sc_hs__nand2_1_25/B
+ prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_39/a_376_368# prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_63/X
+ prbs_generator_syn_17/m3_13600_3481# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_69/a_1178_124#
+ prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_21/a_138_385# prbs_generator_syn_17/sky130_fd_sc_hs__nor2b_1_8/Y
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_19/a_1178_124# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_49/a_27_74#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_45/a_437_503# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_27/a_651_503#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_71/a_1141_508# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_65/a_651_503#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_29/a_544_485# prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_3/a_138_385#
+ prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_55/X prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_43/a_735_102#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_41/a_1034_424# prbs_generator_syn_17/sky130_fd_sc_hs__nand2_1_9/B
+ prbs_generator_syn_17/sky130_fd_sc_hs__nor2b_1_9/Y prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_59/a_1034_424#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_39/a_1141_508# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_33/a_1226_296#
+ prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_49/a_52_123# prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_47/Y
+ prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_43/Y prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_4/a_651_503#
+ prbs_generator_syn_17/sky130_fd_sc_hs__nand2_1_49/B prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_19/A
+ prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_11/a_138_385# prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_5/X
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_63/a_206_368# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_17/a_651_503#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_19/a_544_485# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_55/a_651_503#
+ prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_9/Y prbs_generator_syn_17/sky130_fd_sc_hs__nand2_1_17/B
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_57/a_544_485# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_67/a_696_458#
+ prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_35/X prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_19/a_27_74#
+ prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_45/a_222_392# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_32/a_1226_296#
+ prbs_generator_syn_17/sky130_fd_sc_hs__nand2_1_43/B prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_25/A
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_1/a_206_368# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_49/a_1226_296#
+ prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_1/a_112_119# prbs_generator_syn_17/sky130_fd_sc_hs__or2_1_1/X
+ prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_59/a_376_368# prbs_generator_syn_17/sky130_fd_sc_hs__nand2_1_19/B
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_5/a_696_458# prbs_generator_syn_17/sky130_fd_sc_hs__nor2b_1_1/Y
+ prbs_generator_syn_17/sky130_fd_sc_hs__nor2b_1_5/a_278_368# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_17/a_1178_124#
+ prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_39/X prbs_generator_syn_17/m3_13600_5433#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_63/a_437_503# prbs_generator_syn_17/sky130_fd_sc_hs__nand2_2_5/B
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_23/a_735_102# prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_53/A
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_61/a_735_102# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_57/a_1034_424#
+ prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_63/B prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_37/a_1141_508#
+ prbs_generator_syn_17/sky130_fd_sc_hs__nand2_1_47/B prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_29/X
+ prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_65/Y prbs_generator_syn_17/m3_13600_4701#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_1/a_437_503# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_67/a_1178_124#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_9/a_735_102# prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_13/a_132_392#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_15/a_1178_124# prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_15/A
+ prbs_generator_syn_17/sky130_fd_sc_hs__nand2_1_1/B prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_43/B
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_35/a_651_503# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_8/D
+ prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_29/A prbs_generator_syn_17/sky130_fd_sc_hs__nand2_1_7/B
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_13/a_735_102# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_47/a_696_458#
+ prbs_generator_syn_17/sky130_fd_sc_hs__nand2_1_31/B prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_51/a_735_102#
+ prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_59/X prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_35/a_1141_508#
+ prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_25/a_222_392# prbs_generator_syn_17/sky130_fd_sc_hs__sdlclkp_2_1/a_288_48#
+ prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_55/B prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_17/B
+ prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_43/A prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_7/A
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_65/a_1178_124# prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_59/Y
+ prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_41/X prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_21/a_230_79#
+ prbs_generator_syn_17/sky130_fd_sc_hs__nand2_1_57/a_117_74# prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_1/a_222_392#
+ prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_19/B prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_35/a_293_74#
+ prbs_generator_syn_17/sky130_fd_sc_hs__nand2_1_23/a_117_74# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_73/a_206_368#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_25/a_651_503# prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_1/a_138_385#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_37/a_696_458# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_67/a_544_485#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_43/a_27_74# prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_9/X
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_55/a_1034_424# prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_39/a_112_119#
+ prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_15/a_222_392# prbs_generator_syn_17/sky130_fd_sc_hs__conb_1_1/HI
+ prbs_generator_syn_17/sky130_fd_sc_hs__nand2_1_23/B prbs_generator_syn_17/sky130_fd_sc_hs__nand2_1_53/B
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_9/a_1178_124# prbs_generator_syn_17/sky130_fd_sc_hs__nor2b_1_4/A
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_47/a_1226_296# prbs_generator_syn_17/m3_13600_11045#
+ prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_17/X prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_29/a_376_368#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_5/a_544_485# prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_3/X
+ prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_31/a_132_392# prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_61/A
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_15/a_651_503# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_73/a_437_503#
+ prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_25/a_230_79# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_27/a_696_458#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_65/a_696_458# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_33/a_735_102#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_71/a_735_102# prbs_generator_syn_17/m3_13600_7263#
+ prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_43/a_222_392# prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_50/Y
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_8/a_1178_124# prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_53/B
+ prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_19/a_376_368# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_63/a_1178_124#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_4/a_696_458# prbs_generator_syn_17/sky130_fd_sc_hs__nor2b_1_4/a_278_368#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_13/a_1178_124# prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_61/a_132_392#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_53/a_206_368# prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_21/a_52_123#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_45/a_651_503# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_17/a_696_458#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_47/a_544_485# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_55/a_696_458#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_21/a_735_102# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_37/a_27_74#
+ prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_61/B prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_61/X
+ prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_59/a_112_119# prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_31/A
+ prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_33/a_222_392# prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_29/a_230_79#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_45/a_1226_296# prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_9/a_132_392#
+ prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_5/A prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_57/Y
+ prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_31/X prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_51/a_27_74#
+ prbs_generator_syn_17/sky130_fd_sc_hs__nor2b_1_8/a_27_112# prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_47/a_376_368#
+ prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_53/a_293_74# prbs_generator_syn_17/sky130_fd_sc_hs__nand2_1_43/a_117_74#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_8/a_735_102# prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_21/a_293_74#
+ prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_39/a_138_385# prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_63/Y
+ prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_51/a_132_392# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_43/a_206_368#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_53/a_437_503# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_37/a_544_485#
+ prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_57/X prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_53/a_1034_424#
+ prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_25/a_52_123# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_33/a_1141_508#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_63/Q prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_23/a_222_392#
+ prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_63/a_222_392# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_7/a_1178_124#
+ prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_53/X prbs_generator_syn_17/sky130_fd_sc_hs__nand2_2_5/Y
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_61/a_1178_124# prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_1/a_230_79#
+ prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_43/a_230_79# prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_11/a_230_79#
+ prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_41/a_132_392# prbs_generator_syn_17/sky130_fd_sc_hs__nand2_1_13/a_117_74#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_43/a_437_503# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_27/a_544_485#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_63/a_651_503# prbs_generator_syn_17/sky130_fd_sc_hs__nand2_1_7/a_117_74#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_35/a_696_458# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_65/a_544_485#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_51/a_1034_424# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_41/a_735_102#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_32/a_1141_508# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_49/a_1141_508#
+ prbs_generator_syn_17/sky130_fd_sc_hs__nand2_1_55/B prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_53/a_222_392#
+ prbs_generator_syn_17/sky130_fd_sc_hs__sdlclkp_2_1/a_114_112# prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_9/a_293_74#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_43/a_1226_296# prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_29/a_52_123#
+ prbs_generator_syn_17/sky130_fd_sc_hs__nand2_1_37/B prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_1/a_651_503#
+ prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_27/a_376_368# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_4/a_544_485#
+ prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_67/a_376_368# prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_27/X
+ prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_1/X prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_59/a_138_385#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_29/a_1178_124# prbs_generator_syn_17/m3_13600_2871#
+ prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_5/a_230_79# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_23/a_206_368#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_61/a_206_368# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_17/a_544_485#
+ prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_15/a_230_79# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_25/a_696_458#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_55/a_544_485# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_32/a_735_102#
+ prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_29/a_293_74# prbs_generator_syn_17/sky130_fd_sc_hs__nand2_1_17/a_117_74#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_69/a_1034_424# prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_29/a_112_119#
+ prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_37/X prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_31/B
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_19/a_1034_424# prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_33/A
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_9/a_206_368# prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_57/a_376_368#
+ prbs_generator_syn_17/sky130_fd_sc_hs__sdlclkp_2_1/a_706_317# prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_11/B
+ prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_1/a_52_123# prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_39/B
+ prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_21/a_132_392# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_13/a_206_368#
+ prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_43/a_52_123# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_51/a_206_368#
+ prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_47/X prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_23/a_437_503#
+ prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_11/a_52_123# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_61/a_437_503#
+ prbs_generator_syn_17/sky130_fd_sc_hs__nor2b_1_7/Y prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_51/A
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_15/a_696_458# prbs_generator_syn_17/sky130_fd_sc_hs__nor2b_1_5/Y
+ prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_9/a_230_79# prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_25/X
+ prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_19/a_112_119# prbs_generator_syn_17/sky130_fd_sc_hs__nand2_1_45/B
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_5/a_1178_124# prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_19/a_230_79#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_41/a_1226_296# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_59/a_1226_296#
+ prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_63/a_230_79# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_51/Q
+ prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_7/a_132_392# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_9/a_437_503#
+ prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_46/a_376_368# prbs_generator_syn_17/sky130_fd_sc_hs__nand2_1_33/a_117_74#
+ prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_11/a_293_74# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_27/a_1178_124#
+ prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_11/a_132_392# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_13/a_437_503#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_51/a_437_503# prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_5/a_52_123#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_35/a_544_485# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_73/a_651_503#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_45/a_696_458# prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_15/a_52_123#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_47/a_1141_508# prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_47/a_112_119#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_4/a_1178_124# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_17/a_1034_424#
+ prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_23/B prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_37/a_376_368#
+ prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_15/B prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_7/Y
+ prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_29/a_138_385# prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_33/a_230_79#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_25/a_1178_124# prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_47/a_293_74#
+ prbs_generator_syn_17/sky130_fd_sc_hs__nand2_1_37/a_117_74# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_33/a_206_368#
+ prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_15/a_293_74# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_71/a_206_368#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_25/a_544_485# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_67/a_1034_424#
+ prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_13/a_222_392# prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_9/a_52_123#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_15/a_1034_424# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_57/a_1226_296#
+ prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_19/a_52_123# prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_23/X
+ prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_63/a_52_123# prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_19/a_138_385#
+ prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_9/a_376_368# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_21/a_206_368#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_33/a_437_503# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_71/a_437_503#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_53/a_651_503# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_15/a_544_485#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_63/a_696_458# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_65/a_1034_424#
+ prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_19/a_293_74# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_45/a_1141_508#
+ prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_27/a_112_119# prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_67/a_112_119#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_1/a_1178_124# prbs_generator_syn_17/sky130_fd_sc_hs__conb_1_1/a_21_290#
+ prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_63/a_293_74# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_8/a_206_368#
+ prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_17/a_376_368# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_63/a_27_74#
+ prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_21/A prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_55/a_376_368#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_1/a_696_458# prbs_generator_syn_17/sky130_fd_sc_hs__nor2b_1_1/a_278_368#
+ prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_47/a_138_385# prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_33/a_52_123#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_9/a_1034_424# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_21/a_437_503#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_1/a_27_74# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_43/a_651_503#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_1/Q prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_45/a_544_485#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_69/a_735_102# prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_57/a_112_119#
+ prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_31/a_222_392# prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_13/A
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_55/a_1226_296# prbs_generator_syn_17/sky130_fd_sc_hs__nand2_2_5/a_27_74#
+ prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_53/a_230_79# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_8/a_437_503#
+ prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_67/a_293_74# prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_33/a_293_74#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_7/a_735_102# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_23/a_1178_124#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_41/a_206_368# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_8/a_1034_424#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_63/a_1034_424# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_59/a_735_102#
+ prbs_generator_syn_17/sky130_fd_sc_hs__nand2_1_5/B prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_43/a_1141_508#
+ prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_46/a_112_119# prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_61/a_222_392#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_13/a_1034_424# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_73/a_1178_124#
+ prbs_generator_syn_17/sky130_fd_sc_hs__nand2_1_27/B prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_13/B
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_57/a_27_74# prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_57/a_230_79#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_21/a_1178_124# prbs_generator_syn_17/sky130_fd_sc_hs__nor2b_1_1/a_27_112#
+ prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_27/a_138_385# prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_23/a_230_79#
+ prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_67/a_138_385# prbs_generator_syn_17/sky130_fd_sc_hs__nand2_1_41/B
+ prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_9/a_222_392# prbs_generator_syn_17/sky130_fd_sc_hs__nand2_1_27/a_117_74#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_32/a_206_368# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_23/a_651_503#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_41/a_437_503# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_73/a_27_74#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_61/a_651_503# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_63/a_544_485#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_49/a_735_102# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_73/a_696_458#
+ prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_37/a_112_119# prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_51/a_222_392#
+ prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_43/X prbs_generator_syn_17/sky130_fd_sc_hs__nand2_2_1/B
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_9/a_651_503# prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_53/a_52_123#
+ prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_49/X prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_25/a_376_368#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_1/a_544_485# prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_65/a_376_368#
+ prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_57/a_138_385# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_27/a_27_74#
+ prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_39/a_132_392# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_7/a_1034_424#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_13/a_651_503# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_32/a_437_503#
+ prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_27/a_230_79# prbs_generator_syn_17/m3_13600_12265#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_51/a_651_503# prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_59/B
+ prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_47/A prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_61/a_1034_424#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_41/a_1141_508# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_59/a_1141_508#
+ prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_41/a_222_392# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_53/a_1226_296#
+ prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_3/A prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_71/a_1178_124#
+ prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_9/a_112_119# prbs_generator_syn_17/sky130_fd_sc_hs__nand2_1_3/a_117_74#
+ prbs_generator_syn_17/m3_13600_8483# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_39/a_1178_124#
+ prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_57/a_52_123# prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_46/a_138_385#
+ prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_23/a_52_123# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_67/a_27_74#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_53/a_696_458# prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_17/a_112_119#
+ prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_11/A prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_55/a_112_119#
+ prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_1/A prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_51/a_1226_296#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_29/a_1034_424# prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_59/A
+ prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_23/A prbs_generator_syn_17/sky130_fd_sc_hs__nand2_1_39/B
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_5/a_27_74# prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_57/a_293_74#
+ prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_37/a_138_385# prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_59/a_132_392#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_33/a_651_503# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_71/a_651_503#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_43/a_696_458# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_73/a_544_485#
+ prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_27/a_52_123# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_57/a_1141_508#
+ prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_21/a_222_392# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_35/a_27_74#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_69/a_1226_296# prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_37/B
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_19/a_1226_296# prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_35/a_376_368#
+ prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_47/a_230_79# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_37/a_1178_124#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_5/a_1034_424# prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_49/a_132_392#
+ prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_7/a_222_392# prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_27/a_293_74#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_21/a_651_503# prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_9/a_138_385#
+ prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_11/a_222_392# prbs_generator_syn_17/m3_13600_14095#
+ prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_50/A prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_27/a_1034_424#
+ prbs_generator_syn_17/sky130_fd_sc_hs__nand2_1_13/B prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_8/a_651_503#
+ prbs_generator_syn_17/m3_13600_9703# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_35/a_1178_124#
+ prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_17/a_138_385# prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_55/a_138_385#
+ prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_7/a_230_79# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_4/a_1034_424#
+ prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_7/a_376_368# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_69/a_206_368#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_23/a_696_458# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_53/a_544_485#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_39/a_735_102# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_61/a_696_458#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_55/a_1141_508# prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_25/a_112_119#
+ prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_65/a_112_119# prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_43/a_293_74#
+ prbs_generator_syn_17/sky130_fd_sc_hs__nand2_1_57/B prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_25/a_1034_424#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_7/a_206_368# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_17/a_1226_296#
+ prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_15/a_376_368# prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_53/a_376_368#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_9/a_696_458# prbs_generator_syn_17/m3_13600_431#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_45/a_27_74# prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_47/a_52_123#
+ prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_29/a_132_392# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_59/a_206_368#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_69/a_437_503# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_41/a_651_503#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_43/a_544_485# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_13/a_696_458#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_29/a_735_102# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_51/a_696_458#
+ prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_61/Y prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_67/a_1226_296#
+ prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_5/a_132_392# prbs_generator_syn_17/sky130_fd_sc_hs__and2b_2_1/a_198_48#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_7/a_437_503# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_15/a_1226_296#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_69/a_27_74# prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_46/a_293_74#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_1/a_1034_424# prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_19/a_132_392#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_49/a_206_368# prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_7/a_52_123#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_59/a_437_503# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_32/a_651_503#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_7/a_27_74# prbs_generator_syn_17/sky130_fd_sc_hs__nand2_2_1/a_27_74#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_19/a_735_102# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_57/a_735_102#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_65/a_1226_296# prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_37/A
+ prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_33/a_376_368# prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_37/a_230_79#
+ prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_25/a_138_385# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_39/a_27_74#
+ prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_65/a_138_385# prbs_generator_syn_17/sky130_fd_sc_hs__nor2b_1_9/a_278_368#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_49/a_437_503# prbs_generator_syn_17/sky130_fd_sc_hs__and2b_2_1/a_505_74#
+ prbs_generator_syn_17/sky130_fd_sc_hs__nand2_1_51/a_117_74# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_23/a_544_485#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_33/a_696_458# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_61/a_544_485#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_9/a_1226_296# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_53/a_1141_508#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_71/a_696_458# prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_35/a_112_119#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_23/a_1034_424# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_9/a_544_485#
+ prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_63/a_376_368# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_33/a_1178_124#
+ prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_5/a_376_368# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_13/a_544_485#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_73/a_1034_424# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_21/a_696_458#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_51/a_544_485# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_8/a_1226_296#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_51/a_1141_508# prbs_generator_syn_17/sky130_fd_sc_hs__nand2_1_55/a_117_74#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_21/a_1034_424# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_63/a_1226_296#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_23/a_27_74# prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_7/a_112_119#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_13/a_1226_296# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_8/a_696_458#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_32/a_1178_124# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_49/a_1178_124#
+ prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_37/a_52_123# prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_27/a_132_392#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_71/Q prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_67/a_735_102#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_69/a_1141_508# prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_15/a_112_119#
+ prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_53/a_112_119# prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_39/a_222_392#
+ prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_55/a_230_79# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_19/a_1141_508#
+ prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_37/a_293_74# prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_43/a_376_368#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_5/a_735_102# prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_35/a_138_385#
+ prbs_generator_syn_17/sky130_fd_sc_hs__sdlclkp_2_1/a_114_424# prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_57/a_132_392#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_71/a_1034_424# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_7/a_1226_296#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_33/a_544_485# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_41/a_696_458#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_71/a_544_485# prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_21/B
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_61/a_1226_296# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_39/a_1034_424#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_17/a_27_74# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_9/a_27_74#
+ prbs_generator_syn_17/sky130_fd_sc_hs__nor2b_1_5/a_27_112# prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_47/a_132_392#
+ prbs_generator_syn_17/sky130_fd_sc_hs__nor2b_1_8/a_278_368# prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_9/B
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_39/a_206_368# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_33/a_27_74#
+ prbs_generator_syn_17/sky130_fd_sc_hs__nand2_1_41/a_117_74# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_69/a_651_503#
+ prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_51/a_293_74# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_21/a_544_485#
+ prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_7/a_138_385# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_32/a_696_458#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_47/a_735_102# prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_33/a_112_119#
+ prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_59/a_222_392# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_17/a_1141_508#
+ prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_55/a_52_123# prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_3/a_293_74#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_7/a_651_503# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_29/a_1226_296#
+ prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_23/a_376_368# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_8/a_544_485#
+ prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_47/B prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_47/a_1178_124#
+ prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_15/a_138_385# prbs_generator_syn_17/sky130_fd_sc_hs__sdlclkp_2_1/a_1195_374#
+ prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_53/a_138_385# prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_37/a_132_392#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_29/a_206_368# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_39/a_437_503#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_59/a_651_503# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_37/a_735_102#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_67/a_1141_508# prbs_generator_syn_17/sky130_fd_sc_hs__and2b_2_1/a_27_74#
+ prbs_generator_syn_17/sky130_fd_sc_hs__conb_1_1/a_165_290# prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_55/a_293_74#
+ prbs_generator_syn_17/sky130_fd_sc_hs__nand2_1_45/a_117_74# prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_63/a_112_119#
+ prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_49/a_222_392# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_37/a_1034_424#
+ prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_23/a_293_74# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_15/a_1141_508#
+ prbs_generator_syn_17/sky130_fd_sc_hs__nand2_1_5/a_117_74# prbs_generator_syn_17/m3_13600_13485#
+ prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_5/a_112_119# prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_13/a_376_368#
+ prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_51/a_376_368# prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_7/a_293_74#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_19/a_206_368# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_57/a_206_368#
+ prbs_generator_syn_17/sky130_fd_sc_hs__sdlclkp_2_1/a_318_74# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_29/a_437_503#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_49/a_651_503# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_25/a_27_74#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_5/a_1226_296# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_41/a_544_485#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_27/a_735_102# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_65/a_1141_508#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_65/a_735_102# prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_3/a_230_79#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_35/a_1034_424# prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_13/a_230_79#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_41/a_27_74# prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_3/a_132_392#
+ prbs_generator_syn_17/sky130_fd_sc_hs__nand2_1_49/a_117_74# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_27/a_1226_296#
+ prbs_generator_syn_17/sky130_fd_sc_hs__nand2_1_15/a_117_74# prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_41/a_376_368#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_45/a_1178_124# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_4/a_735_102#
+ prbs_generator_syn_17/sky130_fd_sc_hs__nand2_1_9/a_117_74# prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_33/a_138_385#
+ prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_17/a_132_392# prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_55/a_132_392#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_9/a_1141_508# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_19/a_437_503#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_57/a_437_503# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_4/a_1226_296#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_32/a_544_485# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_17/a_735_102#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_55/a_735_102# prbs_generator_syn_17/m3_13600_2261#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_65/a_27_74# prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_29/a_222_392#
+ prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_43/a_112_119# prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_19/X
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_25/a_1226_296# prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_31/a_376_368#
+ prbs_generator_syn_17/sky130_fd_sc_hs__or2_1_1/a_63_368# prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_17/a_230_79#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_4/a_27_74# prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_61/a_230_79#
+ prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_63/a_138_385# prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_5/a_222_392#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_8/a_1141_508# prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_41/a_293_74#
+ prbs_generator_syn_17/sky130_fd_sc_hs__nand2_1_31/a_117_74# prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_5/a_138_385#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_63/a_1141_508# prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_19/a_222_392#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_13/a_1141_508# prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_3/a_52_123#
+ prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_13/a_52_123# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_43/a_1178_124#
+ prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_61/a_376_368# prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_35/a_132_392#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_67/a_206_368# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_1/a_1226_296#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_69/a_696_458# prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_31/a_230_79#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_35/a_735_102# prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_23/a_112_119#
+ prbs_generator_syn_17/sky130_fd_sc_hs__nand2_1_35/a_117_74# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_59/a_27_74#
+ prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_13/a_293_74# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_5/a_206_368#
+ prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_50/a_376_368# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_7/a_696_458#
+ prbs_generator_syn_17/sky130_fd_sc_hs__nor2b_1_7/a_278_368# prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_17/a_52_123#
+ prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_43/a_138_385# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_7/a_1141_508#
+ prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_61/a_52_123# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_67/a_437_503#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_61/a_1141_508# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_25/a_735_102#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_59/a_696_458# prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_13/a_112_119#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_33/a_1034_424# prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_51/a_112_119#
+ prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_35/a_230_79# prbs_generator_syn_17/m3_13600_4091#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_23/a_1226_296# prbs_generator_syn_17/sky130_fd_sc_hs__nand2_1_39/a_117_74#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_29/a_27_74# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_5/a_437_503#
+ prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_17/a_293_74# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_41/a_1178_124#
+ prbs_generator_syn_17/sky130_fd_sc_hs__or2_1_1/a_152_368# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_59/a_1178_124#
+ prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_61/a_293_74# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_47/a_206_368#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_39/a_651_503# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_49/a_696_458#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_15/a_735_102# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_32/a_1034_424#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_73/a_1226_296# prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_27/a_222_392#
+ prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_41/a_112_119# prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_31/a_52_123#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_49/a_1034_424# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_29/a_1141_508#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_21/a_1226_296# prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_39/a_230_79#
+ prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_23/a_138_385# prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_51/a_230_79#
+ prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_45/a_132_392# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_37/a_206_368#
+ prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_65/a_293_74# prbs_generator_syn_17/sky130_fd_sc_hs__nand2_1_53/a_117_74#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_47/a_437_503# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_29/a_651_503#
+ prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_31/a_293_74# prbs_generator_syn_17/sky130_fd_sc_hs__nand2_1_21/a_117_74#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_69/a_544_485# prbs_generator_syn_17/sky130_fd_sc_hs__clkbuf_16_1/a_114_74#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_45/a_735_102# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_13/a_27_74#
+ prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_31/a_112_119# prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_57/a_222_392#
+ prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_35/a_52_123# prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_21/a_376_368#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_7/a_544_485# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_57/a_1178_124#
+ prbs_generator_syn_17/m3_13600_6043# prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_13/a_138_385#
+ prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_51/a_138_385# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_5/a_1141_508#
+ prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_3/a_376_368# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_27/a_206_368#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_65/a_206_368# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_37/a_437_503#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_19/a_651_503# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_57/a_651_503#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_59/a_544_485# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_71/a_1226_296#
+ prbs_generator_syn_17/sky130_fd_sc_hs__nand2_1_25/a_117_74# prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_61/a_112_119#
+ prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_47/a_222_392# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_27/a_1141_508#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_53/a_27_74# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_4/a_206_368#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_39/a_1226_296# prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_11/a_376_368#
+ prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_39/a_52_123# prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_41/a_138_385#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_4/a_1141_508# prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_25/a_132_392#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_17/a_206_368# prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_41/A
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_55/a_206_368# prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_51/a_52_123#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_27/a_437_503# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_65/a_437_503#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_49/a_544_485# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_63/a_735_102#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_47/a_1034_424# prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_50/a_112_119#
+ prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_37/a_222_392# prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_59/a_230_79#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_25/a_1141_508# prbs_generator_syn_17/sky130_fd_sc_hs__nor2b_1_4/a_27_112#
+ prbs_generator_syn_17/sky130_fd_sc_hs__sdlclkp_2_1/a_685_81# prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_1/a_132_392#
+ prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_39/a_293_74# prbs_generator_syn_17/sky130_fd_sc_hs__nand2_1_29/a_117_74#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_4/a_437_503# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_55/a_1178_124#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_21/a_27_74# prbs_generator_syn_17/m3_13600_12875#
+ prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_50/a_293_74# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_1/a_735_102#
+ prbs_generator_syn_17/sky130_fd_sc_hs__xnor2_1_31/a_138_385# prbs_generator_syn_17/sky130_fd_sc_hs__a22o_1_15/a_132_392#
+ prbs_generator_syn_17/sky130_fd_sc_hs__nand2_1_1/a_117_74# prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_17/a_437_503#
+ prbs_generator_syn_17/sky130_fd_sc_hs__dfxtp_4_55/a_437_503# prbs_generator_syn
Xprbs_generator_syn_28 prbs_generator_syn_31/clk prbs_generator_syn_31/rst prbs_generator_syn_29/cke
+ sky130_fd_sc_hs__conb_1_265/LO sky130_fd_sc_hs__conb_1_265/LO sky130_fd_sc_hs__conb_1_265/LO
+ sky130_fd_sc_hs__conb_1_265/LO prbs_generator_syn_31/eqn[8] prbs_generator_syn_31/eqn[8]
+ sky130_fd_sc_hs__conb_1_265/LO sky130_fd_sc_hs__conb_1_265/LO sky130_fd_sc_hs__conb_1_265/LO
+ sky130_fd_sc_hs__conb_1_265/LO sky130_fd_sc_hs__conb_1_241/LO sky130_fd_sc_hs__conb_1_241/LO
+ sky130_fd_sc_hs__conb_1_241/LO sky130_fd_sc_hs__conb_1_241/LO sky130_fd_sc_hs__conb_1_241/LO
+ sky130_fd_sc_hs__conb_1_241/LO sky130_fd_sc_hs__conb_1_241/LO sky130_fd_sc_hs__conb_1_241/LO
+ prbs_generator_syn_29/eqn[2] prbs_generator_syn_29/eqn[2] prbs_generator_syn_29/eqn[2]
+ prbs_generator_syn_29/eqn[1] prbs_generator_syn_29/eqn[2] prbs_generator_syn_29/eqn[1]
+ sky130_fd_sc_hs__conb_1_263/LO sky130_fd_sc_hs__conb_1_263/HI sky130_fd_sc_hs__conb_1_263/LO
+ sky130_fd_sc_hs__conb_1_263/HI sky130_fd_sc_hs__conb_1_263/LO sky130_fd_sc_hs__conb_1_263/HI
+ sky130_fd_sc_hs__conb_1_263/LO sky130_fd_sc_hs__conb_1_263/HI prbs_generator_syn_29/eqn[31]
+ prbs_generator_syn_29/eqn[31] prbs_generator_syn_29/eqn[31] prbs_generator_syn_29/eqn[28]
+ prbs_generator_syn_29/eqn[28] prbs_generator_syn_29/eqn[28] prbs_generator_syn_29/eqn[28]
+ prbs_generator_syn_29/eqn[28] prbs_generator_syn_29/eqn[28] prbs_generator_syn_29/eqn[22]
+ prbs_generator_syn_29/eqn[22] prbs_generator_syn_29/eqn[20] prbs_generator_syn_29/eqn[22]
+ prbs_generator_syn_29/eqn[22] prbs_generator_syn_29/eqn[22] prbs_generator_syn_29/eqn[22]
+ prbs_generator_syn_23/eqn[0] prbs_generator_syn_23/eqn[0] prbs_generator_syn_23/eqn[0]
+ prbs_generator_syn_23/eqn[0] prbs_generator_syn_23/eqn[0] prbs_generator_syn_23/eqn[0]
+ prbs_generator_syn_29/eqn[9] prbs_generator_syn_29/eqn[9] prbs_generator_syn_29/eqn[9]
+ prbs_generator_syn_29/eqn[9] prbs_generator_syn_29/eqn[9] prbs_generator_syn_29/eqn[9]
+ prbs_generator_syn_29/eqn[9] prbs_generator_syn_29/eqn[2] prbs_generator_syn_29/eqn[1]
+ prbs_generator_syn_29/eqn[2] prbs_generator_syn_31/inj_err prbs_generator_syn_29/eqn[31]
+ prbs_generator_syn_29/eqn[31] hr_16t4_mux_top_1/din[6] DVSS: DVDD: prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_1/a_293_74#
+ prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_15/X prbs_generator_syn_29/sky130_fd_sc_hs__nand2_1_35/B
+ prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_51/Y prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_9/A
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_9/CLK prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_47/a_27_74#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_37/a_1226_296# prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_3/B
+ prbs_generator_syn_29/sky130_fd_sc_hs__nor2b_1_7/a_27_112# prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_29/B
+ prbs_generator_syn_29/sky130_fd_sc_hs__sdlclkp_2_1/a_580_74# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_1/a_1141_508#
+ prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_5/Y prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_41/a_230_79#
+ prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_61/a_138_385# prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_43/a_132_392#
+ prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_3/a_222_392# prbs_generator_syn_29/sky130_fd_sc_hs__nor2b_1_9/a_27_112#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_61/a_27_74# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_35/a_206_368#
+ prbs_generator_syn_29/sky130_fd_sc_hs__nand2_2_3/Y prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_25/B
+ prbs_generator_syn_29/sky130_fd_sc_hs__nand2_1_11/a_117_74# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_67/a_651_503#
+ prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_45/X prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_39/a_696_458#
+ prbs_generator_syn_29/sky130_fd_sc_hs__sdlclkp_2_1/a_1198_74# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_45/a_1034_424#
+ prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_17/a_222_392# prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_55/a_222_392#
+ prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_53/Y prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_35/A
+ prbs_generator_syn_29/m3_13600_1651# prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_59/a_52_123#
+ prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_5/a_293_74# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_35/a_1226_296#
+ prbs_generator_syn_29/sky130_fd_sc_hs__nand2_1_51/B prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_5/a_651_503#
+ prbs_generator_syn_29/sky130_fd_sc_hs__nand2_1_21/B prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_8/a_27_74#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_15/a_27_74# prbs_generator_syn_29/sky130_fd_sc_hs__and2b_2_1/X
+ prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_13/X prbs_generator_syn_29/sky130_fd_sc_hs__nand2_2_3/a_27_74#
+ prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_50/a_138_385# prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_33/a_132_392#
+ prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_1/a_376_368# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_25/a_206_368#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_35/a_437_503# prbs_generator_syn_29/sky130_fd_sc_hs__sdlclkp_2_1/a_708_451#
+ prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_45/a_230_79# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_29/a_696_458#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_32/a_27_74# prbs_generator_syn_29/sky130_fd_sc_hs__nor2b_1_4/Y
+ prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_59/a_293_74# prbs_generator_syn_29/sky130_fd_sc_hs__nand2_1_47/a_117_74#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_73/a_735_102# prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_21/a_112_119#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_23/a_1141_508# prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_25/a_293_74#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_7/Q prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_3/a_112_119#
+ prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_35/B prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_51/X
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_53/a_1178_124# prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_23/a_132_392#
+ prbs_generator_syn_29/sky130_fd_sc_hs__nand2_1_3/B prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_15/a_206_368#
+ prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_63/a_132_392# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_55/a_27_74#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_25/a_437_503# prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_41/a_52_123#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_47/a_651_503# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_73/a_1141_508#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_19/a_696_458# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_57/a_696_458#
+ prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_7/X prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_43/a_1034_424#
+ prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_55/A prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_11/a_112_119#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_21/a_1141_508# prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_35/a_222_392#
+ prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_49/a_230_79# prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_67/Y
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_71/a_27_74# prbs_generator_syn_29/sky130_fd_sc_hs__nand2_1_33/B
+ prbs_generator_syn_29/sky130_fd_sc_hs__conb_1_1/LO prbs_generator_syn_29/sky130_fd_sc_hs__nand2_1_19/a_117_74#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_51/a_1178_124# prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_33/X
+ prbs_generator_syn_29/sky130_fd_sc_hs__nand2_1_29/B prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_41/Y
+ prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_53/a_132_392# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_45/a_206_368#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_15/a_437_503# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_37/a_651_503#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_39/a_544_485# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_53/a_735_102#
+ prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_45/a_52_123# prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_1/B
+ prbs_generator_syn_29/sky130_fd_sc_hs__nand2_2_3/B prbs_generator_syn_29/sky130_fd_sc_hs__clkbuf_16_1/A
+ prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_21/X prbs_generator_syn_29/sky130_fd_sc_hs__nand2_1_25/B
+ prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_39/a_376_368# prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_63/X
+ prbs_generator_syn_29/m3_13600_3481# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_69/a_1178_124#
+ prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_21/a_138_385# prbs_generator_syn_29/sky130_fd_sc_hs__nor2b_1_8/Y
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_19/a_1178_124# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_49/a_27_74#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_45/a_437_503# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_27/a_651_503#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_71/a_1141_508# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_65/a_651_503#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_29/a_544_485# prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_3/a_138_385#
+ prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_55/X prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_43/a_735_102#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_41/a_1034_424# prbs_generator_syn_29/sky130_fd_sc_hs__nand2_1_9/B
+ prbs_generator_syn_29/sky130_fd_sc_hs__nor2b_1_9/Y prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_59/a_1034_424#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_39/a_1141_508# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_33/a_1226_296#
+ prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_49/a_52_123# prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_47/Y
+ prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_43/Y prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_4/a_651_503#
+ prbs_generator_syn_29/sky130_fd_sc_hs__nand2_1_49/B prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_19/A
+ prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_11/a_138_385# prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_5/X
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_63/a_206_368# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_17/a_651_503#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_19/a_544_485# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_55/a_651_503#
+ prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_9/Y prbs_generator_syn_29/sky130_fd_sc_hs__nand2_1_17/B
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_57/a_544_485# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_67/a_696_458#
+ prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_35/X prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_19/a_27_74#
+ prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_45/a_222_392# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_32/a_1226_296#
+ prbs_generator_syn_29/sky130_fd_sc_hs__nand2_1_43/B prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_25/A
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_1/a_206_368# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_49/a_1226_296#
+ prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_1/a_112_119# prbs_generator_syn_29/sky130_fd_sc_hs__or2_1_1/X
+ prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_59/a_376_368# prbs_generator_syn_29/sky130_fd_sc_hs__nand2_1_19/B
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_5/a_696_458# prbs_generator_syn_29/sky130_fd_sc_hs__nor2b_1_1/Y
+ prbs_generator_syn_29/sky130_fd_sc_hs__nor2b_1_5/a_278_368# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_17/a_1178_124#
+ prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_39/X prbs_generator_syn_29/m3_13600_5433#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_63/a_437_503# prbs_generator_syn_29/sky130_fd_sc_hs__nand2_2_5/B
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_23/a_735_102# prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_53/A
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_61/a_735_102# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_57/a_1034_424#
+ prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_63/B prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_37/a_1141_508#
+ prbs_generator_syn_29/sky130_fd_sc_hs__nand2_1_47/B prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_29/X
+ prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_65/Y prbs_generator_syn_29/m3_13600_4701#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_1/a_437_503# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_67/a_1178_124#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_9/a_735_102# prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_13/a_132_392#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_15/a_1178_124# prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_15/A
+ prbs_generator_syn_29/sky130_fd_sc_hs__nand2_1_1/B prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_43/B
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_35/a_651_503# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_8/D
+ prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_29/A prbs_generator_syn_29/sky130_fd_sc_hs__nand2_1_7/B
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_13/a_735_102# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_47/a_696_458#
+ prbs_generator_syn_29/sky130_fd_sc_hs__nand2_1_31/B prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_51/a_735_102#
+ prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_59/X prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_35/a_1141_508#
+ prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_25/a_222_392# prbs_generator_syn_29/sky130_fd_sc_hs__sdlclkp_2_1/a_288_48#
+ prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_55/B prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_17/B
+ prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_43/A prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_7/A
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_65/a_1178_124# prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_59/Y
+ prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_41/X prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_21/a_230_79#
+ prbs_generator_syn_29/sky130_fd_sc_hs__nand2_1_57/a_117_74# prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_1/a_222_392#
+ prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_19/B prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_35/a_293_74#
+ prbs_generator_syn_29/sky130_fd_sc_hs__nand2_1_23/a_117_74# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_73/a_206_368#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_25/a_651_503# prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_1/a_138_385#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_37/a_696_458# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_67/a_544_485#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_43/a_27_74# prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_9/X
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_55/a_1034_424# prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_39/a_112_119#
+ prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_15/a_222_392# prbs_generator_syn_29/sky130_fd_sc_hs__conb_1_1/HI
+ prbs_generator_syn_29/sky130_fd_sc_hs__nand2_1_23/B prbs_generator_syn_29/sky130_fd_sc_hs__nand2_1_53/B
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_9/a_1178_124# prbs_generator_syn_29/sky130_fd_sc_hs__nor2b_1_4/A
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_47/a_1226_296# prbs_generator_syn_29/m3_13600_11045#
+ prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_17/X prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_29/a_376_368#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_5/a_544_485# prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_3/X
+ prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_31/a_132_392# prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_61/A
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_15/a_651_503# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_73/a_437_503#
+ prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_25/a_230_79# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_27/a_696_458#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_65/a_696_458# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_33/a_735_102#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_71/a_735_102# prbs_generator_syn_29/m3_13600_7263#
+ prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_43/a_222_392# prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_50/Y
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_8/a_1178_124# prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_53/B
+ prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_19/a_376_368# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_63/a_1178_124#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_4/a_696_458# prbs_generator_syn_29/sky130_fd_sc_hs__nor2b_1_4/a_278_368#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_13/a_1178_124# prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_61/a_132_392#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_53/a_206_368# prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_21/a_52_123#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_45/a_651_503# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_17/a_696_458#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_47/a_544_485# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_55/a_696_458#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_21/a_735_102# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_37/a_27_74#
+ prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_61/B prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_61/X
+ prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_59/a_112_119# prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_31/A
+ prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_33/a_222_392# prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_29/a_230_79#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_45/a_1226_296# prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_9/a_132_392#
+ prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_5/A prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_57/Y
+ prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_31/X prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_51/a_27_74#
+ prbs_generator_syn_29/sky130_fd_sc_hs__nor2b_1_8/a_27_112# prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_47/a_376_368#
+ prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_53/a_293_74# prbs_generator_syn_29/sky130_fd_sc_hs__nand2_1_43/a_117_74#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_8/a_735_102# prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_21/a_293_74#
+ prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_39/a_138_385# prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_63/Y
+ prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_51/a_132_392# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_43/a_206_368#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_53/a_437_503# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_37/a_544_485#
+ prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_57/X prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_53/a_1034_424#
+ prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_25/a_52_123# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_33/a_1141_508#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_63/Q prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_23/a_222_392#
+ prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_63/a_222_392# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_7/a_1178_124#
+ prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_53/X prbs_generator_syn_29/sky130_fd_sc_hs__nand2_2_5/Y
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_61/a_1178_124# prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_1/a_230_79#
+ prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_43/a_230_79# prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_11/a_230_79#
+ prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_41/a_132_392# prbs_generator_syn_29/sky130_fd_sc_hs__nand2_1_13/a_117_74#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_43/a_437_503# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_27/a_544_485#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_63/a_651_503# prbs_generator_syn_29/sky130_fd_sc_hs__nand2_1_7/a_117_74#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_35/a_696_458# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_65/a_544_485#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_51/a_1034_424# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_41/a_735_102#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_32/a_1141_508# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_49/a_1141_508#
+ prbs_generator_syn_29/sky130_fd_sc_hs__nand2_1_55/B prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_53/a_222_392#
+ prbs_generator_syn_29/sky130_fd_sc_hs__sdlclkp_2_1/a_114_112# prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_9/a_293_74#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_43/a_1226_296# prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_29/a_52_123#
+ prbs_generator_syn_29/sky130_fd_sc_hs__nand2_1_37/B prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_1/a_651_503#
+ prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_27/a_376_368# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_4/a_544_485#
+ prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_67/a_376_368# prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_27/X
+ prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_1/X prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_59/a_138_385#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_29/a_1178_124# prbs_generator_syn_29/m3_13600_2871#
+ prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_5/a_230_79# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_23/a_206_368#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_61/a_206_368# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_17/a_544_485#
+ prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_15/a_230_79# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_25/a_696_458#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_55/a_544_485# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_32/a_735_102#
+ prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_29/a_293_74# prbs_generator_syn_29/sky130_fd_sc_hs__nand2_1_17/a_117_74#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_69/a_1034_424# prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_29/a_112_119#
+ prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_37/X prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_31/B
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_19/a_1034_424# prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_33/A
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_9/a_206_368# prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_57/a_376_368#
+ prbs_generator_syn_29/sky130_fd_sc_hs__sdlclkp_2_1/a_706_317# prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_11/B
+ prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_1/a_52_123# prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_39/B
+ prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_21/a_132_392# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_13/a_206_368#
+ prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_43/a_52_123# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_51/a_206_368#
+ prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_47/X prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_23/a_437_503#
+ prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_11/a_52_123# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_61/a_437_503#
+ prbs_generator_syn_29/sky130_fd_sc_hs__nor2b_1_7/Y prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_51/A
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_15/a_696_458# prbs_generator_syn_29/sky130_fd_sc_hs__nor2b_1_5/Y
+ prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_9/a_230_79# prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_25/X
+ prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_19/a_112_119# prbs_generator_syn_29/sky130_fd_sc_hs__nand2_1_45/B
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_5/a_1178_124# prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_19/a_230_79#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_41/a_1226_296# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_59/a_1226_296#
+ prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_63/a_230_79# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_51/Q
+ prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_7/a_132_392# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_9/a_437_503#
+ prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_46/a_376_368# prbs_generator_syn_29/sky130_fd_sc_hs__nand2_1_33/a_117_74#
+ prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_11/a_293_74# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_27/a_1178_124#
+ prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_11/a_132_392# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_13/a_437_503#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_51/a_437_503# prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_5/a_52_123#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_35/a_544_485# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_73/a_651_503#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_45/a_696_458# prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_15/a_52_123#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_47/a_1141_508# prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_47/a_112_119#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_4/a_1178_124# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_17/a_1034_424#
+ prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_23/B prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_37/a_376_368#
+ prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_15/B prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_7/Y
+ prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_29/a_138_385# prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_33/a_230_79#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_25/a_1178_124# prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_47/a_293_74#
+ prbs_generator_syn_29/sky130_fd_sc_hs__nand2_1_37/a_117_74# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_33/a_206_368#
+ prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_15/a_293_74# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_71/a_206_368#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_25/a_544_485# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_67/a_1034_424#
+ prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_13/a_222_392# prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_9/a_52_123#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_15/a_1034_424# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_57/a_1226_296#
+ prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_19/a_52_123# prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_23/X
+ prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_63/a_52_123# prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_19/a_138_385#
+ prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_9/a_376_368# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_21/a_206_368#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_33/a_437_503# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_71/a_437_503#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_53/a_651_503# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_15/a_544_485#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_63/a_696_458# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_65/a_1034_424#
+ prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_19/a_293_74# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_45/a_1141_508#
+ prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_27/a_112_119# prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_67/a_112_119#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_1/a_1178_124# prbs_generator_syn_29/sky130_fd_sc_hs__conb_1_1/a_21_290#
+ prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_63/a_293_74# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_8/a_206_368#
+ prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_17/a_376_368# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_63/a_27_74#
+ prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_21/A prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_55/a_376_368#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_1/a_696_458# prbs_generator_syn_29/sky130_fd_sc_hs__nor2b_1_1/a_278_368#
+ prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_47/a_138_385# prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_33/a_52_123#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_9/a_1034_424# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_21/a_437_503#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_1/a_27_74# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_43/a_651_503#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_1/Q prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_45/a_544_485#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_69/a_735_102# prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_57/a_112_119#
+ prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_31/a_222_392# prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_13/A
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_55/a_1226_296# prbs_generator_syn_29/sky130_fd_sc_hs__nand2_2_5/a_27_74#
+ prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_53/a_230_79# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_8/a_437_503#
+ prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_67/a_293_74# prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_33/a_293_74#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_7/a_735_102# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_23/a_1178_124#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_41/a_206_368# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_8/a_1034_424#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_63/a_1034_424# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_59/a_735_102#
+ prbs_generator_syn_29/sky130_fd_sc_hs__nand2_1_5/B prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_43/a_1141_508#
+ prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_46/a_112_119# prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_61/a_222_392#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_13/a_1034_424# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_73/a_1178_124#
+ prbs_generator_syn_29/sky130_fd_sc_hs__nand2_1_27/B prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_13/B
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_57/a_27_74# prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_57/a_230_79#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_21/a_1178_124# prbs_generator_syn_29/sky130_fd_sc_hs__nor2b_1_1/a_27_112#
+ prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_27/a_138_385# prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_23/a_230_79#
+ prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_67/a_138_385# prbs_generator_syn_29/sky130_fd_sc_hs__nand2_1_41/B
+ prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_9/a_222_392# prbs_generator_syn_29/sky130_fd_sc_hs__nand2_1_27/a_117_74#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_32/a_206_368# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_23/a_651_503#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_41/a_437_503# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_73/a_27_74#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_61/a_651_503# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_63/a_544_485#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_49/a_735_102# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_73/a_696_458#
+ prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_37/a_112_119# prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_51/a_222_392#
+ prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_43/X prbs_generator_syn_29/sky130_fd_sc_hs__nand2_2_1/B
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_9/a_651_503# prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_53/a_52_123#
+ prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_49/X prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_25/a_376_368#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_1/a_544_485# prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_65/a_376_368#
+ prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_57/a_138_385# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_27/a_27_74#
+ prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_39/a_132_392# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_7/a_1034_424#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_13/a_651_503# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_32/a_437_503#
+ prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_27/a_230_79# prbs_generator_syn_29/m3_13600_12265#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_51/a_651_503# prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_59/B
+ prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_47/A prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_61/a_1034_424#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_41/a_1141_508# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_59/a_1141_508#
+ prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_41/a_222_392# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_53/a_1226_296#
+ prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_3/A prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_71/a_1178_124#
+ prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_9/a_112_119# prbs_generator_syn_29/sky130_fd_sc_hs__nand2_1_3/a_117_74#
+ prbs_generator_syn_29/m3_13600_8483# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_39/a_1178_124#
+ prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_57/a_52_123# prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_46/a_138_385#
+ prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_23/a_52_123# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_67/a_27_74#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_53/a_696_458# prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_17/a_112_119#
+ prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_11/A prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_55/a_112_119#
+ prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_1/A prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_51/a_1226_296#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_29/a_1034_424# prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_59/A
+ prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_23/A prbs_generator_syn_29/sky130_fd_sc_hs__nand2_1_39/B
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_5/a_27_74# prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_57/a_293_74#
+ prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_37/a_138_385# prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_59/a_132_392#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_33/a_651_503# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_71/a_651_503#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_43/a_696_458# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_73/a_544_485#
+ prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_27/a_52_123# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_57/a_1141_508#
+ prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_21/a_222_392# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_35/a_27_74#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_69/a_1226_296# prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_37/B
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_19/a_1226_296# prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_35/a_376_368#
+ prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_47/a_230_79# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_37/a_1178_124#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_5/a_1034_424# prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_49/a_132_392#
+ prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_7/a_222_392# prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_27/a_293_74#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_21/a_651_503# prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_9/a_138_385#
+ prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_11/a_222_392# prbs_generator_syn_29/m3_13600_14095#
+ prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_50/A prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_27/a_1034_424#
+ prbs_generator_syn_29/sky130_fd_sc_hs__nand2_1_13/B prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_8/a_651_503#
+ prbs_generator_syn_29/m3_13600_9703# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_35/a_1178_124#
+ prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_17/a_138_385# prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_55/a_138_385#
+ prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_7/a_230_79# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_4/a_1034_424#
+ prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_7/a_376_368# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_69/a_206_368#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_23/a_696_458# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_53/a_544_485#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_39/a_735_102# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_61/a_696_458#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_55/a_1141_508# prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_25/a_112_119#
+ prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_65/a_112_119# prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_43/a_293_74#
+ prbs_generator_syn_29/sky130_fd_sc_hs__nand2_1_57/B prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_25/a_1034_424#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_7/a_206_368# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_17/a_1226_296#
+ prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_15/a_376_368# prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_53/a_376_368#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_9/a_696_458# prbs_generator_syn_29/m3_13600_431#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_45/a_27_74# prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_47/a_52_123#
+ prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_29/a_132_392# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_59/a_206_368#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_69/a_437_503# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_41/a_651_503#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_43/a_544_485# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_13/a_696_458#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_29/a_735_102# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_51/a_696_458#
+ prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_61/Y prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_67/a_1226_296#
+ prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_5/a_132_392# prbs_generator_syn_29/sky130_fd_sc_hs__and2b_2_1/a_198_48#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_7/a_437_503# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_15/a_1226_296#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_69/a_27_74# prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_46/a_293_74#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_1/a_1034_424# prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_19/a_132_392#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_49/a_206_368# prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_7/a_52_123#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_59/a_437_503# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_32/a_651_503#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_7/a_27_74# prbs_generator_syn_29/sky130_fd_sc_hs__nand2_2_1/a_27_74#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_19/a_735_102# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_57/a_735_102#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_65/a_1226_296# prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_37/A
+ prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_33/a_376_368# prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_37/a_230_79#
+ prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_25/a_138_385# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_39/a_27_74#
+ prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_65/a_138_385# prbs_generator_syn_29/sky130_fd_sc_hs__nor2b_1_9/a_278_368#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_49/a_437_503# prbs_generator_syn_29/sky130_fd_sc_hs__and2b_2_1/a_505_74#
+ prbs_generator_syn_29/sky130_fd_sc_hs__nand2_1_51/a_117_74# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_23/a_544_485#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_33/a_696_458# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_61/a_544_485#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_9/a_1226_296# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_53/a_1141_508#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_71/a_696_458# prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_35/a_112_119#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_23/a_1034_424# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_9/a_544_485#
+ prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_63/a_376_368# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_33/a_1178_124#
+ prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_5/a_376_368# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_13/a_544_485#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_73/a_1034_424# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_21/a_696_458#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_51/a_544_485# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_8/a_1226_296#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_51/a_1141_508# prbs_generator_syn_29/sky130_fd_sc_hs__nand2_1_55/a_117_74#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_21/a_1034_424# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_63/a_1226_296#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_23/a_27_74# prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_7/a_112_119#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_13/a_1226_296# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_8/a_696_458#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_32/a_1178_124# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_49/a_1178_124#
+ prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_37/a_52_123# prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_27/a_132_392#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_71/Q prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_67/a_735_102#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_69/a_1141_508# prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_15/a_112_119#
+ prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_53/a_112_119# prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_39/a_222_392#
+ prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_55/a_230_79# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_19/a_1141_508#
+ prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_37/a_293_74# prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_43/a_376_368#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_5/a_735_102# prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_35/a_138_385#
+ prbs_generator_syn_29/sky130_fd_sc_hs__sdlclkp_2_1/a_114_424# prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_57/a_132_392#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_71/a_1034_424# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_7/a_1226_296#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_33/a_544_485# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_41/a_696_458#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_71/a_544_485# prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_21/B
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_61/a_1226_296# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_39/a_1034_424#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_17/a_27_74# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_9/a_27_74#
+ prbs_generator_syn_29/sky130_fd_sc_hs__nor2b_1_5/a_27_112# prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_47/a_132_392#
+ prbs_generator_syn_29/sky130_fd_sc_hs__nor2b_1_8/a_278_368# prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_9/B
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_39/a_206_368# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_33/a_27_74#
+ prbs_generator_syn_29/sky130_fd_sc_hs__nand2_1_41/a_117_74# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_69/a_651_503#
+ prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_51/a_293_74# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_21/a_544_485#
+ prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_7/a_138_385# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_32/a_696_458#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_47/a_735_102# prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_33/a_112_119#
+ prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_59/a_222_392# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_17/a_1141_508#
+ prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_55/a_52_123# prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_3/a_293_74#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_7/a_651_503# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_29/a_1226_296#
+ prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_23/a_376_368# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_8/a_544_485#
+ prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_47/B prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_47/a_1178_124#
+ prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_15/a_138_385# prbs_generator_syn_29/sky130_fd_sc_hs__sdlclkp_2_1/a_1195_374#
+ prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_53/a_138_385# prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_37/a_132_392#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_29/a_206_368# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_39/a_437_503#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_59/a_651_503# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_37/a_735_102#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_67/a_1141_508# prbs_generator_syn_29/sky130_fd_sc_hs__and2b_2_1/a_27_74#
+ prbs_generator_syn_29/sky130_fd_sc_hs__conb_1_1/a_165_290# prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_55/a_293_74#
+ prbs_generator_syn_29/sky130_fd_sc_hs__nand2_1_45/a_117_74# prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_63/a_112_119#
+ prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_49/a_222_392# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_37/a_1034_424#
+ prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_23/a_293_74# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_15/a_1141_508#
+ prbs_generator_syn_29/sky130_fd_sc_hs__nand2_1_5/a_117_74# prbs_generator_syn_29/m3_13600_13485#
+ prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_5/a_112_119# prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_13/a_376_368#
+ prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_51/a_376_368# prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_7/a_293_74#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_19/a_206_368# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_57/a_206_368#
+ prbs_generator_syn_29/sky130_fd_sc_hs__sdlclkp_2_1/a_318_74# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_29/a_437_503#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_49/a_651_503# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_25/a_27_74#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_5/a_1226_296# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_41/a_544_485#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_27/a_735_102# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_65/a_1141_508#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_65/a_735_102# prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_3/a_230_79#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_35/a_1034_424# prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_13/a_230_79#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_41/a_27_74# prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_3/a_132_392#
+ prbs_generator_syn_29/sky130_fd_sc_hs__nand2_1_49/a_117_74# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_27/a_1226_296#
+ prbs_generator_syn_29/sky130_fd_sc_hs__nand2_1_15/a_117_74# prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_41/a_376_368#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_45/a_1178_124# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_4/a_735_102#
+ prbs_generator_syn_29/sky130_fd_sc_hs__nand2_1_9/a_117_74# prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_33/a_138_385#
+ prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_17/a_132_392# prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_55/a_132_392#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_9/a_1141_508# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_19/a_437_503#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_57/a_437_503# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_4/a_1226_296#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_32/a_544_485# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_17/a_735_102#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_55/a_735_102# prbs_generator_syn_29/m3_13600_2261#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_65/a_27_74# prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_29/a_222_392#
+ prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_43/a_112_119# prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_19/X
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_25/a_1226_296# prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_31/a_376_368#
+ prbs_generator_syn_29/sky130_fd_sc_hs__or2_1_1/a_63_368# prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_17/a_230_79#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_4/a_27_74# prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_61/a_230_79#
+ prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_63/a_138_385# prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_5/a_222_392#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_8/a_1141_508# prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_41/a_293_74#
+ prbs_generator_syn_29/sky130_fd_sc_hs__nand2_1_31/a_117_74# prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_5/a_138_385#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_63/a_1141_508# prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_19/a_222_392#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_13/a_1141_508# prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_3/a_52_123#
+ prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_13/a_52_123# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_43/a_1178_124#
+ prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_61/a_376_368# prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_35/a_132_392#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_67/a_206_368# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_1/a_1226_296#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_69/a_696_458# prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_31/a_230_79#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_35/a_735_102# prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_23/a_112_119#
+ prbs_generator_syn_29/sky130_fd_sc_hs__nand2_1_35/a_117_74# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_59/a_27_74#
+ prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_13/a_293_74# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_5/a_206_368#
+ prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_50/a_376_368# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_7/a_696_458#
+ prbs_generator_syn_29/sky130_fd_sc_hs__nor2b_1_7/a_278_368# prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_17/a_52_123#
+ prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_43/a_138_385# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_7/a_1141_508#
+ prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_61/a_52_123# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_67/a_437_503#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_61/a_1141_508# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_25/a_735_102#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_59/a_696_458# prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_13/a_112_119#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_33/a_1034_424# prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_51/a_112_119#
+ prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_35/a_230_79# prbs_generator_syn_29/m3_13600_4091#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_23/a_1226_296# prbs_generator_syn_29/sky130_fd_sc_hs__nand2_1_39/a_117_74#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_29/a_27_74# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_5/a_437_503#
+ prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_17/a_293_74# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_41/a_1178_124#
+ prbs_generator_syn_29/sky130_fd_sc_hs__or2_1_1/a_152_368# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_59/a_1178_124#
+ prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_61/a_293_74# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_47/a_206_368#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_39/a_651_503# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_49/a_696_458#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_15/a_735_102# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_32/a_1034_424#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_73/a_1226_296# prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_27/a_222_392#
+ prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_41/a_112_119# prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_31/a_52_123#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_49/a_1034_424# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_29/a_1141_508#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_21/a_1226_296# prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_39/a_230_79#
+ prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_23/a_138_385# prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_51/a_230_79#
+ prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_45/a_132_392# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_37/a_206_368#
+ prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_65/a_293_74# prbs_generator_syn_29/sky130_fd_sc_hs__nand2_1_53/a_117_74#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_47/a_437_503# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_29/a_651_503#
+ prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_31/a_293_74# prbs_generator_syn_29/sky130_fd_sc_hs__nand2_1_21/a_117_74#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_69/a_544_485# prbs_generator_syn_29/sky130_fd_sc_hs__clkbuf_16_1/a_114_74#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_45/a_735_102# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_13/a_27_74#
+ prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_31/a_112_119# prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_57/a_222_392#
+ prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_35/a_52_123# prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_21/a_376_368#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_7/a_544_485# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_57/a_1178_124#
+ prbs_generator_syn_29/m3_13600_6043# prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_13/a_138_385#
+ prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_51/a_138_385# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_5/a_1141_508#
+ prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_3/a_376_368# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_27/a_206_368#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_65/a_206_368# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_37/a_437_503#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_19/a_651_503# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_57/a_651_503#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_59/a_544_485# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_71/a_1226_296#
+ prbs_generator_syn_29/sky130_fd_sc_hs__nand2_1_25/a_117_74# prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_61/a_112_119#
+ prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_47/a_222_392# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_27/a_1141_508#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_53/a_27_74# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_4/a_206_368#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_39/a_1226_296# prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_11/a_376_368#
+ prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_39/a_52_123# prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_41/a_138_385#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_4/a_1141_508# prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_25/a_132_392#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_17/a_206_368# prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_41/A
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_55/a_206_368# prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_51/a_52_123#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_27/a_437_503# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_65/a_437_503#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_49/a_544_485# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_63/a_735_102#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_47/a_1034_424# prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_50/a_112_119#
+ prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_37/a_222_392# prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_59/a_230_79#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_25/a_1141_508# prbs_generator_syn_29/sky130_fd_sc_hs__nor2b_1_4/a_27_112#
+ prbs_generator_syn_29/sky130_fd_sc_hs__sdlclkp_2_1/a_685_81# prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_1/a_132_392#
+ prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_39/a_293_74# prbs_generator_syn_29/sky130_fd_sc_hs__nand2_1_29/a_117_74#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_4/a_437_503# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_55/a_1178_124#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_21/a_27_74# prbs_generator_syn_29/m3_13600_12875#
+ prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_50/a_293_74# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_1/a_735_102#
+ prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_31/a_138_385# prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_15/a_132_392#
+ prbs_generator_syn_29/sky130_fd_sc_hs__nand2_1_1/a_117_74# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_17/a_437_503#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_55/a_437_503# prbs_generator_syn
Xsky130_fd_sc_hs__conb_1_8 DVSS: DVDD: DVDD: DVSS: prbs_generator_syn_3/eqn[8] sky130_fd_sc_hs__conb_1_9/HI
+ sky130_fd_sc_hs__conb_1_9/a_165_290# sky130_fd_sc_hs__conb_1_9/a_21_290# sky130_fd_sc_hs__conb_1
Xsky130_fd_sc_hs__buf_2_104 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__buf_2_105/A sky130_fd_sc_hs__buf_2_105/X
+ sky130_fd_sc_hs__buf_2_105/a_21_260# sky130_fd_sc_hs__buf_2
Xsky130_fd_sc_hs__buf_2_115 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__buf_2_115/A sky130_fd_sc_hs__buf_2_115/X
+ sky130_fd_sc_hs__buf_2_115/a_21_260# sky130_fd_sc_hs__buf_2
Xsky130_fd_sc_hs__buf_2_126 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__buf_2_127/A sky130_fd_sc_hs__buf_2_15/A
+ sky130_fd_sc_hs__buf_2_127/a_21_260# sky130_fd_sc_hs__buf_2
Xsky130_fd_sc_hs__buf_2_137 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__buf_2_137/A sky130_fd_sc_hs__buf_2_137/X
+ sky130_fd_sc_hs__buf_2_137/a_21_260# sky130_fd_sc_hs__buf_2
Xsky130_fd_sc_hs__buf_2_148 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__buf_2_149/A sky130_fd_sc_hs__buf_2_153/A
+ sky130_fd_sc_hs__buf_2_149/a_21_260# sky130_fd_sc_hs__buf_2
Xsky130_fd_sc_hs__buf_2_159 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__buf_2_159/A sky130_fd_sc_hs__buf_2_159/X
+ sky130_fd_sc_hs__buf_2_159/a_21_260# sky130_fd_sc_hs__buf_2
Xsky130_fd_sc_hs__einvp_2_16 DVSS: DVDD: DVDD: DVSS: dout_n sky130_fd_sc_hs__einvp_2_9/A
+ sky130_fd_sc_hs__dlrtp_1_5/Q sky130_fd_sc_hs__einvp_2_17/a_263_323# sky130_fd_sc_hs__einvp_2_17/a_36_74#
+ sky130_fd_sc_hs__einvp_2_17/a_27_368# sky130_fd_sc_hs__einvp_2
Xsky130_fd_sc_hs__einvp_2_27 DVSS: DVDD: DVDD: DVSS: dout_n sky130_fd_sc_hs__einvp_2_9/A
+ sky130_fd_sc_hs__einvp_2_27/TE sky130_fd_sc_hs__einvp_2_27/a_263_323# sky130_fd_sc_hs__einvp_2_27/a_36_74#
+ sky130_fd_sc_hs__einvp_2_27/a_27_368# sky130_fd_sc_hs__einvp_2
Xsky130_fd_sc_hs__einvp_2_38 DVSS: DVDD: DVDD: DVSS: dout_n sky130_fd_sc_hs__buf_8_1/A
+ sky130_fd_sc_hs__buf_2_17/X sky130_fd_sc_hs__einvp_2_39/a_263_323# sky130_fd_sc_hs__einvp_2_39/a_36_74#
+ sky130_fd_sc_hs__einvp_2_39/a_27_368# sky130_fd_sc_hs__einvp_2
Xsky130_fd_sc_hs__einvp_2_49 DVSS: DVDD: DVDD: DVSS: dout_n sky130_fd_sc_hs__buf_8_1/A
+ sky130_fd_sc_hs__einvp_2_49/TE sky130_fd_sc_hs__einvp_2_49/a_263_323# sky130_fd_sc_hs__einvp_2_49/a_36_74#
+ sky130_fd_sc_hs__einvp_2_49/a_27_368# sky130_fd_sc_hs__einvp_2
Xsky130_fd_sc_hs__conb_1_15 DVSS: DVDD: DVDD: DVSS: prbs_generator_syn_9/eqn[16] sky130_fd_sc_hs__conb_1_15/HI
+ sky130_fd_sc_hs__conb_1_15/a_165_290# sky130_fd_sc_hs__conb_1_15/a_21_290# sky130_fd_sc_hs__conb_1
Xsky130_fd_sc_hs__conb_1_26 DVSS: DVDD: DVDD: DVSS: prbs_generator_syn_5/eqn[13] sky130_fd_sc_hs__conb_1_27/HI
+ sky130_fd_sc_hs__conb_1_27/a_165_290# sky130_fd_sc_hs__conb_1_27/a_21_290# sky130_fd_sc_hs__conb_1
Xsky130_fd_sc_hs__conb_1_37 DVSS: DVDD: DVDD: DVSS: prbs_generator_syn_3/eqn[28] sky130_fd_sc_hs__conb_1_37/HI
+ sky130_fd_sc_hs__conb_1_37/a_165_290# sky130_fd_sc_hs__conb_1_37/a_21_290# sky130_fd_sc_hs__conb_1
Xsky130_fd_sc_hs__conb_1_48 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__conb_1_49/LO
+ sky130_fd_sc_hs__conb_1_49/HI sky130_fd_sc_hs__conb_1_49/a_165_290# sky130_fd_sc_hs__conb_1_49/a_21_290#
+ sky130_fd_sc_hs__conb_1
Xsky130_fd_sc_hs__conb_1_59 DVSS: DVDD: DVDD: DVSS: prbs_generator_syn_11/eqn[9] sky130_fd_sc_hs__conb_1_59/HI
+ sky130_fd_sc_hs__conb_1_59/a_165_290# sky130_fd_sc_hs__conb_1_59/a_21_290# sky130_fd_sc_hs__conb_1
Xsky130_fd_sc_hs__inv_4_11 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__inv_4_11/Y sky130_fd_sc_hs__inv_4_11/A
+ sky130_fd_sc_hs__inv_4
Xsky130_fd_sc_hs__inv_4_22 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__inv_4_23/Y sky130_fd_sc_hs__inv_4_23/A
+ sky130_fd_sc_hs__inv_4
Xsky130_fd_sc_hs__inv_4_33 DVSS: DVDD: DVDD: DVSS: osc_core_1/pi1_r[1] osc_core_1/pi1_l[1]
+ sky130_fd_sc_hs__inv_4
Xsky130_fd_sc_hs__inv_4_44 DVSS: DVDD: DVDD: DVSS: osc_core_1/pi3_r[3] osc_core_1/pi3_l[3]
+ sky130_fd_sc_hs__inv_4
Xsky130_fd_sc_hs__inv_4_55 DVSS: DVDD: DVDD: DVSS: osc_core_1/pi4_r[0] osc_core_1/pi4_l[0]
+ sky130_fd_sc_hs__inv_4
Xsky130_fd_sc_hs__inv_4_66 DVSS: DVDD: DVDD: DVSS: hr_16t4_mux_top_3/din[1] hr_16t4_mux_top_1/din[1]
+ sky130_fd_sc_hs__inv_4
Xsky130_fd_sc_hs__inv_4_77 DVSS: DVDD: DVDD: DVSS: hr_16t4_mux_top_3/din[10] prbs_generator_syn_19/out
+ sky130_fd_sc_hs__inv_4
Xsky130_fd_sc_hs__inv_4_88 DVSS: DVDD: DVDD: DVSS: hr_16t4_mux_top_3/din[0] hr_16t4_mux_top_1/din[0]
+ sky130_fd_sc_hs__inv_4
Xsky130_fd_sc_hs__dlrtp_1_17 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__dlrtp_1_17/Q
+ sky130_fd_sc_hs__dlrtp_1_9/GATE sky130_fd_sc_hs__conb_1_119/HI sky130_fd_sc_hs__dlrtp_1_17/D
+ sky130_fd_sc_hs__dlrtp_1_17/a_216_424# sky130_fd_sc_hs__dlrtp_1_17/a_759_508# sky130_fd_sc_hs__dlrtp_1_17/a_565_74#
+ sky130_fd_sc_hs__dlrtp_1_17/a_27_424# sky130_fd_sc_hs__dlrtp_1_17/a_1045_74# sky130_fd_sc_hs__dlrtp_1_17/a_643_74#
+ sky130_fd_sc_hs__dlrtp_1_17/a_817_48# sky130_fd_sc_hs__dlrtp_1_17/a_568_392# sky130_fd_sc_hs__dlrtp_1_17/a_363_74#
+ sky130_fd_sc_hs__dlrtp_1_17/a_769_74# sky130_fd_sc_hs__dlrtp_1
Xsky130_fd_sc_hs__dlrtp_1_28 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__dlrtp_1_29/Q
+ sky130_fd_sc_hs__clkbuf_2_3/A sky130_fd_sc_hs__conb_1_123/HI sky130_fd_sc_hs__dlrtp_1_29/D
+ sky130_fd_sc_hs__dlrtp_1_29/a_216_424# sky130_fd_sc_hs__dlrtp_1_29/a_759_508# sky130_fd_sc_hs__dlrtp_1_29/a_565_74#
+ sky130_fd_sc_hs__dlrtp_1_29/a_27_424# sky130_fd_sc_hs__dlrtp_1_29/a_1045_74# sky130_fd_sc_hs__dlrtp_1_29/a_643_74#
+ sky130_fd_sc_hs__dlrtp_1_29/a_817_48# sky130_fd_sc_hs__dlrtp_1_29/a_568_392# sky130_fd_sc_hs__dlrtp_1_29/a_363_74#
+ sky130_fd_sc_hs__dlrtp_1_29/a_769_74# sky130_fd_sc_hs__dlrtp_1
Xsky130_fd_sc_hs__dlrtp_1_39 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__dlrtp_1_39/Q
+ sky130_fd_sc_hs__clkbuf_16_53/A sky130_fd_sc_hs__conb_1_123/HI sky130_fd_sc_hs__buf_2_30/X
+ sky130_fd_sc_hs__dlrtp_1_39/a_216_424# sky130_fd_sc_hs__dlrtp_1_39/a_759_508# sky130_fd_sc_hs__dlrtp_1_39/a_565_74#
+ sky130_fd_sc_hs__dlrtp_1_39/a_27_424# sky130_fd_sc_hs__dlrtp_1_39/a_1045_74# sky130_fd_sc_hs__dlrtp_1_39/a_643_74#
+ sky130_fd_sc_hs__dlrtp_1_39/a_817_48# sky130_fd_sc_hs__dlrtp_1_39/a_568_392# sky130_fd_sc_hs__dlrtp_1_39/a_363_74#
+ sky130_fd_sc_hs__dlrtp_1_39/a_769_74# sky130_fd_sc_hs__dlrtp_1
Xsky130_fd_sc_hs__clkbuf_16_60 DVSS: DVDD: DVDD: DVSS: qr_4t1_mux_top_3/clk_I sky130_fd_sc_hs__einvn_2_1/Z
+ sky130_fd_sc_hs__clkbuf_16_61/a_114_74# sky130_fd_sc_hs__clkbuf_16
Xsky130_fd_sc_hs__clkbuf_16_71 DVSS: DVDD: DVDD: DVSS: prbs_generator_syn_13/rst prbs_generator_syn_19/rst
+ sky130_fd_sc_hs__clkbuf_16_71/a_114_74# sky130_fd_sc_hs__clkbuf_16
Xsky130_fd_sc_hs__clkbuf_16_82 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__nor2_4_1/A
+ sky130_fd_sc_hs__clkbuf_4_113/X sky130_fd_sc_hs__clkbuf_16_83/a_114_74# sky130_fd_sc_hs__clkbuf_16
Xsky130_fd_sc_hs__clkbuf_16_93 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__clkbuf_16_93/X
+ sky130_fd_sc_hs__clkbuf_4_115/X sky130_fd_sc_hs__clkbuf_16_93/a_114_74# sky130_fd_sc_hs__clkbuf_16
Xsky130_fd_sc_hs__clkbuf_8_101 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__clkinv_8_19/A
+ rst sky130_fd_sc_hs__clkbuf_8_101/a_125_368# sky130_fd_sc_hs__clkbuf_8
Xsky130_fd_sc_hs__nand2_2_12 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__buf_2_87/A sky130_fd_sc_hs__buf_8_3/X
+ sky130_fd_sc_hs__inv_4_21/Y sky130_fd_sc_hs__nand2_2_13/a_27_74# sky130_fd_sc_hs__nand2_2
Xsky130_fd_sc_hs__nand2_2_23 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__nand2_2_23/Y
+ sky130_fd_sc_hs__nor4_2_1/C sky130_fd_sc_hs__nor4_2_1/B sky130_fd_sc_hs__nand2_2_23/a_27_74#
+ sky130_fd_sc_hs__nand2_2
Xsky130_fd_sc_hs__conb_1_209 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__conb_1_209/LO
+ sky130_fd_sc_hs__conb_1_209/HI sky130_fd_sc_hs__conb_1_209/a_165_290# sky130_fd_sc_hs__conb_1_209/a_21_290#
+ sky130_fd_sc_hs__conb_1
Xprbs_generator_syn_1 prbs_generator_syn_9/clk prbs_generator_syn_9/rst prbs_generator_syn_1/cke
+ sky130_fd_sc_hs__conb_1_41/LO prbs_generator_syn_5/eqn[5] prbs_generator_syn_5/eqn[1]
+ prbs_generator_syn_5/eqn[1] prbs_generator_syn_5/eqn[1] prbs_generator_syn_5/eqn[1]
+ sky130_fd_sc_hs__conb_1_41/HI sky130_fd_sc_hs__conb_1_41/LO sky130_fd_sc_hs__conb_1_41/LO
+ sky130_fd_sc_hs__conb_1_41/LO sky130_fd_sc_hs__conb_1_41/LO prbs_generator_syn_1/eqn[31]
+ prbs_generator_syn_5/eqn[13] sky130_fd_sc_hs__conb_1_27/HI prbs_generator_syn_5/eqn[13]
+ sky130_fd_sc_hs__conb_1_27/HI prbs_generator_syn_5/eqn[13] sky130_fd_sc_hs__conb_1_27/HI
+ prbs_generator_syn_3/eqn[9] prbs_generator_syn_3/eqn[20] prbs_generator_syn_3/eqn[20]
+ prbs_generator_syn_3/eqn[20] prbs_generator_syn_3/eqn[20] prbs_generator_syn_3/eqn[28]
+ prbs_generator_syn_3/eqn[28] sky130_fd_sc_hs__conb_1_37/HI sky130_fd_sc_hs__conb_1_37/HI
+ prbs_generator_syn_3/eqn[30] sky130_fd_sc_hs__conb_1_45/HI prbs_generator_syn_3/eqn[30]
+ sky130_fd_sc_hs__conb_1_45/HI prbs_generator_syn_3/eqn[30] prbs_generator_syn_1/eqn[31]
+ prbs_generator_syn_1/eqn[30] prbs_generator_syn_1/eqn[30] prbs_generator_syn_1/eqn[30]
+ prbs_generator_syn_1/eqn[30] prbs_generator_syn_1/eqn[30] prbs_generator_syn_1/eqn[30]
+ prbs_generator_syn_1/eqn[30] prbs_generator_syn_1/eqn[30] sky130_fd_sc_hs__conb_1_3/LO
+ sky130_fd_sc_hs__conb_1_3/LO sky130_fd_sc_hs__conb_1_3/HI sky130_fd_sc_hs__conb_1_3/LO
+ sky130_fd_sc_hs__conb_1_3/LO sky130_fd_sc_hs__conb_1_3/LO sky130_fd_sc_hs__conb_1_3/LO
+ sky130_fd_sc_hs__conb_1_3/LO sky130_fd_sc_hs__conb_1_3/LO prbs_generator_syn_1/eqn[9]
+ prbs_generator_syn_1/eqn[9] prbs_generator_syn_1/eqn[9] prbs_generator_syn_1/eqn[9]
+ prbs_generator_syn_1/eqn[9] prbs_generator_syn_1/eqn[8] prbs_generator_syn_1/eqn[8]
+ prbs_generator_syn_1/eqn[8] prbs_generator_syn_1/eqn[8] prbs_generator_syn_1/eqn[8]
+ prbs_generator_syn_1/eqn[8] prbs_generator_syn_1/eqn[8] prbs_generator_syn_1/eqn[1]
+ prbs_generator_syn_3/eqn[9] prbs_generator_syn_9/inj_err prbs_generator_syn_1/eqn[31]
+ prbs_generator_syn_1/eqn[31] prbs_generator_syn_1/out DVSS: DVDD: prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_1/a_293_74#
+ prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_15/X prbs_generator_syn_1/sky130_fd_sc_hs__nand2_1_35/B
+ prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_51/Y prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_9/A
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_9/CLK prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_47/a_27_74#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_37/a_1226_296# prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_3/B
+ prbs_generator_syn_1/sky130_fd_sc_hs__nor2b_1_7/a_27_112# prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_29/B
+ prbs_generator_syn_1/sky130_fd_sc_hs__sdlclkp_2_1/a_580_74# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_1/a_1141_508#
+ prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_5/Y prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_41/a_230_79#
+ prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_61/a_138_385# prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_43/a_132_392#
+ prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_3/a_222_392# prbs_generator_syn_1/sky130_fd_sc_hs__nor2b_1_9/a_27_112#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_61/a_27_74# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_35/a_206_368#
+ prbs_generator_syn_1/sky130_fd_sc_hs__nand2_2_3/Y prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_25/B
+ prbs_generator_syn_1/sky130_fd_sc_hs__nand2_1_11/a_117_74# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_67/a_651_503#
+ prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_45/X prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_39/a_696_458#
+ prbs_generator_syn_1/sky130_fd_sc_hs__sdlclkp_2_1/a_1198_74# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_45/a_1034_424#
+ prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_17/a_222_392# prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_55/a_222_392#
+ prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_53/Y prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_35/A
+ prbs_generator_syn_1/m3_13600_1651# prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_59/a_52_123#
+ prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_5/a_293_74# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_35/a_1226_296#
+ prbs_generator_syn_1/sky130_fd_sc_hs__nand2_1_51/B prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_5/a_651_503#
+ prbs_generator_syn_1/sky130_fd_sc_hs__nand2_1_21/B prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_8/a_27_74#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_15/a_27_74# prbs_generator_syn_1/sky130_fd_sc_hs__and2b_2_1/X
+ prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_13/X prbs_generator_syn_1/sky130_fd_sc_hs__nand2_2_3/a_27_74#
+ prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_50/a_138_385# prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_33/a_132_392#
+ prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_1/a_376_368# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_25/a_206_368#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_35/a_437_503# prbs_generator_syn_1/sky130_fd_sc_hs__sdlclkp_2_1/a_708_451#
+ prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_45/a_230_79# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_29/a_696_458#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_32/a_27_74# prbs_generator_syn_1/sky130_fd_sc_hs__nor2b_1_4/Y
+ prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_59/a_293_74# prbs_generator_syn_1/sky130_fd_sc_hs__nand2_1_47/a_117_74#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_73/a_735_102# prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_21/a_112_119#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_23/a_1141_508# prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_25/a_293_74#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_7/Q prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_3/a_112_119#
+ prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_35/B prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_51/X
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_53/a_1178_124# prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_23/a_132_392#
+ prbs_generator_syn_1/sky130_fd_sc_hs__nand2_1_3/B prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_15/a_206_368#
+ prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_63/a_132_392# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_55/a_27_74#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_25/a_437_503# prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_41/a_52_123#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_47/a_651_503# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_73/a_1141_508#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_19/a_696_458# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_57/a_696_458#
+ prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_7/X prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_43/a_1034_424#
+ prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_55/A prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_11/a_112_119#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_21/a_1141_508# prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_35/a_222_392#
+ prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_49/a_230_79# prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_67/Y
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_71/a_27_74# prbs_generator_syn_1/sky130_fd_sc_hs__nand2_1_33/B
+ prbs_generator_syn_1/sky130_fd_sc_hs__conb_1_1/LO prbs_generator_syn_1/sky130_fd_sc_hs__nand2_1_19/a_117_74#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_51/a_1178_124# prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_33/X
+ prbs_generator_syn_1/sky130_fd_sc_hs__nand2_1_29/B prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_41/Y
+ prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_53/a_132_392# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_45/a_206_368#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_15/a_437_503# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_37/a_651_503#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_39/a_544_485# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_53/a_735_102#
+ prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_45/a_52_123# prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_1/B
+ prbs_generator_syn_1/sky130_fd_sc_hs__nand2_2_3/B prbs_generator_syn_1/sky130_fd_sc_hs__clkbuf_16_1/A
+ prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_21/X prbs_generator_syn_1/sky130_fd_sc_hs__nand2_1_25/B
+ prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_39/a_376_368# prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_63/X
+ prbs_generator_syn_1/m3_13600_3481# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_69/a_1178_124#
+ prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_21/a_138_385# prbs_generator_syn_1/sky130_fd_sc_hs__nor2b_1_8/Y
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_19/a_1178_124# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_49/a_27_74#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_45/a_437_503# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_27/a_651_503#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_71/a_1141_508# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_65/a_651_503#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_29/a_544_485# prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_3/a_138_385#
+ prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_55/X prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_43/a_735_102#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_41/a_1034_424# prbs_generator_syn_1/sky130_fd_sc_hs__nand2_1_9/B
+ prbs_generator_syn_1/sky130_fd_sc_hs__nor2b_1_9/Y prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_59/a_1034_424#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_39/a_1141_508# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_33/a_1226_296#
+ prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_49/a_52_123# prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_47/Y
+ prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_43/Y prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_4/a_651_503#
+ prbs_generator_syn_1/sky130_fd_sc_hs__nand2_1_49/B prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_19/A
+ prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_11/a_138_385# prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_5/X
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_63/a_206_368# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_17/a_651_503#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_19/a_544_485# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_55/a_651_503#
+ prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_9/Y prbs_generator_syn_1/sky130_fd_sc_hs__nand2_1_17/B
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_57/a_544_485# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_67/a_696_458#
+ prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_35/X prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_19/a_27_74#
+ prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_45/a_222_392# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_32/a_1226_296#
+ prbs_generator_syn_1/sky130_fd_sc_hs__nand2_1_43/B prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_25/A
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_1/a_206_368# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_49/a_1226_296#
+ prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_1/a_112_119# prbs_generator_syn_1/sky130_fd_sc_hs__or2_1_1/X
+ prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_59/a_376_368# prbs_generator_syn_1/sky130_fd_sc_hs__nand2_1_19/B
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_5/a_696_458# prbs_generator_syn_1/sky130_fd_sc_hs__nor2b_1_1/Y
+ prbs_generator_syn_1/sky130_fd_sc_hs__nor2b_1_5/a_278_368# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_17/a_1178_124#
+ prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_39/X prbs_generator_syn_1/m3_13600_5433#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_63/a_437_503# prbs_generator_syn_1/sky130_fd_sc_hs__nand2_2_5/B
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_23/a_735_102# prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_53/A
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_61/a_735_102# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_57/a_1034_424#
+ prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_63/B prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_37/a_1141_508#
+ prbs_generator_syn_1/sky130_fd_sc_hs__nand2_1_47/B prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_29/X
+ prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_65/Y prbs_generator_syn_1/m3_13600_4701#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_1/a_437_503# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_67/a_1178_124#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_9/a_735_102# prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_13/a_132_392#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_15/a_1178_124# prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_15/A
+ prbs_generator_syn_1/sky130_fd_sc_hs__nand2_1_1/B prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_43/B
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_35/a_651_503# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_8/D
+ prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_29/A prbs_generator_syn_1/sky130_fd_sc_hs__nand2_1_7/B
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_13/a_735_102# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_47/a_696_458#
+ prbs_generator_syn_1/sky130_fd_sc_hs__nand2_1_31/B prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_51/a_735_102#
+ prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_59/X prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_35/a_1141_508#
+ prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_25/a_222_392# prbs_generator_syn_1/sky130_fd_sc_hs__sdlclkp_2_1/a_288_48#
+ prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_55/B prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_17/B
+ prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_43/A prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_7/A
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_65/a_1178_124# prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_59/Y
+ prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_41/X prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_21/a_230_79#
+ prbs_generator_syn_1/sky130_fd_sc_hs__nand2_1_57/a_117_74# prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_1/a_222_392#
+ prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_19/B prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_35/a_293_74#
+ prbs_generator_syn_1/sky130_fd_sc_hs__nand2_1_23/a_117_74# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_73/a_206_368#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_25/a_651_503# prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_1/a_138_385#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_37/a_696_458# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_67/a_544_485#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_43/a_27_74# prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_9/X
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_55/a_1034_424# prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_39/a_112_119#
+ prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_15/a_222_392# prbs_generator_syn_1/sky130_fd_sc_hs__conb_1_1/HI
+ prbs_generator_syn_1/sky130_fd_sc_hs__nand2_1_23/B prbs_generator_syn_1/sky130_fd_sc_hs__nand2_1_53/B
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_9/a_1178_124# prbs_generator_syn_1/sky130_fd_sc_hs__nor2b_1_4/A
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_47/a_1226_296# prbs_generator_syn_1/m3_13600_11045#
+ prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_17/X prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_29/a_376_368#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_5/a_544_485# prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_3/X
+ prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_31/a_132_392# prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_61/A
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_15/a_651_503# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_73/a_437_503#
+ prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_25/a_230_79# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_27/a_696_458#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_65/a_696_458# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_33/a_735_102#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_71/a_735_102# prbs_generator_syn_1/m3_13600_7263#
+ prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_43/a_222_392# prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_50/Y
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_8/a_1178_124# prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_53/B
+ prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_19/a_376_368# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_63/a_1178_124#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_4/a_696_458# prbs_generator_syn_1/sky130_fd_sc_hs__nor2b_1_4/a_278_368#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_13/a_1178_124# prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_61/a_132_392#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_53/a_206_368# prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_21/a_52_123#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_45/a_651_503# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_17/a_696_458#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_47/a_544_485# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_55/a_696_458#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_21/a_735_102# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_37/a_27_74#
+ prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_61/B prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_61/X
+ prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_59/a_112_119# prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_31/A
+ prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_33/a_222_392# prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_29/a_230_79#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_45/a_1226_296# prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_9/a_132_392#
+ prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_5/A prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_57/Y
+ prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_31/X prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_51/a_27_74#
+ prbs_generator_syn_1/sky130_fd_sc_hs__nor2b_1_8/a_27_112# prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_47/a_376_368#
+ prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_53/a_293_74# prbs_generator_syn_1/sky130_fd_sc_hs__nand2_1_43/a_117_74#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_8/a_735_102# prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_21/a_293_74#
+ prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_39/a_138_385# prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_63/Y
+ prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_51/a_132_392# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_43/a_206_368#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_53/a_437_503# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_37/a_544_485#
+ prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_57/X prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_53/a_1034_424#
+ prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_25/a_52_123# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_33/a_1141_508#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_63/Q prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_23/a_222_392#
+ prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_63/a_222_392# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_7/a_1178_124#
+ prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_53/X prbs_generator_syn_1/sky130_fd_sc_hs__nand2_2_5/Y
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_61/a_1178_124# prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_1/a_230_79#
+ prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_43/a_230_79# prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_11/a_230_79#
+ prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_41/a_132_392# prbs_generator_syn_1/sky130_fd_sc_hs__nand2_1_13/a_117_74#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_43/a_437_503# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_27/a_544_485#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_63/a_651_503# prbs_generator_syn_1/sky130_fd_sc_hs__nand2_1_7/a_117_74#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_35/a_696_458# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_65/a_544_485#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_51/a_1034_424# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_41/a_735_102#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_32/a_1141_508# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_49/a_1141_508#
+ prbs_generator_syn_1/sky130_fd_sc_hs__nand2_1_55/B prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_53/a_222_392#
+ prbs_generator_syn_1/sky130_fd_sc_hs__sdlclkp_2_1/a_114_112# prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_9/a_293_74#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_43/a_1226_296# prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_29/a_52_123#
+ prbs_generator_syn_1/sky130_fd_sc_hs__nand2_1_37/B prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_1/a_651_503#
+ prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_27/a_376_368# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_4/a_544_485#
+ prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_67/a_376_368# prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_27/X
+ prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_1/X prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_59/a_138_385#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_29/a_1178_124# prbs_generator_syn_1/m3_13600_2871#
+ prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_5/a_230_79# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_23/a_206_368#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_61/a_206_368# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_17/a_544_485#
+ prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_15/a_230_79# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_25/a_696_458#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_55/a_544_485# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_32/a_735_102#
+ prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_29/a_293_74# prbs_generator_syn_1/sky130_fd_sc_hs__nand2_1_17/a_117_74#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_69/a_1034_424# prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_29/a_112_119#
+ prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_37/X prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_31/B
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_19/a_1034_424# prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_33/A
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_9/a_206_368# prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_57/a_376_368#
+ prbs_generator_syn_1/sky130_fd_sc_hs__sdlclkp_2_1/a_706_317# prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_11/B
+ prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_1/a_52_123# prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_39/B
+ prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_21/a_132_392# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_13/a_206_368#
+ prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_43/a_52_123# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_51/a_206_368#
+ prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_47/X prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_23/a_437_503#
+ prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_11/a_52_123# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_61/a_437_503#
+ prbs_generator_syn_1/sky130_fd_sc_hs__nor2b_1_7/Y prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_51/A
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_15/a_696_458# prbs_generator_syn_1/sky130_fd_sc_hs__nor2b_1_5/Y
+ prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_9/a_230_79# prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_25/X
+ prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_19/a_112_119# prbs_generator_syn_1/sky130_fd_sc_hs__nand2_1_45/B
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_5/a_1178_124# prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_19/a_230_79#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_41/a_1226_296# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_59/a_1226_296#
+ prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_63/a_230_79# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_51/Q
+ prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_7/a_132_392# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_9/a_437_503#
+ prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_46/a_376_368# prbs_generator_syn_1/sky130_fd_sc_hs__nand2_1_33/a_117_74#
+ prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_11/a_293_74# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_27/a_1178_124#
+ prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_11/a_132_392# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_13/a_437_503#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_51/a_437_503# prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_5/a_52_123#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_35/a_544_485# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_73/a_651_503#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_45/a_696_458# prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_15/a_52_123#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_47/a_1141_508# prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_47/a_112_119#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_4/a_1178_124# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_17/a_1034_424#
+ prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_23/B prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_37/a_376_368#
+ prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_15/B prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_7/Y
+ prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_29/a_138_385# prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_33/a_230_79#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_25/a_1178_124# prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_47/a_293_74#
+ prbs_generator_syn_1/sky130_fd_sc_hs__nand2_1_37/a_117_74# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_33/a_206_368#
+ prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_15/a_293_74# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_71/a_206_368#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_25/a_544_485# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_67/a_1034_424#
+ prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_13/a_222_392# prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_9/a_52_123#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_15/a_1034_424# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_57/a_1226_296#
+ prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_19/a_52_123# prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_23/X
+ prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_63/a_52_123# prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_19/a_138_385#
+ prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_9/a_376_368# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_21/a_206_368#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_33/a_437_503# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_71/a_437_503#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_53/a_651_503# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_15/a_544_485#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_63/a_696_458# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_65/a_1034_424#
+ prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_19/a_293_74# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_45/a_1141_508#
+ prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_27/a_112_119# prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_67/a_112_119#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_1/a_1178_124# prbs_generator_syn_1/sky130_fd_sc_hs__conb_1_1/a_21_290#
+ prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_63/a_293_74# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_8/a_206_368#
+ prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_17/a_376_368# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_63/a_27_74#
+ prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_21/A prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_55/a_376_368#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_1/a_696_458# prbs_generator_syn_1/sky130_fd_sc_hs__nor2b_1_1/a_278_368#
+ prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_47/a_138_385# prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_33/a_52_123#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_9/a_1034_424# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_21/a_437_503#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_1/a_27_74# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_43/a_651_503#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_1/Q prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_45/a_544_485#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_69/a_735_102# prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_57/a_112_119#
+ prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_31/a_222_392# prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_13/A
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_55/a_1226_296# prbs_generator_syn_1/sky130_fd_sc_hs__nand2_2_5/a_27_74#
+ prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_53/a_230_79# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_8/a_437_503#
+ prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_67/a_293_74# prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_33/a_293_74#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_7/a_735_102# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_23/a_1178_124#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_41/a_206_368# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_8/a_1034_424#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_63/a_1034_424# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_59/a_735_102#
+ prbs_generator_syn_1/sky130_fd_sc_hs__nand2_1_5/B prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_43/a_1141_508#
+ prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_46/a_112_119# prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_61/a_222_392#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_13/a_1034_424# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_73/a_1178_124#
+ prbs_generator_syn_1/sky130_fd_sc_hs__nand2_1_27/B prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_13/B
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_57/a_27_74# prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_57/a_230_79#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_21/a_1178_124# prbs_generator_syn_1/sky130_fd_sc_hs__nor2b_1_1/a_27_112#
+ prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_27/a_138_385# prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_23/a_230_79#
+ prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_67/a_138_385# prbs_generator_syn_1/sky130_fd_sc_hs__nand2_1_41/B
+ prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_9/a_222_392# prbs_generator_syn_1/sky130_fd_sc_hs__nand2_1_27/a_117_74#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_32/a_206_368# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_23/a_651_503#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_41/a_437_503# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_73/a_27_74#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_61/a_651_503# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_63/a_544_485#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_49/a_735_102# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_73/a_696_458#
+ prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_37/a_112_119# prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_51/a_222_392#
+ prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_43/X prbs_generator_syn_1/sky130_fd_sc_hs__nand2_2_1/B
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_9/a_651_503# prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_53/a_52_123#
+ prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_49/X prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_25/a_376_368#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_1/a_544_485# prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_65/a_376_368#
+ prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_57/a_138_385# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_27/a_27_74#
+ prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_39/a_132_392# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_7/a_1034_424#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_13/a_651_503# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_32/a_437_503#
+ prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_27/a_230_79# prbs_generator_syn_1/m3_13600_12265#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_51/a_651_503# prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_59/B
+ prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_47/A prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_61/a_1034_424#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_41/a_1141_508# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_59/a_1141_508#
+ prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_41/a_222_392# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_53/a_1226_296#
+ prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_3/A prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_71/a_1178_124#
+ prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_9/a_112_119# prbs_generator_syn_1/sky130_fd_sc_hs__nand2_1_3/a_117_74#
+ prbs_generator_syn_1/m3_13600_8483# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_39/a_1178_124#
+ prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_57/a_52_123# prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_46/a_138_385#
+ prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_23/a_52_123# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_67/a_27_74#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_53/a_696_458# prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_17/a_112_119#
+ prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_11/A prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_55/a_112_119#
+ prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_1/A prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_51/a_1226_296#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_29/a_1034_424# prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_59/A
+ prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_23/A prbs_generator_syn_1/sky130_fd_sc_hs__nand2_1_39/B
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_5/a_27_74# prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_57/a_293_74#
+ prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_37/a_138_385# prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_59/a_132_392#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_33/a_651_503# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_71/a_651_503#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_43/a_696_458# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_73/a_544_485#
+ prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_27/a_52_123# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_57/a_1141_508#
+ prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_21/a_222_392# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_35/a_27_74#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_69/a_1226_296# prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_37/B
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_19/a_1226_296# prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_35/a_376_368#
+ prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_47/a_230_79# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_37/a_1178_124#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_5/a_1034_424# prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_49/a_132_392#
+ prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_7/a_222_392# prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_27/a_293_74#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_21/a_651_503# prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_9/a_138_385#
+ prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_11/a_222_392# prbs_generator_syn_1/m3_13600_14095#
+ prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_50/A prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_27/a_1034_424#
+ prbs_generator_syn_1/sky130_fd_sc_hs__nand2_1_13/B prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_8/a_651_503#
+ prbs_generator_syn_1/m3_13600_9703# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_35/a_1178_124#
+ prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_17/a_138_385# prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_55/a_138_385#
+ prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_7/a_230_79# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_4/a_1034_424#
+ prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_7/a_376_368# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_69/a_206_368#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_23/a_696_458# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_53/a_544_485#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_39/a_735_102# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_61/a_696_458#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_55/a_1141_508# prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_25/a_112_119#
+ prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_65/a_112_119# prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_43/a_293_74#
+ prbs_generator_syn_1/sky130_fd_sc_hs__nand2_1_57/B prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_25/a_1034_424#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_7/a_206_368# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_17/a_1226_296#
+ prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_15/a_376_368# prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_53/a_376_368#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_9/a_696_458# prbs_generator_syn_1/m3_13600_431#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_45/a_27_74# prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_47/a_52_123#
+ prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_29/a_132_392# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_59/a_206_368#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_69/a_437_503# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_41/a_651_503#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_43/a_544_485# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_13/a_696_458#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_29/a_735_102# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_51/a_696_458#
+ prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_61/Y prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_67/a_1226_296#
+ prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_5/a_132_392# prbs_generator_syn_1/sky130_fd_sc_hs__and2b_2_1/a_198_48#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_7/a_437_503# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_15/a_1226_296#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_69/a_27_74# prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_46/a_293_74#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_1/a_1034_424# prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_19/a_132_392#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_49/a_206_368# prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_7/a_52_123#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_59/a_437_503# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_32/a_651_503#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_7/a_27_74# prbs_generator_syn_1/sky130_fd_sc_hs__nand2_2_1/a_27_74#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_19/a_735_102# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_57/a_735_102#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_65/a_1226_296# prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_37/A
+ prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_33/a_376_368# prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_37/a_230_79#
+ prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_25/a_138_385# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_39/a_27_74#
+ prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_65/a_138_385# prbs_generator_syn_1/sky130_fd_sc_hs__nor2b_1_9/a_278_368#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_49/a_437_503# prbs_generator_syn_1/sky130_fd_sc_hs__and2b_2_1/a_505_74#
+ prbs_generator_syn_1/sky130_fd_sc_hs__nand2_1_51/a_117_74# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_23/a_544_485#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_33/a_696_458# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_61/a_544_485#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_9/a_1226_296# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_53/a_1141_508#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_71/a_696_458# prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_35/a_112_119#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_23/a_1034_424# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_9/a_544_485#
+ prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_63/a_376_368# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_33/a_1178_124#
+ prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_5/a_376_368# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_13/a_544_485#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_73/a_1034_424# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_21/a_696_458#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_51/a_544_485# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_8/a_1226_296#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_51/a_1141_508# prbs_generator_syn_1/sky130_fd_sc_hs__nand2_1_55/a_117_74#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_21/a_1034_424# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_63/a_1226_296#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_23/a_27_74# prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_7/a_112_119#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_13/a_1226_296# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_8/a_696_458#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_32/a_1178_124# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_49/a_1178_124#
+ prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_37/a_52_123# prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_27/a_132_392#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_71/Q prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_67/a_735_102#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_69/a_1141_508# prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_15/a_112_119#
+ prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_53/a_112_119# prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_39/a_222_392#
+ prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_55/a_230_79# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_19/a_1141_508#
+ prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_37/a_293_74# prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_43/a_376_368#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_5/a_735_102# prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_35/a_138_385#
+ prbs_generator_syn_1/sky130_fd_sc_hs__sdlclkp_2_1/a_114_424# prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_57/a_132_392#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_71/a_1034_424# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_7/a_1226_296#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_33/a_544_485# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_41/a_696_458#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_71/a_544_485# prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_21/B
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_61/a_1226_296# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_39/a_1034_424#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_17/a_27_74# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_9/a_27_74#
+ prbs_generator_syn_1/sky130_fd_sc_hs__nor2b_1_5/a_27_112# prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_47/a_132_392#
+ prbs_generator_syn_1/sky130_fd_sc_hs__nor2b_1_8/a_278_368# prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_9/B
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_39/a_206_368# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_33/a_27_74#
+ prbs_generator_syn_1/sky130_fd_sc_hs__nand2_1_41/a_117_74# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_69/a_651_503#
+ prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_51/a_293_74# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_21/a_544_485#
+ prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_7/a_138_385# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_32/a_696_458#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_47/a_735_102# prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_33/a_112_119#
+ prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_59/a_222_392# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_17/a_1141_508#
+ prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_55/a_52_123# prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_3/a_293_74#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_7/a_651_503# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_29/a_1226_296#
+ prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_23/a_376_368# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_8/a_544_485#
+ prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_47/B prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_47/a_1178_124#
+ prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_15/a_138_385# prbs_generator_syn_1/sky130_fd_sc_hs__sdlclkp_2_1/a_1195_374#
+ prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_53/a_138_385# prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_37/a_132_392#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_29/a_206_368# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_39/a_437_503#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_59/a_651_503# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_37/a_735_102#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_67/a_1141_508# prbs_generator_syn_1/sky130_fd_sc_hs__and2b_2_1/a_27_74#
+ prbs_generator_syn_1/sky130_fd_sc_hs__conb_1_1/a_165_290# prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_55/a_293_74#
+ prbs_generator_syn_1/sky130_fd_sc_hs__nand2_1_45/a_117_74# prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_63/a_112_119#
+ prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_49/a_222_392# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_37/a_1034_424#
+ prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_23/a_293_74# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_15/a_1141_508#
+ prbs_generator_syn_1/sky130_fd_sc_hs__nand2_1_5/a_117_74# prbs_generator_syn_1/m3_13600_13485#
+ prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_5/a_112_119# prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_13/a_376_368#
+ prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_51/a_376_368# prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_7/a_293_74#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_19/a_206_368# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_57/a_206_368#
+ prbs_generator_syn_1/sky130_fd_sc_hs__sdlclkp_2_1/a_318_74# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_29/a_437_503#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_49/a_651_503# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_25/a_27_74#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_5/a_1226_296# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_41/a_544_485#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_27/a_735_102# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_65/a_1141_508#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_65/a_735_102# prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_3/a_230_79#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_35/a_1034_424# prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_13/a_230_79#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_41/a_27_74# prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_3/a_132_392#
+ prbs_generator_syn_1/sky130_fd_sc_hs__nand2_1_49/a_117_74# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_27/a_1226_296#
+ prbs_generator_syn_1/sky130_fd_sc_hs__nand2_1_15/a_117_74# prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_41/a_376_368#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_45/a_1178_124# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_4/a_735_102#
+ prbs_generator_syn_1/sky130_fd_sc_hs__nand2_1_9/a_117_74# prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_33/a_138_385#
+ prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_17/a_132_392# prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_55/a_132_392#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_9/a_1141_508# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_19/a_437_503#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_57/a_437_503# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_4/a_1226_296#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_32/a_544_485# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_17/a_735_102#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_55/a_735_102# prbs_generator_syn_1/m3_13600_2261#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_65/a_27_74# prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_29/a_222_392#
+ prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_43/a_112_119# prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_19/X
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_25/a_1226_296# prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_31/a_376_368#
+ prbs_generator_syn_1/sky130_fd_sc_hs__or2_1_1/a_63_368# prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_17/a_230_79#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_4/a_27_74# prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_61/a_230_79#
+ prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_63/a_138_385# prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_5/a_222_392#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_8/a_1141_508# prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_41/a_293_74#
+ prbs_generator_syn_1/sky130_fd_sc_hs__nand2_1_31/a_117_74# prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_5/a_138_385#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_63/a_1141_508# prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_19/a_222_392#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_13/a_1141_508# prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_3/a_52_123#
+ prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_13/a_52_123# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_43/a_1178_124#
+ prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_61/a_376_368# prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_35/a_132_392#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_67/a_206_368# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_1/a_1226_296#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_69/a_696_458# prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_31/a_230_79#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_35/a_735_102# prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_23/a_112_119#
+ prbs_generator_syn_1/sky130_fd_sc_hs__nand2_1_35/a_117_74# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_59/a_27_74#
+ prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_13/a_293_74# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_5/a_206_368#
+ prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_50/a_376_368# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_7/a_696_458#
+ prbs_generator_syn_1/sky130_fd_sc_hs__nor2b_1_7/a_278_368# prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_17/a_52_123#
+ prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_43/a_138_385# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_7/a_1141_508#
+ prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_61/a_52_123# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_67/a_437_503#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_61/a_1141_508# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_25/a_735_102#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_59/a_696_458# prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_13/a_112_119#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_33/a_1034_424# prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_51/a_112_119#
+ prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_35/a_230_79# prbs_generator_syn_1/m3_13600_4091#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_23/a_1226_296# prbs_generator_syn_1/sky130_fd_sc_hs__nand2_1_39/a_117_74#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_29/a_27_74# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_5/a_437_503#
+ prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_17/a_293_74# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_41/a_1178_124#
+ prbs_generator_syn_1/sky130_fd_sc_hs__or2_1_1/a_152_368# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_59/a_1178_124#
+ prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_61/a_293_74# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_47/a_206_368#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_39/a_651_503# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_49/a_696_458#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_15/a_735_102# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_32/a_1034_424#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_73/a_1226_296# prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_27/a_222_392#
+ prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_41/a_112_119# prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_31/a_52_123#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_49/a_1034_424# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_29/a_1141_508#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_21/a_1226_296# prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_39/a_230_79#
+ prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_23/a_138_385# prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_51/a_230_79#
+ prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_45/a_132_392# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_37/a_206_368#
+ prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_65/a_293_74# prbs_generator_syn_1/sky130_fd_sc_hs__nand2_1_53/a_117_74#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_47/a_437_503# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_29/a_651_503#
+ prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_31/a_293_74# prbs_generator_syn_1/sky130_fd_sc_hs__nand2_1_21/a_117_74#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_69/a_544_485# prbs_generator_syn_1/sky130_fd_sc_hs__clkbuf_16_1/a_114_74#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_45/a_735_102# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_13/a_27_74#
+ prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_31/a_112_119# prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_57/a_222_392#
+ prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_35/a_52_123# prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_21/a_376_368#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_7/a_544_485# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_57/a_1178_124#
+ prbs_generator_syn_1/m3_13600_6043# prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_13/a_138_385#
+ prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_51/a_138_385# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_5/a_1141_508#
+ prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_3/a_376_368# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_27/a_206_368#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_65/a_206_368# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_37/a_437_503#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_19/a_651_503# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_57/a_651_503#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_59/a_544_485# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_71/a_1226_296#
+ prbs_generator_syn_1/sky130_fd_sc_hs__nand2_1_25/a_117_74# prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_61/a_112_119#
+ prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_47/a_222_392# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_27/a_1141_508#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_53/a_27_74# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_4/a_206_368#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_39/a_1226_296# prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_11/a_376_368#
+ prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_39/a_52_123# prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_41/a_138_385#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_4/a_1141_508# prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_25/a_132_392#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_17/a_206_368# prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_41/A
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_55/a_206_368# prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_51/a_52_123#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_27/a_437_503# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_65/a_437_503#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_49/a_544_485# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_63/a_735_102#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_47/a_1034_424# prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_50/a_112_119#
+ prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_37/a_222_392# prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_59/a_230_79#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_25/a_1141_508# prbs_generator_syn_1/sky130_fd_sc_hs__nor2b_1_4/a_27_112#
+ prbs_generator_syn_1/sky130_fd_sc_hs__sdlclkp_2_1/a_685_81# prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_1/a_132_392#
+ prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_39/a_293_74# prbs_generator_syn_1/sky130_fd_sc_hs__nand2_1_29/a_117_74#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_4/a_437_503# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_55/a_1178_124#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_21/a_27_74# prbs_generator_syn_1/m3_13600_12875#
+ prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_50/a_293_74# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_1/a_735_102#
+ prbs_generator_syn_1/sky130_fd_sc_hs__xnor2_1_31/a_138_385# prbs_generator_syn_1/sky130_fd_sc_hs__a22o_1_15/a_132_392#
+ prbs_generator_syn_1/sky130_fd_sc_hs__nand2_1_1/a_117_74# prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_17/a_437_503#
+ prbs_generator_syn_1/sky130_fd_sc_hs__dfxtp_4_55/a_437_503# prbs_generator_syn
Xsky130_fd_sc_hs__clkdlyinv5sd2_1_0 DVSS: DVDD: DVSS: DVDD: dout_p sky130_fd_sc_hs__nand2_2_1/B
+ sky130_fd_sc_hs__clkdlyinv5sd2_1_1/a_28_74# sky130_fd_sc_hs__clkdlyinv5sd2_1_1/a_682_74#
+ sky130_fd_sc_hs__clkdlyinv5sd2_1_1/a_549_74# sky130_fd_sc_hs__clkdlyinv5sd2_1_1/a_288_74#
+ sky130_fd_sc_hs__clkdlyinv5sd2_1
Xsky130_fd_sc_hs__o21bai_2_8 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__nand2_2_7/A
+ sky130_fd_sc_hs__o21bai_4_7/A1 sky130_fd_sc_hs__dlrtp_1_65/D sky130_fd_sc_hs__buf_2_57/A
+ sky130_fd_sc_hs__o21bai_2_9/a_27_74# sky130_fd_sc_hs__o21bai_2_9/a_225_74# sky130_fd_sc_hs__o21bai_2_9/a_507_368#
+ sky130_fd_sc_hs__o21bai_2
Xsky130_fd_sc_hs__o21ai_2_13 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__inv_4_13/Y sky130_fd_sc_hs__nand2_2_9/B
+ sky130_fd_sc_hs__o21ai_2_55/A1 sky130_fd_sc_hs__buf_2_47/A sky130_fd_sc_hs__o21ai_2_13/a_116_368#
+ sky130_fd_sc_hs__o21ai_2_13/a_27_74# sky130_fd_sc_hs__o21ai_2
Xsky130_fd_sc_hs__o21ai_2_24 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__inv_4_15/Y sky130_fd_sc_hs__nand2_2_11/B
+ sky130_fd_sc_hs__o21ai_2_55/A1 sky130_fd_sc_hs__o21ai_2_25/Y sky130_fd_sc_hs__o21ai_2_25/a_116_368#
+ sky130_fd_sc_hs__o21ai_2_25/a_27_74# sky130_fd_sc_hs__o21ai_2
Xsky130_fd_sc_hs__o21ai_2_35 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__inv_4_21/Y sky130_fd_sc_hs__buf_8_3/X
+ sky130_fd_sc_hs__clkinv_4_7/Y sky130_fd_sc_hs__buf_2_91/A sky130_fd_sc_hs__o21ai_2_35/a_116_368#
+ sky130_fd_sc_hs__o21ai_2_35/a_27_74# sky130_fd_sc_hs__o21ai_2
Xsky130_fd_sc_hs__o21ai_2_46 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__nand2_2_27/B
+ sky130_fd_sc_hs__nand2_2_21/B sky130_fd_sc_hs__clkinv_4_7/Y sky130_fd_sc_hs__o21ai_2_47/Y
+ sky130_fd_sc_hs__o21ai_2_47/a_116_368# sky130_fd_sc_hs__o21ai_2_47/a_27_74# sky130_fd_sc_hs__o21ai_2
Xsky130_fd_sc_hs__o21ai_2_57 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__inv_4_29/A sky130_fd_sc_hs__o21ai_2_3/A2
+ sky130_fd_sc_hs__or2b_4_3/X sky130_fd_sc_hs__buf_2_157/A sky130_fd_sc_hs__o21ai_2_57/a_116_368#
+ sky130_fd_sc_hs__o21ai_2_57/a_27_74# sky130_fd_sc_hs__o21ai_2
Xsky130_fd_sc_hs__clkinv_4_16 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__nor2_4_3/B
+ sky130_fd_sc_hs__nand2_2_7/A sky130_fd_sc_hs__clkinv_4
Xprbs_generator_syn_18 prbs_generator_syn_19/clk prbs_generator_syn_19/rst prbs_generator_syn_19/cke
+ sky130_fd_sc_hs__conb_1_209/LO sky130_fd_sc_hs__conb_1_209/LO sky130_fd_sc_hs__conb_1_209/HI
+ sky130_fd_sc_hs__conb_1_209/HI sky130_fd_sc_hs__conb_1_209/LO sky130_fd_sc_hs__conb_1_209/LO
+ sky130_fd_sc_hs__conb_1_209/LO sky130_fd_sc_hs__conb_1_209/HI sky130_fd_sc_hs__conb_1_209/HI
+ sky130_fd_sc_hs__conb_1_209/HI sky130_fd_sc_hs__conb_1_209/HI prbs_generator_syn_19/cke
+ prbs_generator_syn_19/eqn[31] prbs_generator_syn_19/cke prbs_generator_syn_19/eqn[31]
+ prbs_generator_syn_19/eqn[31] prbs_generator_syn_19/eqn[31] prbs_generator_syn_19/eqn[31]
+ prbs_generator_syn_19/eqn[2] prbs_generator_syn_19/eqn[2] prbs_generator_syn_19/eqn[2]
+ prbs_generator_syn_19/eqn[2] prbs_generator_syn_19/eqn[2] prbs_generator_syn_19/eqn[1]
+ sky130_fd_sc_hs__conb_1_203/HI sky130_fd_sc_hs__conb_1_203/HI sky130_fd_sc_hs__conb_1_203/HI
+ sky130_fd_sc_hs__conb_1_203/HI sky130_fd_sc_hs__conb_1_203/LO sky130_fd_sc_hs__conb_1_203/LO
+ sky130_fd_sc_hs__conb_1_203/HI sky130_fd_sc_hs__conb_1_203/HI prbs_generator_syn_19/eqn[31]
+ prbs_generator_syn_19/eqn[30] prbs_generator_syn_19/eqn[30] prbs_generator_syn_19/eqn[30]
+ prbs_generator_syn_19/eqn[30] prbs_generator_syn_19/eqn[30] prbs_generator_syn_19/eqn[30]
+ prbs_generator_syn_19/eqn[30] prbs_generator_syn_19/eqn[30] prbs_generator_syn_19/eqn[22]
+ prbs_generator_syn_19/eqn[22] prbs_generator_syn_19/eqn[20] prbs_generator_syn_19/eqn[22]
+ prbs_generator_syn_19/eqn[22] prbs_generator_syn_19/eqn[22] prbs_generator_syn_19/eqn[22]
+ prbs_generator_syn_19/eqn[22] prbs_generator_syn_19/eqn[22] prbs_generator_syn_19/eqn[13]
+ prbs_generator_syn_19/eqn[13] prbs_generator_syn_19/eqn[13] prbs_generator_syn_19/eqn[9]
+ prbs_generator_syn_19/eqn[9] prbs_generator_syn_19/eqn[9] prbs_generator_syn_19/eqn[9]
+ prbs_generator_syn_19/eqn[9] prbs_generator_syn_19/eqn[9] prbs_generator_syn_19/eqn[9]
+ prbs_generator_syn_19/eqn[9] prbs_generator_syn_19/eqn[2] prbs_generator_syn_19/eqn[1]
+ prbs_generator_syn_19/eqn[2] prbs_generator_syn_19/inj_err prbs_generator_syn_19/eqn[31]
+ prbs_generator_syn_19/eqn[31] prbs_generator_syn_19/out DVSS: DVDD: prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_1/a_293_74#
+ prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_15/X prbs_generator_syn_19/sky130_fd_sc_hs__nand2_1_35/B
+ prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_51/Y prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_9/A
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_9/CLK prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_47/a_27_74#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_37/a_1226_296# prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_3/B
+ prbs_generator_syn_19/sky130_fd_sc_hs__nor2b_1_7/a_27_112# prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_29/B
+ prbs_generator_syn_19/sky130_fd_sc_hs__sdlclkp_2_1/a_580_74# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_1/a_1141_508#
+ prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_5/Y prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_41/a_230_79#
+ prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_61/a_138_385# prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_43/a_132_392#
+ prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_3/a_222_392# prbs_generator_syn_19/sky130_fd_sc_hs__nor2b_1_9/a_27_112#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_61/a_27_74# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_35/a_206_368#
+ prbs_generator_syn_19/sky130_fd_sc_hs__nand2_2_3/Y prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_25/B
+ prbs_generator_syn_19/sky130_fd_sc_hs__nand2_1_11/a_117_74# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_67/a_651_503#
+ prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_45/X prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_39/a_696_458#
+ prbs_generator_syn_19/sky130_fd_sc_hs__sdlclkp_2_1/a_1198_74# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_45/a_1034_424#
+ prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_17/a_222_392# prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_55/a_222_392#
+ prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_53/Y prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_35/A
+ prbs_generator_syn_19/m3_13600_1651# prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_59/a_52_123#
+ prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_5/a_293_74# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_35/a_1226_296#
+ prbs_generator_syn_19/sky130_fd_sc_hs__nand2_1_51/B prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_5/a_651_503#
+ prbs_generator_syn_19/sky130_fd_sc_hs__nand2_1_21/B prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_8/a_27_74#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_15/a_27_74# prbs_generator_syn_19/sky130_fd_sc_hs__and2b_2_1/X
+ prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_13/X prbs_generator_syn_19/sky130_fd_sc_hs__nand2_2_3/a_27_74#
+ prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_50/a_138_385# prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_33/a_132_392#
+ prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_1/a_376_368# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_25/a_206_368#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_35/a_437_503# prbs_generator_syn_19/sky130_fd_sc_hs__sdlclkp_2_1/a_708_451#
+ prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_45/a_230_79# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_29/a_696_458#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_32/a_27_74# prbs_generator_syn_19/sky130_fd_sc_hs__nor2b_1_4/Y
+ prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_59/a_293_74# prbs_generator_syn_19/sky130_fd_sc_hs__nand2_1_47/a_117_74#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_73/a_735_102# prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_21/a_112_119#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_23/a_1141_508# prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_25/a_293_74#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_7/Q prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_3/a_112_119#
+ prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_35/B prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_51/X
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_53/a_1178_124# prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_23/a_132_392#
+ prbs_generator_syn_19/sky130_fd_sc_hs__nand2_1_3/B prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_15/a_206_368#
+ prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_63/a_132_392# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_55/a_27_74#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_25/a_437_503# prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_41/a_52_123#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_47/a_651_503# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_73/a_1141_508#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_19/a_696_458# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_57/a_696_458#
+ prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_7/X prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_43/a_1034_424#
+ prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_55/A prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_11/a_112_119#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_21/a_1141_508# prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_35/a_222_392#
+ prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_49/a_230_79# prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_67/Y
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_71/a_27_74# prbs_generator_syn_19/sky130_fd_sc_hs__nand2_1_33/B
+ prbs_generator_syn_19/sky130_fd_sc_hs__conb_1_1/LO prbs_generator_syn_19/sky130_fd_sc_hs__nand2_1_19/a_117_74#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_51/a_1178_124# prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_33/X
+ prbs_generator_syn_19/sky130_fd_sc_hs__nand2_1_29/B prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_41/Y
+ prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_53/a_132_392# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_45/a_206_368#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_15/a_437_503# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_37/a_651_503#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_39/a_544_485# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_53/a_735_102#
+ prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_45/a_52_123# prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_1/B
+ prbs_generator_syn_19/sky130_fd_sc_hs__nand2_2_3/B prbs_generator_syn_19/sky130_fd_sc_hs__clkbuf_16_1/A
+ prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_21/X prbs_generator_syn_19/sky130_fd_sc_hs__nand2_1_25/B
+ prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_39/a_376_368# prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_63/X
+ prbs_generator_syn_19/m3_13600_3481# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_69/a_1178_124#
+ prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_21/a_138_385# prbs_generator_syn_19/sky130_fd_sc_hs__nor2b_1_8/Y
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_19/a_1178_124# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_49/a_27_74#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_45/a_437_503# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_27/a_651_503#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_71/a_1141_508# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_65/a_651_503#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_29/a_544_485# prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_3/a_138_385#
+ prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_55/X prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_43/a_735_102#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_41/a_1034_424# prbs_generator_syn_19/sky130_fd_sc_hs__nand2_1_9/B
+ prbs_generator_syn_19/sky130_fd_sc_hs__nor2b_1_9/Y prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_59/a_1034_424#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_39/a_1141_508# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_33/a_1226_296#
+ prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_49/a_52_123# prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_47/Y
+ prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_43/Y prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_4/a_651_503#
+ prbs_generator_syn_19/sky130_fd_sc_hs__nand2_1_49/B prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_19/A
+ prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_11/a_138_385# prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_5/X
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_63/a_206_368# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_17/a_651_503#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_19/a_544_485# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_55/a_651_503#
+ prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_9/Y prbs_generator_syn_19/sky130_fd_sc_hs__nand2_1_17/B
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_57/a_544_485# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_67/a_696_458#
+ prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_35/X prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_19/a_27_74#
+ prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_45/a_222_392# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_32/a_1226_296#
+ prbs_generator_syn_19/sky130_fd_sc_hs__nand2_1_43/B prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_25/A
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_1/a_206_368# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_49/a_1226_296#
+ prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_1/a_112_119# prbs_generator_syn_19/sky130_fd_sc_hs__or2_1_1/X
+ prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_59/a_376_368# prbs_generator_syn_19/sky130_fd_sc_hs__nand2_1_19/B
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_5/a_696_458# prbs_generator_syn_19/sky130_fd_sc_hs__nor2b_1_1/Y
+ prbs_generator_syn_19/sky130_fd_sc_hs__nor2b_1_5/a_278_368# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_17/a_1178_124#
+ prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_39/X prbs_generator_syn_19/m3_13600_5433#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_63/a_437_503# prbs_generator_syn_19/sky130_fd_sc_hs__nand2_2_5/B
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_23/a_735_102# prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_53/A
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_61/a_735_102# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_57/a_1034_424#
+ prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_63/B prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_37/a_1141_508#
+ prbs_generator_syn_19/sky130_fd_sc_hs__nand2_1_47/B prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_29/X
+ prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_65/Y prbs_generator_syn_19/m3_13600_4701#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_1/a_437_503# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_67/a_1178_124#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_9/a_735_102# prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_13/a_132_392#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_15/a_1178_124# prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_15/A
+ prbs_generator_syn_19/sky130_fd_sc_hs__nand2_1_1/B prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_43/B
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_35/a_651_503# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_8/D
+ prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_29/A prbs_generator_syn_19/sky130_fd_sc_hs__nand2_1_7/B
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_13/a_735_102# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_47/a_696_458#
+ prbs_generator_syn_19/sky130_fd_sc_hs__nand2_1_31/B prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_51/a_735_102#
+ prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_59/X prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_35/a_1141_508#
+ prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_25/a_222_392# prbs_generator_syn_19/sky130_fd_sc_hs__sdlclkp_2_1/a_288_48#
+ prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_55/B prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_17/B
+ prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_43/A prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_7/A
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_65/a_1178_124# prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_59/Y
+ prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_41/X prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_21/a_230_79#
+ prbs_generator_syn_19/sky130_fd_sc_hs__nand2_1_57/a_117_74# prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_1/a_222_392#
+ prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_19/B prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_35/a_293_74#
+ prbs_generator_syn_19/sky130_fd_sc_hs__nand2_1_23/a_117_74# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_73/a_206_368#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_25/a_651_503# prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_1/a_138_385#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_37/a_696_458# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_67/a_544_485#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_43/a_27_74# prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_9/X
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_55/a_1034_424# prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_39/a_112_119#
+ prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_15/a_222_392# prbs_generator_syn_19/sky130_fd_sc_hs__conb_1_1/HI
+ prbs_generator_syn_19/sky130_fd_sc_hs__nand2_1_23/B prbs_generator_syn_19/sky130_fd_sc_hs__nand2_1_53/B
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_9/a_1178_124# prbs_generator_syn_19/sky130_fd_sc_hs__nor2b_1_4/A
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_47/a_1226_296# prbs_generator_syn_19/m3_13600_11045#
+ prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_17/X prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_29/a_376_368#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_5/a_544_485# prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_3/X
+ prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_31/a_132_392# prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_61/A
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_15/a_651_503# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_73/a_437_503#
+ prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_25/a_230_79# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_27/a_696_458#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_65/a_696_458# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_33/a_735_102#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_71/a_735_102# prbs_generator_syn_19/m3_13600_7263#
+ prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_43/a_222_392# prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_50/Y
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_8/a_1178_124# prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_53/B
+ prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_19/a_376_368# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_63/a_1178_124#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_4/a_696_458# prbs_generator_syn_19/sky130_fd_sc_hs__nor2b_1_4/a_278_368#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_13/a_1178_124# prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_61/a_132_392#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_53/a_206_368# prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_21/a_52_123#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_45/a_651_503# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_17/a_696_458#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_47/a_544_485# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_55/a_696_458#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_21/a_735_102# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_37/a_27_74#
+ prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_61/B prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_61/X
+ prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_59/a_112_119# prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_31/A
+ prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_33/a_222_392# prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_29/a_230_79#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_45/a_1226_296# prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_9/a_132_392#
+ prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_5/A prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_57/Y
+ prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_31/X prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_51/a_27_74#
+ prbs_generator_syn_19/sky130_fd_sc_hs__nor2b_1_8/a_27_112# prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_47/a_376_368#
+ prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_53/a_293_74# prbs_generator_syn_19/sky130_fd_sc_hs__nand2_1_43/a_117_74#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_8/a_735_102# prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_21/a_293_74#
+ prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_39/a_138_385# prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_63/Y
+ prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_51/a_132_392# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_43/a_206_368#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_53/a_437_503# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_37/a_544_485#
+ prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_57/X prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_53/a_1034_424#
+ prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_25/a_52_123# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_33/a_1141_508#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_63/Q prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_23/a_222_392#
+ prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_63/a_222_392# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_7/a_1178_124#
+ prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_53/X prbs_generator_syn_19/sky130_fd_sc_hs__nand2_2_5/Y
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_61/a_1178_124# prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_1/a_230_79#
+ prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_43/a_230_79# prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_11/a_230_79#
+ prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_41/a_132_392# prbs_generator_syn_19/sky130_fd_sc_hs__nand2_1_13/a_117_74#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_43/a_437_503# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_27/a_544_485#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_63/a_651_503# prbs_generator_syn_19/sky130_fd_sc_hs__nand2_1_7/a_117_74#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_35/a_696_458# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_65/a_544_485#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_51/a_1034_424# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_41/a_735_102#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_32/a_1141_508# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_49/a_1141_508#
+ prbs_generator_syn_19/sky130_fd_sc_hs__nand2_1_55/B prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_53/a_222_392#
+ prbs_generator_syn_19/sky130_fd_sc_hs__sdlclkp_2_1/a_114_112# prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_9/a_293_74#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_43/a_1226_296# prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_29/a_52_123#
+ prbs_generator_syn_19/sky130_fd_sc_hs__nand2_1_37/B prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_1/a_651_503#
+ prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_27/a_376_368# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_4/a_544_485#
+ prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_67/a_376_368# prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_27/X
+ prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_1/X prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_59/a_138_385#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_29/a_1178_124# prbs_generator_syn_19/m3_13600_2871#
+ prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_5/a_230_79# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_23/a_206_368#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_61/a_206_368# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_17/a_544_485#
+ prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_15/a_230_79# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_25/a_696_458#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_55/a_544_485# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_32/a_735_102#
+ prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_29/a_293_74# prbs_generator_syn_19/sky130_fd_sc_hs__nand2_1_17/a_117_74#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_69/a_1034_424# prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_29/a_112_119#
+ prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_37/X prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_31/B
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_19/a_1034_424# prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_33/A
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_9/a_206_368# prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_57/a_376_368#
+ prbs_generator_syn_19/sky130_fd_sc_hs__sdlclkp_2_1/a_706_317# prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_11/B
+ prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_1/a_52_123# prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_39/B
+ prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_21/a_132_392# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_13/a_206_368#
+ prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_43/a_52_123# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_51/a_206_368#
+ prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_47/X prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_23/a_437_503#
+ prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_11/a_52_123# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_61/a_437_503#
+ prbs_generator_syn_19/sky130_fd_sc_hs__nor2b_1_7/Y prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_51/A
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_15/a_696_458# prbs_generator_syn_19/sky130_fd_sc_hs__nor2b_1_5/Y
+ prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_9/a_230_79# prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_25/X
+ prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_19/a_112_119# prbs_generator_syn_19/sky130_fd_sc_hs__nand2_1_45/B
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_5/a_1178_124# prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_19/a_230_79#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_41/a_1226_296# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_59/a_1226_296#
+ prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_63/a_230_79# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_51/Q
+ prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_7/a_132_392# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_9/a_437_503#
+ prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_46/a_376_368# prbs_generator_syn_19/sky130_fd_sc_hs__nand2_1_33/a_117_74#
+ prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_11/a_293_74# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_27/a_1178_124#
+ prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_11/a_132_392# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_13/a_437_503#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_51/a_437_503# prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_5/a_52_123#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_35/a_544_485# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_73/a_651_503#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_45/a_696_458# prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_15/a_52_123#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_47/a_1141_508# prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_47/a_112_119#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_4/a_1178_124# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_17/a_1034_424#
+ prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_23/B prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_37/a_376_368#
+ prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_15/B prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_7/Y
+ prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_29/a_138_385# prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_33/a_230_79#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_25/a_1178_124# prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_47/a_293_74#
+ prbs_generator_syn_19/sky130_fd_sc_hs__nand2_1_37/a_117_74# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_33/a_206_368#
+ prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_15/a_293_74# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_71/a_206_368#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_25/a_544_485# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_67/a_1034_424#
+ prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_13/a_222_392# prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_9/a_52_123#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_15/a_1034_424# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_57/a_1226_296#
+ prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_19/a_52_123# prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_23/X
+ prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_63/a_52_123# prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_19/a_138_385#
+ prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_9/a_376_368# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_21/a_206_368#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_33/a_437_503# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_71/a_437_503#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_53/a_651_503# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_15/a_544_485#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_63/a_696_458# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_65/a_1034_424#
+ prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_19/a_293_74# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_45/a_1141_508#
+ prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_27/a_112_119# prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_67/a_112_119#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_1/a_1178_124# prbs_generator_syn_19/sky130_fd_sc_hs__conb_1_1/a_21_290#
+ prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_63/a_293_74# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_8/a_206_368#
+ prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_17/a_376_368# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_63/a_27_74#
+ prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_21/A prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_55/a_376_368#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_1/a_696_458# prbs_generator_syn_19/sky130_fd_sc_hs__nor2b_1_1/a_278_368#
+ prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_47/a_138_385# prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_33/a_52_123#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_9/a_1034_424# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_21/a_437_503#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_1/a_27_74# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_43/a_651_503#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_1/Q prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_45/a_544_485#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_69/a_735_102# prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_57/a_112_119#
+ prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_31/a_222_392# prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_13/A
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_55/a_1226_296# prbs_generator_syn_19/sky130_fd_sc_hs__nand2_2_5/a_27_74#
+ prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_53/a_230_79# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_8/a_437_503#
+ prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_67/a_293_74# prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_33/a_293_74#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_7/a_735_102# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_23/a_1178_124#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_41/a_206_368# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_8/a_1034_424#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_63/a_1034_424# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_59/a_735_102#
+ prbs_generator_syn_19/sky130_fd_sc_hs__nand2_1_5/B prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_43/a_1141_508#
+ prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_46/a_112_119# prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_61/a_222_392#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_13/a_1034_424# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_73/a_1178_124#
+ prbs_generator_syn_19/sky130_fd_sc_hs__nand2_1_27/B prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_13/B
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_57/a_27_74# prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_57/a_230_79#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_21/a_1178_124# prbs_generator_syn_19/sky130_fd_sc_hs__nor2b_1_1/a_27_112#
+ prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_27/a_138_385# prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_23/a_230_79#
+ prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_67/a_138_385# prbs_generator_syn_19/sky130_fd_sc_hs__nand2_1_41/B
+ prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_9/a_222_392# prbs_generator_syn_19/sky130_fd_sc_hs__nand2_1_27/a_117_74#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_32/a_206_368# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_23/a_651_503#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_41/a_437_503# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_73/a_27_74#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_61/a_651_503# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_63/a_544_485#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_49/a_735_102# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_73/a_696_458#
+ prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_37/a_112_119# prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_51/a_222_392#
+ prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_43/X prbs_generator_syn_19/sky130_fd_sc_hs__nand2_2_1/B
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_9/a_651_503# prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_53/a_52_123#
+ prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_49/X prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_25/a_376_368#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_1/a_544_485# prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_65/a_376_368#
+ prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_57/a_138_385# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_27/a_27_74#
+ prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_39/a_132_392# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_7/a_1034_424#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_13/a_651_503# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_32/a_437_503#
+ prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_27/a_230_79# prbs_generator_syn_19/m3_13600_12265#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_51/a_651_503# prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_59/B
+ prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_47/A prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_61/a_1034_424#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_41/a_1141_508# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_59/a_1141_508#
+ prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_41/a_222_392# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_53/a_1226_296#
+ prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_3/A prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_71/a_1178_124#
+ prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_9/a_112_119# prbs_generator_syn_19/sky130_fd_sc_hs__nand2_1_3/a_117_74#
+ prbs_generator_syn_19/m3_13600_8483# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_39/a_1178_124#
+ prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_57/a_52_123# prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_46/a_138_385#
+ prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_23/a_52_123# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_67/a_27_74#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_53/a_696_458# prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_17/a_112_119#
+ prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_11/A prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_55/a_112_119#
+ prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_1/A prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_51/a_1226_296#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_29/a_1034_424# prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_59/A
+ prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_23/A prbs_generator_syn_19/sky130_fd_sc_hs__nand2_1_39/B
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_5/a_27_74# prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_57/a_293_74#
+ prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_37/a_138_385# prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_59/a_132_392#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_33/a_651_503# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_71/a_651_503#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_43/a_696_458# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_73/a_544_485#
+ prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_27/a_52_123# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_57/a_1141_508#
+ prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_21/a_222_392# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_35/a_27_74#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_69/a_1226_296# prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_37/B
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_19/a_1226_296# prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_35/a_376_368#
+ prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_47/a_230_79# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_37/a_1178_124#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_5/a_1034_424# prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_49/a_132_392#
+ prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_7/a_222_392# prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_27/a_293_74#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_21/a_651_503# prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_9/a_138_385#
+ prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_11/a_222_392# prbs_generator_syn_19/m3_13600_14095#
+ prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_50/A prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_27/a_1034_424#
+ prbs_generator_syn_19/sky130_fd_sc_hs__nand2_1_13/B prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_8/a_651_503#
+ prbs_generator_syn_19/m3_13600_9703# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_35/a_1178_124#
+ prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_17/a_138_385# prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_55/a_138_385#
+ prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_7/a_230_79# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_4/a_1034_424#
+ prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_7/a_376_368# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_69/a_206_368#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_23/a_696_458# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_53/a_544_485#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_39/a_735_102# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_61/a_696_458#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_55/a_1141_508# prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_25/a_112_119#
+ prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_65/a_112_119# prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_43/a_293_74#
+ prbs_generator_syn_19/sky130_fd_sc_hs__nand2_1_57/B prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_25/a_1034_424#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_7/a_206_368# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_17/a_1226_296#
+ prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_15/a_376_368# prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_53/a_376_368#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_9/a_696_458# prbs_generator_syn_19/m3_13600_431#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_45/a_27_74# prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_47/a_52_123#
+ prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_29/a_132_392# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_59/a_206_368#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_69/a_437_503# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_41/a_651_503#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_43/a_544_485# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_13/a_696_458#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_29/a_735_102# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_51/a_696_458#
+ prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_61/Y prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_67/a_1226_296#
+ prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_5/a_132_392# prbs_generator_syn_19/sky130_fd_sc_hs__and2b_2_1/a_198_48#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_7/a_437_503# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_15/a_1226_296#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_69/a_27_74# prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_46/a_293_74#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_1/a_1034_424# prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_19/a_132_392#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_49/a_206_368# prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_7/a_52_123#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_59/a_437_503# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_32/a_651_503#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_7/a_27_74# prbs_generator_syn_19/sky130_fd_sc_hs__nand2_2_1/a_27_74#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_19/a_735_102# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_57/a_735_102#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_65/a_1226_296# prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_37/A
+ prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_33/a_376_368# prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_37/a_230_79#
+ prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_25/a_138_385# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_39/a_27_74#
+ prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_65/a_138_385# prbs_generator_syn_19/sky130_fd_sc_hs__nor2b_1_9/a_278_368#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_49/a_437_503# prbs_generator_syn_19/sky130_fd_sc_hs__and2b_2_1/a_505_74#
+ prbs_generator_syn_19/sky130_fd_sc_hs__nand2_1_51/a_117_74# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_23/a_544_485#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_33/a_696_458# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_61/a_544_485#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_9/a_1226_296# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_53/a_1141_508#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_71/a_696_458# prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_35/a_112_119#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_23/a_1034_424# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_9/a_544_485#
+ prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_63/a_376_368# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_33/a_1178_124#
+ prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_5/a_376_368# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_13/a_544_485#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_73/a_1034_424# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_21/a_696_458#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_51/a_544_485# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_8/a_1226_296#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_51/a_1141_508# prbs_generator_syn_19/sky130_fd_sc_hs__nand2_1_55/a_117_74#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_21/a_1034_424# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_63/a_1226_296#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_23/a_27_74# prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_7/a_112_119#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_13/a_1226_296# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_8/a_696_458#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_32/a_1178_124# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_49/a_1178_124#
+ prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_37/a_52_123# prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_27/a_132_392#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_71/Q prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_67/a_735_102#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_69/a_1141_508# prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_15/a_112_119#
+ prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_53/a_112_119# prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_39/a_222_392#
+ prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_55/a_230_79# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_19/a_1141_508#
+ prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_37/a_293_74# prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_43/a_376_368#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_5/a_735_102# prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_35/a_138_385#
+ prbs_generator_syn_19/sky130_fd_sc_hs__sdlclkp_2_1/a_114_424# prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_57/a_132_392#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_71/a_1034_424# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_7/a_1226_296#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_33/a_544_485# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_41/a_696_458#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_71/a_544_485# prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_21/B
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_61/a_1226_296# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_39/a_1034_424#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_17/a_27_74# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_9/a_27_74#
+ prbs_generator_syn_19/sky130_fd_sc_hs__nor2b_1_5/a_27_112# prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_47/a_132_392#
+ prbs_generator_syn_19/sky130_fd_sc_hs__nor2b_1_8/a_278_368# prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_9/B
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_39/a_206_368# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_33/a_27_74#
+ prbs_generator_syn_19/sky130_fd_sc_hs__nand2_1_41/a_117_74# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_69/a_651_503#
+ prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_51/a_293_74# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_21/a_544_485#
+ prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_7/a_138_385# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_32/a_696_458#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_47/a_735_102# prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_33/a_112_119#
+ prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_59/a_222_392# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_17/a_1141_508#
+ prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_55/a_52_123# prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_3/a_293_74#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_7/a_651_503# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_29/a_1226_296#
+ prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_23/a_376_368# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_8/a_544_485#
+ prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_47/B prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_47/a_1178_124#
+ prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_15/a_138_385# prbs_generator_syn_19/sky130_fd_sc_hs__sdlclkp_2_1/a_1195_374#
+ prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_53/a_138_385# prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_37/a_132_392#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_29/a_206_368# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_39/a_437_503#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_59/a_651_503# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_37/a_735_102#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_67/a_1141_508# prbs_generator_syn_19/sky130_fd_sc_hs__and2b_2_1/a_27_74#
+ prbs_generator_syn_19/sky130_fd_sc_hs__conb_1_1/a_165_290# prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_55/a_293_74#
+ prbs_generator_syn_19/sky130_fd_sc_hs__nand2_1_45/a_117_74# prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_63/a_112_119#
+ prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_49/a_222_392# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_37/a_1034_424#
+ prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_23/a_293_74# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_15/a_1141_508#
+ prbs_generator_syn_19/sky130_fd_sc_hs__nand2_1_5/a_117_74# prbs_generator_syn_19/m3_13600_13485#
+ prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_5/a_112_119# prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_13/a_376_368#
+ prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_51/a_376_368# prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_7/a_293_74#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_19/a_206_368# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_57/a_206_368#
+ prbs_generator_syn_19/sky130_fd_sc_hs__sdlclkp_2_1/a_318_74# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_29/a_437_503#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_49/a_651_503# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_25/a_27_74#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_5/a_1226_296# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_41/a_544_485#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_27/a_735_102# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_65/a_1141_508#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_65/a_735_102# prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_3/a_230_79#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_35/a_1034_424# prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_13/a_230_79#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_41/a_27_74# prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_3/a_132_392#
+ prbs_generator_syn_19/sky130_fd_sc_hs__nand2_1_49/a_117_74# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_27/a_1226_296#
+ prbs_generator_syn_19/sky130_fd_sc_hs__nand2_1_15/a_117_74# prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_41/a_376_368#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_45/a_1178_124# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_4/a_735_102#
+ prbs_generator_syn_19/sky130_fd_sc_hs__nand2_1_9/a_117_74# prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_33/a_138_385#
+ prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_17/a_132_392# prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_55/a_132_392#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_9/a_1141_508# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_19/a_437_503#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_57/a_437_503# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_4/a_1226_296#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_32/a_544_485# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_17/a_735_102#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_55/a_735_102# prbs_generator_syn_19/m3_13600_2261#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_65/a_27_74# prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_29/a_222_392#
+ prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_43/a_112_119# prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_19/X
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_25/a_1226_296# prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_31/a_376_368#
+ prbs_generator_syn_19/sky130_fd_sc_hs__or2_1_1/a_63_368# prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_17/a_230_79#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_4/a_27_74# prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_61/a_230_79#
+ prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_63/a_138_385# prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_5/a_222_392#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_8/a_1141_508# prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_41/a_293_74#
+ prbs_generator_syn_19/sky130_fd_sc_hs__nand2_1_31/a_117_74# prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_5/a_138_385#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_63/a_1141_508# prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_19/a_222_392#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_13/a_1141_508# prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_3/a_52_123#
+ prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_13/a_52_123# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_43/a_1178_124#
+ prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_61/a_376_368# prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_35/a_132_392#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_67/a_206_368# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_1/a_1226_296#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_69/a_696_458# prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_31/a_230_79#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_35/a_735_102# prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_23/a_112_119#
+ prbs_generator_syn_19/sky130_fd_sc_hs__nand2_1_35/a_117_74# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_59/a_27_74#
+ prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_13/a_293_74# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_5/a_206_368#
+ prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_50/a_376_368# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_7/a_696_458#
+ prbs_generator_syn_19/sky130_fd_sc_hs__nor2b_1_7/a_278_368# prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_17/a_52_123#
+ prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_43/a_138_385# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_7/a_1141_508#
+ prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_61/a_52_123# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_67/a_437_503#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_61/a_1141_508# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_25/a_735_102#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_59/a_696_458# prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_13/a_112_119#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_33/a_1034_424# prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_51/a_112_119#
+ prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_35/a_230_79# prbs_generator_syn_19/m3_13600_4091#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_23/a_1226_296# prbs_generator_syn_19/sky130_fd_sc_hs__nand2_1_39/a_117_74#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_29/a_27_74# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_5/a_437_503#
+ prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_17/a_293_74# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_41/a_1178_124#
+ prbs_generator_syn_19/sky130_fd_sc_hs__or2_1_1/a_152_368# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_59/a_1178_124#
+ prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_61/a_293_74# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_47/a_206_368#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_39/a_651_503# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_49/a_696_458#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_15/a_735_102# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_32/a_1034_424#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_73/a_1226_296# prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_27/a_222_392#
+ prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_41/a_112_119# prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_31/a_52_123#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_49/a_1034_424# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_29/a_1141_508#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_21/a_1226_296# prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_39/a_230_79#
+ prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_23/a_138_385# prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_51/a_230_79#
+ prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_45/a_132_392# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_37/a_206_368#
+ prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_65/a_293_74# prbs_generator_syn_19/sky130_fd_sc_hs__nand2_1_53/a_117_74#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_47/a_437_503# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_29/a_651_503#
+ prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_31/a_293_74# prbs_generator_syn_19/sky130_fd_sc_hs__nand2_1_21/a_117_74#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_69/a_544_485# prbs_generator_syn_19/sky130_fd_sc_hs__clkbuf_16_1/a_114_74#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_45/a_735_102# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_13/a_27_74#
+ prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_31/a_112_119# prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_57/a_222_392#
+ prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_35/a_52_123# prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_21/a_376_368#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_7/a_544_485# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_57/a_1178_124#
+ prbs_generator_syn_19/m3_13600_6043# prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_13/a_138_385#
+ prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_51/a_138_385# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_5/a_1141_508#
+ prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_3/a_376_368# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_27/a_206_368#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_65/a_206_368# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_37/a_437_503#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_19/a_651_503# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_57/a_651_503#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_59/a_544_485# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_71/a_1226_296#
+ prbs_generator_syn_19/sky130_fd_sc_hs__nand2_1_25/a_117_74# prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_61/a_112_119#
+ prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_47/a_222_392# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_27/a_1141_508#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_53/a_27_74# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_4/a_206_368#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_39/a_1226_296# prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_11/a_376_368#
+ prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_39/a_52_123# prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_41/a_138_385#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_4/a_1141_508# prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_25/a_132_392#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_17/a_206_368# prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_41/A
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_55/a_206_368# prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_51/a_52_123#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_27/a_437_503# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_65/a_437_503#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_49/a_544_485# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_63/a_735_102#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_47/a_1034_424# prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_50/a_112_119#
+ prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_37/a_222_392# prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_59/a_230_79#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_25/a_1141_508# prbs_generator_syn_19/sky130_fd_sc_hs__nor2b_1_4/a_27_112#
+ prbs_generator_syn_19/sky130_fd_sc_hs__sdlclkp_2_1/a_685_81# prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_1/a_132_392#
+ prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_39/a_293_74# prbs_generator_syn_19/sky130_fd_sc_hs__nand2_1_29/a_117_74#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_4/a_437_503# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_55/a_1178_124#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_21/a_27_74# prbs_generator_syn_19/m3_13600_12875#
+ prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_50/a_293_74# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_1/a_735_102#
+ prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_31/a_138_385# prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_15/a_132_392#
+ prbs_generator_syn_19/sky130_fd_sc_hs__nand2_1_1/a_117_74# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_17/a_437_503#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_55/a_437_503# prbs_generator_syn
Xprbs_generator_syn_29 prbs_generator_syn_31/clk prbs_generator_syn_31/rst prbs_generator_syn_29/cke
+ sky130_fd_sc_hs__conb_1_265/LO sky130_fd_sc_hs__conb_1_265/LO sky130_fd_sc_hs__conb_1_265/LO
+ sky130_fd_sc_hs__conb_1_265/LO prbs_generator_syn_31/eqn[8] prbs_generator_syn_31/eqn[8]
+ sky130_fd_sc_hs__conb_1_265/LO sky130_fd_sc_hs__conb_1_265/LO sky130_fd_sc_hs__conb_1_265/LO
+ sky130_fd_sc_hs__conb_1_265/LO sky130_fd_sc_hs__conb_1_241/LO sky130_fd_sc_hs__conb_1_241/LO
+ sky130_fd_sc_hs__conb_1_241/LO sky130_fd_sc_hs__conb_1_241/LO sky130_fd_sc_hs__conb_1_241/LO
+ sky130_fd_sc_hs__conb_1_241/LO sky130_fd_sc_hs__conb_1_241/LO sky130_fd_sc_hs__conb_1_241/LO
+ prbs_generator_syn_29/eqn[2] prbs_generator_syn_29/eqn[2] prbs_generator_syn_29/eqn[2]
+ prbs_generator_syn_29/eqn[1] prbs_generator_syn_29/eqn[2] prbs_generator_syn_29/eqn[1]
+ sky130_fd_sc_hs__conb_1_263/LO sky130_fd_sc_hs__conb_1_263/HI sky130_fd_sc_hs__conb_1_263/LO
+ sky130_fd_sc_hs__conb_1_263/HI sky130_fd_sc_hs__conb_1_263/LO sky130_fd_sc_hs__conb_1_263/HI
+ sky130_fd_sc_hs__conb_1_263/LO sky130_fd_sc_hs__conb_1_263/HI prbs_generator_syn_29/eqn[31]
+ prbs_generator_syn_29/eqn[31] prbs_generator_syn_29/eqn[31] prbs_generator_syn_29/eqn[28]
+ prbs_generator_syn_29/eqn[28] prbs_generator_syn_29/eqn[28] prbs_generator_syn_29/eqn[28]
+ prbs_generator_syn_29/eqn[28] prbs_generator_syn_29/eqn[28] prbs_generator_syn_29/eqn[22]
+ prbs_generator_syn_29/eqn[22] prbs_generator_syn_29/eqn[20] prbs_generator_syn_29/eqn[22]
+ prbs_generator_syn_29/eqn[22] prbs_generator_syn_29/eqn[22] prbs_generator_syn_29/eqn[22]
+ prbs_generator_syn_23/eqn[0] prbs_generator_syn_23/eqn[0] prbs_generator_syn_23/eqn[0]
+ prbs_generator_syn_23/eqn[0] prbs_generator_syn_23/eqn[0] prbs_generator_syn_23/eqn[0]
+ prbs_generator_syn_29/eqn[9] prbs_generator_syn_29/eqn[9] prbs_generator_syn_29/eqn[9]
+ prbs_generator_syn_29/eqn[9] prbs_generator_syn_29/eqn[9] prbs_generator_syn_29/eqn[9]
+ prbs_generator_syn_29/eqn[9] prbs_generator_syn_29/eqn[2] prbs_generator_syn_29/eqn[1]
+ prbs_generator_syn_29/eqn[2] prbs_generator_syn_31/inj_err prbs_generator_syn_29/eqn[31]
+ prbs_generator_syn_29/eqn[31] hr_16t4_mux_top_1/din[6] DVSS: DVDD: prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_1/a_293_74#
+ prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_15/X prbs_generator_syn_29/sky130_fd_sc_hs__nand2_1_35/B
+ prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_51/Y prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_9/A
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_9/CLK prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_47/a_27_74#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_37/a_1226_296# prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_3/B
+ prbs_generator_syn_29/sky130_fd_sc_hs__nor2b_1_7/a_27_112# prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_29/B
+ prbs_generator_syn_29/sky130_fd_sc_hs__sdlclkp_2_1/a_580_74# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_1/a_1141_508#
+ prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_5/Y prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_41/a_230_79#
+ prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_61/a_138_385# prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_43/a_132_392#
+ prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_3/a_222_392# prbs_generator_syn_29/sky130_fd_sc_hs__nor2b_1_9/a_27_112#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_61/a_27_74# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_35/a_206_368#
+ prbs_generator_syn_29/sky130_fd_sc_hs__nand2_2_3/Y prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_25/B
+ prbs_generator_syn_29/sky130_fd_sc_hs__nand2_1_11/a_117_74# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_67/a_651_503#
+ prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_45/X prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_39/a_696_458#
+ prbs_generator_syn_29/sky130_fd_sc_hs__sdlclkp_2_1/a_1198_74# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_45/a_1034_424#
+ prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_17/a_222_392# prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_55/a_222_392#
+ prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_53/Y prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_35/A
+ prbs_generator_syn_29/m3_13600_1651# prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_59/a_52_123#
+ prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_5/a_293_74# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_35/a_1226_296#
+ prbs_generator_syn_29/sky130_fd_sc_hs__nand2_1_51/B prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_5/a_651_503#
+ prbs_generator_syn_29/sky130_fd_sc_hs__nand2_1_21/B prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_8/a_27_74#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_15/a_27_74# prbs_generator_syn_29/sky130_fd_sc_hs__and2b_2_1/X
+ prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_13/X prbs_generator_syn_29/sky130_fd_sc_hs__nand2_2_3/a_27_74#
+ prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_50/a_138_385# prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_33/a_132_392#
+ prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_1/a_376_368# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_25/a_206_368#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_35/a_437_503# prbs_generator_syn_29/sky130_fd_sc_hs__sdlclkp_2_1/a_708_451#
+ prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_45/a_230_79# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_29/a_696_458#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_32/a_27_74# prbs_generator_syn_29/sky130_fd_sc_hs__nor2b_1_4/Y
+ prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_59/a_293_74# prbs_generator_syn_29/sky130_fd_sc_hs__nand2_1_47/a_117_74#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_73/a_735_102# prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_21/a_112_119#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_23/a_1141_508# prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_25/a_293_74#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_7/Q prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_3/a_112_119#
+ prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_35/B prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_51/X
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_53/a_1178_124# prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_23/a_132_392#
+ prbs_generator_syn_29/sky130_fd_sc_hs__nand2_1_3/B prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_15/a_206_368#
+ prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_63/a_132_392# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_55/a_27_74#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_25/a_437_503# prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_41/a_52_123#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_47/a_651_503# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_73/a_1141_508#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_19/a_696_458# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_57/a_696_458#
+ prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_7/X prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_43/a_1034_424#
+ prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_55/A prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_11/a_112_119#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_21/a_1141_508# prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_35/a_222_392#
+ prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_49/a_230_79# prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_67/Y
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_71/a_27_74# prbs_generator_syn_29/sky130_fd_sc_hs__nand2_1_33/B
+ prbs_generator_syn_29/sky130_fd_sc_hs__conb_1_1/LO prbs_generator_syn_29/sky130_fd_sc_hs__nand2_1_19/a_117_74#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_51/a_1178_124# prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_33/X
+ prbs_generator_syn_29/sky130_fd_sc_hs__nand2_1_29/B prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_41/Y
+ prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_53/a_132_392# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_45/a_206_368#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_15/a_437_503# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_37/a_651_503#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_39/a_544_485# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_53/a_735_102#
+ prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_45/a_52_123# prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_1/B
+ prbs_generator_syn_29/sky130_fd_sc_hs__nand2_2_3/B prbs_generator_syn_29/sky130_fd_sc_hs__clkbuf_16_1/A
+ prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_21/X prbs_generator_syn_29/sky130_fd_sc_hs__nand2_1_25/B
+ prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_39/a_376_368# prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_63/X
+ prbs_generator_syn_29/m3_13600_3481# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_69/a_1178_124#
+ prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_21/a_138_385# prbs_generator_syn_29/sky130_fd_sc_hs__nor2b_1_8/Y
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_19/a_1178_124# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_49/a_27_74#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_45/a_437_503# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_27/a_651_503#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_71/a_1141_508# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_65/a_651_503#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_29/a_544_485# prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_3/a_138_385#
+ prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_55/X prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_43/a_735_102#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_41/a_1034_424# prbs_generator_syn_29/sky130_fd_sc_hs__nand2_1_9/B
+ prbs_generator_syn_29/sky130_fd_sc_hs__nor2b_1_9/Y prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_59/a_1034_424#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_39/a_1141_508# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_33/a_1226_296#
+ prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_49/a_52_123# prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_47/Y
+ prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_43/Y prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_4/a_651_503#
+ prbs_generator_syn_29/sky130_fd_sc_hs__nand2_1_49/B prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_19/A
+ prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_11/a_138_385# prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_5/X
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_63/a_206_368# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_17/a_651_503#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_19/a_544_485# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_55/a_651_503#
+ prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_9/Y prbs_generator_syn_29/sky130_fd_sc_hs__nand2_1_17/B
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_57/a_544_485# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_67/a_696_458#
+ prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_35/X prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_19/a_27_74#
+ prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_45/a_222_392# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_32/a_1226_296#
+ prbs_generator_syn_29/sky130_fd_sc_hs__nand2_1_43/B prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_25/A
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_1/a_206_368# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_49/a_1226_296#
+ prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_1/a_112_119# prbs_generator_syn_29/sky130_fd_sc_hs__or2_1_1/X
+ prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_59/a_376_368# prbs_generator_syn_29/sky130_fd_sc_hs__nand2_1_19/B
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_5/a_696_458# prbs_generator_syn_29/sky130_fd_sc_hs__nor2b_1_1/Y
+ prbs_generator_syn_29/sky130_fd_sc_hs__nor2b_1_5/a_278_368# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_17/a_1178_124#
+ prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_39/X prbs_generator_syn_29/m3_13600_5433#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_63/a_437_503# prbs_generator_syn_29/sky130_fd_sc_hs__nand2_2_5/B
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_23/a_735_102# prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_53/A
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_61/a_735_102# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_57/a_1034_424#
+ prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_63/B prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_37/a_1141_508#
+ prbs_generator_syn_29/sky130_fd_sc_hs__nand2_1_47/B prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_29/X
+ prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_65/Y prbs_generator_syn_29/m3_13600_4701#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_1/a_437_503# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_67/a_1178_124#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_9/a_735_102# prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_13/a_132_392#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_15/a_1178_124# prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_15/A
+ prbs_generator_syn_29/sky130_fd_sc_hs__nand2_1_1/B prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_43/B
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_35/a_651_503# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_8/D
+ prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_29/A prbs_generator_syn_29/sky130_fd_sc_hs__nand2_1_7/B
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_13/a_735_102# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_47/a_696_458#
+ prbs_generator_syn_29/sky130_fd_sc_hs__nand2_1_31/B prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_51/a_735_102#
+ prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_59/X prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_35/a_1141_508#
+ prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_25/a_222_392# prbs_generator_syn_29/sky130_fd_sc_hs__sdlclkp_2_1/a_288_48#
+ prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_55/B prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_17/B
+ prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_43/A prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_7/A
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_65/a_1178_124# prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_59/Y
+ prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_41/X prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_21/a_230_79#
+ prbs_generator_syn_29/sky130_fd_sc_hs__nand2_1_57/a_117_74# prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_1/a_222_392#
+ prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_19/B prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_35/a_293_74#
+ prbs_generator_syn_29/sky130_fd_sc_hs__nand2_1_23/a_117_74# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_73/a_206_368#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_25/a_651_503# prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_1/a_138_385#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_37/a_696_458# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_67/a_544_485#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_43/a_27_74# prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_9/X
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_55/a_1034_424# prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_39/a_112_119#
+ prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_15/a_222_392# prbs_generator_syn_29/sky130_fd_sc_hs__conb_1_1/HI
+ prbs_generator_syn_29/sky130_fd_sc_hs__nand2_1_23/B prbs_generator_syn_29/sky130_fd_sc_hs__nand2_1_53/B
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_9/a_1178_124# prbs_generator_syn_29/sky130_fd_sc_hs__nor2b_1_4/A
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_47/a_1226_296# prbs_generator_syn_29/m3_13600_11045#
+ prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_17/X prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_29/a_376_368#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_5/a_544_485# prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_3/X
+ prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_31/a_132_392# prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_61/A
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_15/a_651_503# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_73/a_437_503#
+ prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_25/a_230_79# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_27/a_696_458#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_65/a_696_458# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_33/a_735_102#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_71/a_735_102# prbs_generator_syn_29/m3_13600_7263#
+ prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_43/a_222_392# prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_50/Y
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_8/a_1178_124# prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_53/B
+ prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_19/a_376_368# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_63/a_1178_124#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_4/a_696_458# prbs_generator_syn_29/sky130_fd_sc_hs__nor2b_1_4/a_278_368#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_13/a_1178_124# prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_61/a_132_392#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_53/a_206_368# prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_21/a_52_123#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_45/a_651_503# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_17/a_696_458#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_47/a_544_485# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_55/a_696_458#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_21/a_735_102# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_37/a_27_74#
+ prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_61/B prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_61/X
+ prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_59/a_112_119# prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_31/A
+ prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_33/a_222_392# prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_29/a_230_79#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_45/a_1226_296# prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_9/a_132_392#
+ prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_5/A prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_57/Y
+ prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_31/X prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_51/a_27_74#
+ prbs_generator_syn_29/sky130_fd_sc_hs__nor2b_1_8/a_27_112# prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_47/a_376_368#
+ prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_53/a_293_74# prbs_generator_syn_29/sky130_fd_sc_hs__nand2_1_43/a_117_74#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_8/a_735_102# prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_21/a_293_74#
+ prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_39/a_138_385# prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_63/Y
+ prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_51/a_132_392# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_43/a_206_368#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_53/a_437_503# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_37/a_544_485#
+ prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_57/X prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_53/a_1034_424#
+ prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_25/a_52_123# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_33/a_1141_508#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_63/Q prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_23/a_222_392#
+ prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_63/a_222_392# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_7/a_1178_124#
+ prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_53/X prbs_generator_syn_29/sky130_fd_sc_hs__nand2_2_5/Y
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_61/a_1178_124# prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_1/a_230_79#
+ prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_43/a_230_79# prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_11/a_230_79#
+ prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_41/a_132_392# prbs_generator_syn_29/sky130_fd_sc_hs__nand2_1_13/a_117_74#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_43/a_437_503# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_27/a_544_485#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_63/a_651_503# prbs_generator_syn_29/sky130_fd_sc_hs__nand2_1_7/a_117_74#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_35/a_696_458# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_65/a_544_485#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_51/a_1034_424# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_41/a_735_102#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_32/a_1141_508# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_49/a_1141_508#
+ prbs_generator_syn_29/sky130_fd_sc_hs__nand2_1_55/B prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_53/a_222_392#
+ prbs_generator_syn_29/sky130_fd_sc_hs__sdlclkp_2_1/a_114_112# prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_9/a_293_74#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_43/a_1226_296# prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_29/a_52_123#
+ prbs_generator_syn_29/sky130_fd_sc_hs__nand2_1_37/B prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_1/a_651_503#
+ prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_27/a_376_368# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_4/a_544_485#
+ prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_67/a_376_368# prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_27/X
+ prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_1/X prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_59/a_138_385#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_29/a_1178_124# prbs_generator_syn_29/m3_13600_2871#
+ prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_5/a_230_79# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_23/a_206_368#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_61/a_206_368# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_17/a_544_485#
+ prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_15/a_230_79# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_25/a_696_458#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_55/a_544_485# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_32/a_735_102#
+ prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_29/a_293_74# prbs_generator_syn_29/sky130_fd_sc_hs__nand2_1_17/a_117_74#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_69/a_1034_424# prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_29/a_112_119#
+ prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_37/X prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_31/B
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_19/a_1034_424# prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_33/A
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_9/a_206_368# prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_57/a_376_368#
+ prbs_generator_syn_29/sky130_fd_sc_hs__sdlclkp_2_1/a_706_317# prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_11/B
+ prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_1/a_52_123# prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_39/B
+ prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_21/a_132_392# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_13/a_206_368#
+ prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_43/a_52_123# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_51/a_206_368#
+ prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_47/X prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_23/a_437_503#
+ prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_11/a_52_123# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_61/a_437_503#
+ prbs_generator_syn_29/sky130_fd_sc_hs__nor2b_1_7/Y prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_51/A
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_15/a_696_458# prbs_generator_syn_29/sky130_fd_sc_hs__nor2b_1_5/Y
+ prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_9/a_230_79# prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_25/X
+ prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_19/a_112_119# prbs_generator_syn_29/sky130_fd_sc_hs__nand2_1_45/B
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_5/a_1178_124# prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_19/a_230_79#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_41/a_1226_296# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_59/a_1226_296#
+ prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_63/a_230_79# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_51/Q
+ prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_7/a_132_392# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_9/a_437_503#
+ prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_46/a_376_368# prbs_generator_syn_29/sky130_fd_sc_hs__nand2_1_33/a_117_74#
+ prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_11/a_293_74# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_27/a_1178_124#
+ prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_11/a_132_392# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_13/a_437_503#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_51/a_437_503# prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_5/a_52_123#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_35/a_544_485# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_73/a_651_503#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_45/a_696_458# prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_15/a_52_123#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_47/a_1141_508# prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_47/a_112_119#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_4/a_1178_124# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_17/a_1034_424#
+ prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_23/B prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_37/a_376_368#
+ prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_15/B prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_7/Y
+ prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_29/a_138_385# prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_33/a_230_79#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_25/a_1178_124# prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_47/a_293_74#
+ prbs_generator_syn_29/sky130_fd_sc_hs__nand2_1_37/a_117_74# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_33/a_206_368#
+ prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_15/a_293_74# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_71/a_206_368#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_25/a_544_485# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_67/a_1034_424#
+ prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_13/a_222_392# prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_9/a_52_123#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_15/a_1034_424# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_57/a_1226_296#
+ prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_19/a_52_123# prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_23/X
+ prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_63/a_52_123# prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_19/a_138_385#
+ prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_9/a_376_368# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_21/a_206_368#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_33/a_437_503# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_71/a_437_503#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_53/a_651_503# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_15/a_544_485#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_63/a_696_458# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_65/a_1034_424#
+ prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_19/a_293_74# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_45/a_1141_508#
+ prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_27/a_112_119# prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_67/a_112_119#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_1/a_1178_124# prbs_generator_syn_29/sky130_fd_sc_hs__conb_1_1/a_21_290#
+ prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_63/a_293_74# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_8/a_206_368#
+ prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_17/a_376_368# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_63/a_27_74#
+ prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_21/A prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_55/a_376_368#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_1/a_696_458# prbs_generator_syn_29/sky130_fd_sc_hs__nor2b_1_1/a_278_368#
+ prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_47/a_138_385# prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_33/a_52_123#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_9/a_1034_424# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_21/a_437_503#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_1/a_27_74# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_43/a_651_503#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_1/Q prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_45/a_544_485#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_69/a_735_102# prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_57/a_112_119#
+ prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_31/a_222_392# prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_13/A
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_55/a_1226_296# prbs_generator_syn_29/sky130_fd_sc_hs__nand2_2_5/a_27_74#
+ prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_53/a_230_79# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_8/a_437_503#
+ prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_67/a_293_74# prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_33/a_293_74#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_7/a_735_102# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_23/a_1178_124#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_41/a_206_368# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_8/a_1034_424#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_63/a_1034_424# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_59/a_735_102#
+ prbs_generator_syn_29/sky130_fd_sc_hs__nand2_1_5/B prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_43/a_1141_508#
+ prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_46/a_112_119# prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_61/a_222_392#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_13/a_1034_424# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_73/a_1178_124#
+ prbs_generator_syn_29/sky130_fd_sc_hs__nand2_1_27/B prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_13/B
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_57/a_27_74# prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_57/a_230_79#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_21/a_1178_124# prbs_generator_syn_29/sky130_fd_sc_hs__nor2b_1_1/a_27_112#
+ prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_27/a_138_385# prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_23/a_230_79#
+ prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_67/a_138_385# prbs_generator_syn_29/sky130_fd_sc_hs__nand2_1_41/B
+ prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_9/a_222_392# prbs_generator_syn_29/sky130_fd_sc_hs__nand2_1_27/a_117_74#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_32/a_206_368# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_23/a_651_503#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_41/a_437_503# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_73/a_27_74#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_61/a_651_503# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_63/a_544_485#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_49/a_735_102# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_73/a_696_458#
+ prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_37/a_112_119# prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_51/a_222_392#
+ prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_43/X prbs_generator_syn_29/sky130_fd_sc_hs__nand2_2_1/B
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_9/a_651_503# prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_53/a_52_123#
+ prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_49/X prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_25/a_376_368#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_1/a_544_485# prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_65/a_376_368#
+ prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_57/a_138_385# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_27/a_27_74#
+ prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_39/a_132_392# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_7/a_1034_424#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_13/a_651_503# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_32/a_437_503#
+ prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_27/a_230_79# prbs_generator_syn_29/m3_13600_12265#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_51/a_651_503# prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_59/B
+ prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_47/A prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_61/a_1034_424#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_41/a_1141_508# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_59/a_1141_508#
+ prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_41/a_222_392# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_53/a_1226_296#
+ prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_3/A prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_71/a_1178_124#
+ prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_9/a_112_119# prbs_generator_syn_29/sky130_fd_sc_hs__nand2_1_3/a_117_74#
+ prbs_generator_syn_29/m3_13600_8483# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_39/a_1178_124#
+ prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_57/a_52_123# prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_46/a_138_385#
+ prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_23/a_52_123# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_67/a_27_74#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_53/a_696_458# prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_17/a_112_119#
+ prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_11/A prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_55/a_112_119#
+ prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_1/A prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_51/a_1226_296#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_29/a_1034_424# prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_59/A
+ prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_23/A prbs_generator_syn_29/sky130_fd_sc_hs__nand2_1_39/B
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_5/a_27_74# prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_57/a_293_74#
+ prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_37/a_138_385# prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_59/a_132_392#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_33/a_651_503# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_71/a_651_503#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_43/a_696_458# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_73/a_544_485#
+ prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_27/a_52_123# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_57/a_1141_508#
+ prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_21/a_222_392# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_35/a_27_74#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_69/a_1226_296# prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_37/B
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_19/a_1226_296# prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_35/a_376_368#
+ prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_47/a_230_79# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_37/a_1178_124#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_5/a_1034_424# prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_49/a_132_392#
+ prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_7/a_222_392# prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_27/a_293_74#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_21/a_651_503# prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_9/a_138_385#
+ prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_11/a_222_392# prbs_generator_syn_29/m3_13600_14095#
+ prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_50/A prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_27/a_1034_424#
+ prbs_generator_syn_29/sky130_fd_sc_hs__nand2_1_13/B prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_8/a_651_503#
+ prbs_generator_syn_29/m3_13600_9703# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_35/a_1178_124#
+ prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_17/a_138_385# prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_55/a_138_385#
+ prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_7/a_230_79# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_4/a_1034_424#
+ prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_7/a_376_368# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_69/a_206_368#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_23/a_696_458# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_53/a_544_485#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_39/a_735_102# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_61/a_696_458#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_55/a_1141_508# prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_25/a_112_119#
+ prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_65/a_112_119# prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_43/a_293_74#
+ prbs_generator_syn_29/sky130_fd_sc_hs__nand2_1_57/B prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_25/a_1034_424#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_7/a_206_368# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_17/a_1226_296#
+ prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_15/a_376_368# prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_53/a_376_368#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_9/a_696_458# prbs_generator_syn_29/m3_13600_431#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_45/a_27_74# prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_47/a_52_123#
+ prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_29/a_132_392# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_59/a_206_368#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_69/a_437_503# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_41/a_651_503#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_43/a_544_485# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_13/a_696_458#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_29/a_735_102# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_51/a_696_458#
+ prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_61/Y prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_67/a_1226_296#
+ prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_5/a_132_392# prbs_generator_syn_29/sky130_fd_sc_hs__and2b_2_1/a_198_48#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_7/a_437_503# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_15/a_1226_296#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_69/a_27_74# prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_46/a_293_74#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_1/a_1034_424# prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_19/a_132_392#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_49/a_206_368# prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_7/a_52_123#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_59/a_437_503# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_32/a_651_503#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_7/a_27_74# prbs_generator_syn_29/sky130_fd_sc_hs__nand2_2_1/a_27_74#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_19/a_735_102# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_57/a_735_102#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_65/a_1226_296# prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_37/A
+ prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_33/a_376_368# prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_37/a_230_79#
+ prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_25/a_138_385# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_39/a_27_74#
+ prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_65/a_138_385# prbs_generator_syn_29/sky130_fd_sc_hs__nor2b_1_9/a_278_368#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_49/a_437_503# prbs_generator_syn_29/sky130_fd_sc_hs__and2b_2_1/a_505_74#
+ prbs_generator_syn_29/sky130_fd_sc_hs__nand2_1_51/a_117_74# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_23/a_544_485#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_33/a_696_458# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_61/a_544_485#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_9/a_1226_296# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_53/a_1141_508#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_71/a_696_458# prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_35/a_112_119#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_23/a_1034_424# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_9/a_544_485#
+ prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_63/a_376_368# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_33/a_1178_124#
+ prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_5/a_376_368# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_13/a_544_485#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_73/a_1034_424# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_21/a_696_458#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_51/a_544_485# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_8/a_1226_296#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_51/a_1141_508# prbs_generator_syn_29/sky130_fd_sc_hs__nand2_1_55/a_117_74#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_21/a_1034_424# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_63/a_1226_296#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_23/a_27_74# prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_7/a_112_119#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_13/a_1226_296# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_8/a_696_458#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_32/a_1178_124# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_49/a_1178_124#
+ prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_37/a_52_123# prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_27/a_132_392#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_71/Q prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_67/a_735_102#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_69/a_1141_508# prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_15/a_112_119#
+ prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_53/a_112_119# prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_39/a_222_392#
+ prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_55/a_230_79# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_19/a_1141_508#
+ prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_37/a_293_74# prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_43/a_376_368#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_5/a_735_102# prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_35/a_138_385#
+ prbs_generator_syn_29/sky130_fd_sc_hs__sdlclkp_2_1/a_114_424# prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_57/a_132_392#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_71/a_1034_424# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_7/a_1226_296#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_33/a_544_485# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_41/a_696_458#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_71/a_544_485# prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_21/B
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_61/a_1226_296# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_39/a_1034_424#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_17/a_27_74# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_9/a_27_74#
+ prbs_generator_syn_29/sky130_fd_sc_hs__nor2b_1_5/a_27_112# prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_47/a_132_392#
+ prbs_generator_syn_29/sky130_fd_sc_hs__nor2b_1_8/a_278_368# prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_9/B
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_39/a_206_368# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_33/a_27_74#
+ prbs_generator_syn_29/sky130_fd_sc_hs__nand2_1_41/a_117_74# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_69/a_651_503#
+ prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_51/a_293_74# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_21/a_544_485#
+ prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_7/a_138_385# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_32/a_696_458#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_47/a_735_102# prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_33/a_112_119#
+ prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_59/a_222_392# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_17/a_1141_508#
+ prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_55/a_52_123# prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_3/a_293_74#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_7/a_651_503# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_29/a_1226_296#
+ prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_23/a_376_368# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_8/a_544_485#
+ prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_47/B prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_47/a_1178_124#
+ prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_15/a_138_385# prbs_generator_syn_29/sky130_fd_sc_hs__sdlclkp_2_1/a_1195_374#
+ prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_53/a_138_385# prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_37/a_132_392#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_29/a_206_368# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_39/a_437_503#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_59/a_651_503# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_37/a_735_102#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_67/a_1141_508# prbs_generator_syn_29/sky130_fd_sc_hs__and2b_2_1/a_27_74#
+ prbs_generator_syn_29/sky130_fd_sc_hs__conb_1_1/a_165_290# prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_55/a_293_74#
+ prbs_generator_syn_29/sky130_fd_sc_hs__nand2_1_45/a_117_74# prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_63/a_112_119#
+ prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_49/a_222_392# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_37/a_1034_424#
+ prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_23/a_293_74# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_15/a_1141_508#
+ prbs_generator_syn_29/sky130_fd_sc_hs__nand2_1_5/a_117_74# prbs_generator_syn_29/m3_13600_13485#
+ prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_5/a_112_119# prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_13/a_376_368#
+ prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_51/a_376_368# prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_7/a_293_74#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_19/a_206_368# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_57/a_206_368#
+ prbs_generator_syn_29/sky130_fd_sc_hs__sdlclkp_2_1/a_318_74# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_29/a_437_503#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_49/a_651_503# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_25/a_27_74#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_5/a_1226_296# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_41/a_544_485#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_27/a_735_102# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_65/a_1141_508#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_65/a_735_102# prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_3/a_230_79#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_35/a_1034_424# prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_13/a_230_79#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_41/a_27_74# prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_3/a_132_392#
+ prbs_generator_syn_29/sky130_fd_sc_hs__nand2_1_49/a_117_74# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_27/a_1226_296#
+ prbs_generator_syn_29/sky130_fd_sc_hs__nand2_1_15/a_117_74# prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_41/a_376_368#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_45/a_1178_124# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_4/a_735_102#
+ prbs_generator_syn_29/sky130_fd_sc_hs__nand2_1_9/a_117_74# prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_33/a_138_385#
+ prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_17/a_132_392# prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_55/a_132_392#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_9/a_1141_508# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_19/a_437_503#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_57/a_437_503# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_4/a_1226_296#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_32/a_544_485# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_17/a_735_102#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_55/a_735_102# prbs_generator_syn_29/m3_13600_2261#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_65/a_27_74# prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_29/a_222_392#
+ prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_43/a_112_119# prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_19/X
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_25/a_1226_296# prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_31/a_376_368#
+ prbs_generator_syn_29/sky130_fd_sc_hs__or2_1_1/a_63_368# prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_17/a_230_79#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_4/a_27_74# prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_61/a_230_79#
+ prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_63/a_138_385# prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_5/a_222_392#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_8/a_1141_508# prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_41/a_293_74#
+ prbs_generator_syn_29/sky130_fd_sc_hs__nand2_1_31/a_117_74# prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_5/a_138_385#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_63/a_1141_508# prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_19/a_222_392#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_13/a_1141_508# prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_3/a_52_123#
+ prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_13/a_52_123# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_43/a_1178_124#
+ prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_61/a_376_368# prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_35/a_132_392#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_67/a_206_368# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_1/a_1226_296#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_69/a_696_458# prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_31/a_230_79#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_35/a_735_102# prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_23/a_112_119#
+ prbs_generator_syn_29/sky130_fd_sc_hs__nand2_1_35/a_117_74# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_59/a_27_74#
+ prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_13/a_293_74# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_5/a_206_368#
+ prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_50/a_376_368# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_7/a_696_458#
+ prbs_generator_syn_29/sky130_fd_sc_hs__nor2b_1_7/a_278_368# prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_17/a_52_123#
+ prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_43/a_138_385# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_7/a_1141_508#
+ prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_61/a_52_123# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_67/a_437_503#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_61/a_1141_508# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_25/a_735_102#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_59/a_696_458# prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_13/a_112_119#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_33/a_1034_424# prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_51/a_112_119#
+ prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_35/a_230_79# prbs_generator_syn_29/m3_13600_4091#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_23/a_1226_296# prbs_generator_syn_29/sky130_fd_sc_hs__nand2_1_39/a_117_74#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_29/a_27_74# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_5/a_437_503#
+ prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_17/a_293_74# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_41/a_1178_124#
+ prbs_generator_syn_29/sky130_fd_sc_hs__or2_1_1/a_152_368# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_59/a_1178_124#
+ prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_61/a_293_74# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_47/a_206_368#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_39/a_651_503# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_49/a_696_458#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_15/a_735_102# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_32/a_1034_424#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_73/a_1226_296# prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_27/a_222_392#
+ prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_41/a_112_119# prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_31/a_52_123#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_49/a_1034_424# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_29/a_1141_508#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_21/a_1226_296# prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_39/a_230_79#
+ prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_23/a_138_385# prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_51/a_230_79#
+ prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_45/a_132_392# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_37/a_206_368#
+ prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_65/a_293_74# prbs_generator_syn_29/sky130_fd_sc_hs__nand2_1_53/a_117_74#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_47/a_437_503# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_29/a_651_503#
+ prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_31/a_293_74# prbs_generator_syn_29/sky130_fd_sc_hs__nand2_1_21/a_117_74#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_69/a_544_485# prbs_generator_syn_29/sky130_fd_sc_hs__clkbuf_16_1/a_114_74#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_45/a_735_102# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_13/a_27_74#
+ prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_31/a_112_119# prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_57/a_222_392#
+ prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_35/a_52_123# prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_21/a_376_368#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_7/a_544_485# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_57/a_1178_124#
+ prbs_generator_syn_29/m3_13600_6043# prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_13/a_138_385#
+ prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_51/a_138_385# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_5/a_1141_508#
+ prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_3/a_376_368# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_27/a_206_368#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_65/a_206_368# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_37/a_437_503#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_19/a_651_503# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_57/a_651_503#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_59/a_544_485# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_71/a_1226_296#
+ prbs_generator_syn_29/sky130_fd_sc_hs__nand2_1_25/a_117_74# prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_61/a_112_119#
+ prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_47/a_222_392# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_27/a_1141_508#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_53/a_27_74# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_4/a_206_368#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_39/a_1226_296# prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_11/a_376_368#
+ prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_39/a_52_123# prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_41/a_138_385#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_4/a_1141_508# prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_25/a_132_392#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_17/a_206_368# prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_41/A
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_55/a_206_368# prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_51/a_52_123#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_27/a_437_503# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_65/a_437_503#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_49/a_544_485# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_63/a_735_102#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_47/a_1034_424# prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_50/a_112_119#
+ prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_37/a_222_392# prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_59/a_230_79#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_25/a_1141_508# prbs_generator_syn_29/sky130_fd_sc_hs__nor2b_1_4/a_27_112#
+ prbs_generator_syn_29/sky130_fd_sc_hs__sdlclkp_2_1/a_685_81# prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_1/a_132_392#
+ prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_39/a_293_74# prbs_generator_syn_29/sky130_fd_sc_hs__nand2_1_29/a_117_74#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_4/a_437_503# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_55/a_1178_124#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_21/a_27_74# prbs_generator_syn_29/m3_13600_12875#
+ prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_50/a_293_74# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_1/a_735_102#
+ prbs_generator_syn_29/sky130_fd_sc_hs__xnor2_1_31/a_138_385# prbs_generator_syn_29/sky130_fd_sc_hs__a22o_1_15/a_132_392#
+ prbs_generator_syn_29/sky130_fd_sc_hs__nand2_1_1/a_117_74# prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_17/a_437_503#
+ prbs_generator_syn_29/sky130_fd_sc_hs__dfxtp_4_55/a_437_503# prbs_generator_syn
Xsky130_fd_sc_hs__conb_1_9 DVSS: DVDD: DVDD: DVSS: prbs_generator_syn_3/eqn[8] sky130_fd_sc_hs__conb_1_9/HI
+ sky130_fd_sc_hs__conb_1_9/a_165_290# sky130_fd_sc_hs__conb_1_9/a_21_290# sky130_fd_sc_hs__conb_1
Xsky130_fd_sc_hs__buf_2_105 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__buf_2_105/A sky130_fd_sc_hs__buf_2_105/X
+ sky130_fd_sc_hs__buf_2_105/a_21_260# sky130_fd_sc_hs__buf_2
Xsky130_fd_sc_hs__buf_2_116 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__buf_2_117/A sky130_fd_sc_hs__buf_2_117/X
+ sky130_fd_sc_hs__buf_2_117/a_21_260# sky130_fd_sc_hs__buf_2
Xsky130_fd_sc_hs__buf_2_127 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__buf_2_127/A sky130_fd_sc_hs__buf_2_15/A
+ sky130_fd_sc_hs__buf_2_127/a_21_260# sky130_fd_sc_hs__buf_2
Xsky130_fd_sc_hs__buf_2_138 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__buf_2_139/A sky130_fd_sc_hs__buf_2_139/X
+ sky130_fd_sc_hs__buf_2_139/a_21_260# sky130_fd_sc_hs__buf_2
Xsky130_fd_sc_hs__buf_2_149 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__buf_2_149/A sky130_fd_sc_hs__buf_2_153/A
+ sky130_fd_sc_hs__buf_2_149/a_21_260# sky130_fd_sc_hs__buf_2
Xsky130_fd_sc_hs__einvp_2_17 DVSS: DVDD: DVDD: DVSS: dout_n sky130_fd_sc_hs__einvp_2_9/A
+ sky130_fd_sc_hs__dlrtp_1_5/Q sky130_fd_sc_hs__einvp_2_17/a_263_323# sky130_fd_sc_hs__einvp_2_17/a_36_74#
+ sky130_fd_sc_hs__einvp_2_17/a_27_368# sky130_fd_sc_hs__einvp_2
Xsky130_fd_sc_hs__einvp_2_28 DVSS: DVDD: DVDD: DVSS: dout_n sky130_fd_sc_hs__buf_8_1/A
+ sky130_fd_sc_hs__dlrtp_1_25/Q sky130_fd_sc_hs__einvp_2_29/a_263_323# sky130_fd_sc_hs__einvp_2_29/a_36_74#
+ sky130_fd_sc_hs__einvp_2_29/a_27_368# sky130_fd_sc_hs__einvp_2
Xsky130_fd_sc_hs__einvp_2_39 DVSS: DVDD: DVDD: DVSS: dout_n sky130_fd_sc_hs__buf_8_1/A
+ sky130_fd_sc_hs__buf_2_17/X sky130_fd_sc_hs__einvp_2_39/a_263_323# sky130_fd_sc_hs__einvp_2_39/a_36_74#
+ sky130_fd_sc_hs__einvp_2_39/a_27_368# sky130_fd_sc_hs__einvp_2
Xsky130_fd_sc_hs__conb_1_16 DVSS: DVDD: DVDD: DVSS: prbs_generator_syn_3/eqn[22] prbs_generator_syn_3/eqn[20]
+ sky130_fd_sc_hs__conb_1_17/a_165_290# sky130_fd_sc_hs__conb_1_17/a_21_290# sky130_fd_sc_hs__conb_1
Xsky130_fd_sc_hs__conb_1_27 DVSS: DVDD: DVDD: DVSS: prbs_generator_syn_5/eqn[13] sky130_fd_sc_hs__conb_1_27/HI
+ sky130_fd_sc_hs__conb_1_27/a_165_290# sky130_fd_sc_hs__conb_1_27/a_21_290# sky130_fd_sc_hs__conb_1
Xsky130_fd_sc_hs__conb_1_38 DVSS: DVDD: DVDD: DVSS: prbs_generator_syn_9/eqn[28] sky130_fd_sc_hs__conb_1_39/HI
+ sky130_fd_sc_hs__conb_1_39/a_165_290# sky130_fd_sc_hs__conb_1_39/a_21_290# sky130_fd_sc_hs__conb_1
Xsky130_fd_sc_hs__conb_1_49 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__conb_1_49/LO
+ sky130_fd_sc_hs__conb_1_49/HI sky130_fd_sc_hs__conb_1_49/a_165_290# sky130_fd_sc_hs__conb_1_49/a_21_290#
+ sky130_fd_sc_hs__conb_1
Xsky130_fd_sc_hs__inv_4_12 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__inv_4_13/Y sky130_fd_sc_hs__inv_4_13/A
+ sky130_fd_sc_hs__inv_4
Xsky130_fd_sc_hs__inv_4_23 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__inv_4_23/Y sky130_fd_sc_hs__inv_4_23/A
+ sky130_fd_sc_hs__inv_4
Xsky130_fd_sc_hs__inv_4_34 DVSS: DVDD: DVDD: DVSS: osc_core_1/pi1_r[0] osc_core_1/pi1_l[0]
+ sky130_fd_sc_hs__inv_4
Xsky130_fd_sc_hs__inv_4_45 DVSS: DVDD: DVDD: DVSS: osc_core_1/pi3_r[3] osc_core_1/pi3_l[3]
+ sky130_fd_sc_hs__inv_4
Xsky130_fd_sc_hs__inv_4_56 DVSS: DVDD: DVDD: DVSS: osc_core_1/pi3_r[0] osc_core_1/pi3_l[0]
+ sky130_fd_sc_hs__inv_4
Xsky130_fd_sc_hs__inv_4_67 DVSS: DVDD: DVDD: DVSS: hr_16t4_mux_top_3/din[1] hr_16t4_mux_top_1/din[1]
+ sky130_fd_sc_hs__inv_4
Xsky130_fd_sc_hs__inv_4_78 DVSS: DVDD: DVDD: DVSS: hr_16t4_mux_top_3/din[12] prbs_generator_syn_21/out
+ sky130_fd_sc_hs__inv_4
Xsky130_fd_sc_hs__inv_4_89 DVSS: DVDD: DVDD: DVSS: hr_16t4_mux_top_3/din[0] hr_16t4_mux_top_1/din[0]
+ sky130_fd_sc_hs__inv_4
Xsky130_fd_sc_hs__dlrtp_1_18 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__dlrtp_1_19/Q
+ sky130_fd_sc_hs__dlrtp_1_9/GATE sky130_fd_sc_hs__conb_1_121/HI sky130_fd_sc_hs__dlrtp_1_19/D
+ sky130_fd_sc_hs__dlrtp_1_19/a_216_424# sky130_fd_sc_hs__dlrtp_1_19/a_759_508# sky130_fd_sc_hs__dlrtp_1_19/a_565_74#
+ sky130_fd_sc_hs__dlrtp_1_19/a_27_424# sky130_fd_sc_hs__dlrtp_1_19/a_1045_74# sky130_fd_sc_hs__dlrtp_1_19/a_643_74#
+ sky130_fd_sc_hs__dlrtp_1_19/a_817_48# sky130_fd_sc_hs__dlrtp_1_19/a_568_392# sky130_fd_sc_hs__dlrtp_1_19/a_363_74#
+ sky130_fd_sc_hs__dlrtp_1_19/a_769_74# sky130_fd_sc_hs__dlrtp_1
Xsky130_fd_sc_hs__dlrtp_1_29 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__dlrtp_1_29/Q
+ sky130_fd_sc_hs__clkbuf_2_3/A sky130_fd_sc_hs__conb_1_123/HI sky130_fd_sc_hs__dlrtp_1_29/D
+ sky130_fd_sc_hs__dlrtp_1_29/a_216_424# sky130_fd_sc_hs__dlrtp_1_29/a_759_508# sky130_fd_sc_hs__dlrtp_1_29/a_565_74#
+ sky130_fd_sc_hs__dlrtp_1_29/a_27_424# sky130_fd_sc_hs__dlrtp_1_29/a_1045_74# sky130_fd_sc_hs__dlrtp_1_29/a_643_74#
+ sky130_fd_sc_hs__dlrtp_1_29/a_817_48# sky130_fd_sc_hs__dlrtp_1_29/a_568_392# sky130_fd_sc_hs__dlrtp_1_29/a_363_74#
+ sky130_fd_sc_hs__dlrtp_1_29/a_769_74# sky130_fd_sc_hs__dlrtp_1
Xsky130_fd_sc_hs__clkbuf_16_50 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__clkbuf_16_53/A
+ sky130_fd_sc_hs__nand2_2_7/Y sky130_fd_sc_hs__clkbuf_16_51/a_114_74# sky130_fd_sc_hs__clkbuf_16
Xsky130_fd_sc_hs__clkbuf_16_61 DVSS: DVDD: DVDD: DVSS: qr_4t1_mux_top_3/clk_I sky130_fd_sc_hs__einvn_2_1/Z
+ sky130_fd_sc_hs__clkbuf_16_61/a_114_74# sky130_fd_sc_hs__clkbuf_16
Xsky130_fd_sc_hs__clkbuf_16_72 DVSS: DVDD: DVDD: DVSS: prbs_generator_syn_19/clk sky130_fd_sc_hs__clkbuf_16_75/X
+ sky130_fd_sc_hs__clkbuf_16_73/a_114_74# sky130_fd_sc_hs__clkbuf_16
Xsky130_fd_sc_hs__clkbuf_16_83 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__nor2_4_1/A
+ sky130_fd_sc_hs__clkbuf_4_113/X sky130_fd_sc_hs__clkbuf_16_83/a_114_74# sky130_fd_sc_hs__clkbuf_16
Xsky130_fd_sc_hs__clkbuf_16_94 DVSS: DVDD: DVDD: DVSS: osc_core_1/glob_en osc_en sky130_fd_sc_hs__clkbuf_16_95/a_114_74#
+ sky130_fd_sc_hs__clkbuf_16
Xsky130_fd_sc_hs__nand2_2_13 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__buf_2_87/A sky130_fd_sc_hs__buf_8_3/X
+ sky130_fd_sc_hs__inv_4_21/Y sky130_fd_sc_hs__nand2_2_13/a_27_74# sky130_fd_sc_hs__nand2_2
Xsky130_fd_sc_hs__nand2_2_24 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__nand2_2_25/Y
+ sky130_fd_sc_hs__nor4_2_1/B sky130_fd_sc_hs__nor4_2_1/A sky130_fd_sc_hs__nand2_2_25/a_27_74#
+ sky130_fd_sc_hs__nand2_2
Xprbs_generator_syn_2 prbs_generator_syn_9/clk prbs_generator_syn_9/rst prbs_generator_syn_3/cke
+ sky130_fd_sc_hs__conb_1_49/LO sky130_fd_sc_hs__conb_1_49/LO sky130_fd_sc_hs__conb_1_49/LO
+ prbs_generator_syn_7/eqn[1] prbs_generator_syn_7/eqn[1] prbs_generator_syn_7/eqn[1]
+ prbs_generator_syn_7/eqn[1] prbs_generator_syn_7/eqn[1] sky130_fd_sc_hs__conb_1_49/HI
+ sky130_fd_sc_hs__conb_1_49/HI sky130_fd_sc_hs__conb_1_49/HI prbs_generator_syn_3/cke
+ prbs_generator_syn_3/cke prbs_generator_syn_3/cke prbs_generator_syn_7/eqn[9] sky130_fd_sc_hs__conb_1_51/HI
+ prbs_generator_syn_7/eqn[9] sky130_fd_sc_hs__conb_1_51/HI prbs_generator_syn_9/eqn[16]
+ prbs_generator_syn_9/eqn[16] prbs_generator_syn_9/eqn[22] prbs_generator_syn_9/eqn[22]
+ prbs_generator_syn_9/eqn[22] prbs_generator_syn_9/eqn[28] sky130_fd_sc_hs__conb_1_39/HI
+ sky130_fd_sc_hs__conb_1_39/HI prbs_generator_syn_9/eqn[28] prbs_generator_syn_9/eqn[30]
+ sky130_fd_sc_hs__conb_1_55/HI sky130_fd_sc_hs__conb_1_55/HI prbs_generator_syn_9/eqn[30]
+ prbs_generator_syn_9/eqn[30] prbs_generator_syn_3/eqn[31] prbs_generator_syn_3/eqn[30]
+ prbs_generator_syn_3/eqn[30] prbs_generator_syn_3/eqn[28] prbs_generator_syn_3/eqn[28]
+ prbs_generator_syn_3/eqn[28] prbs_generator_syn_3/eqn[28] prbs_generator_syn_3/eqn[28]
+ prbs_generator_syn_3/eqn[28] prbs_generator_syn_3/eqn[22] prbs_generator_syn_3/eqn[22]
+ prbs_generator_syn_3/eqn[20] prbs_generator_syn_3/eqn[22] prbs_generator_syn_3/eqn[22]
+ prbs_generator_syn_3/eqn[22] prbs_generator_syn_3/eqn[22] prbs_generator_syn_3/eqn[22]
+ prbs_generator_syn_3/eqn[9] prbs_generator_syn_3/eqn[9] prbs_generator_syn_3/eqn[9]
+ prbs_generator_syn_3/eqn[9] prbs_generator_syn_3/eqn[9] prbs_generator_syn_3/eqn[9]
+ prbs_generator_syn_3/eqn[8] prbs_generator_syn_3/eqn[8] prbs_generator_syn_3/eqn[8]
+ prbs_generator_syn_3/eqn[8] prbs_generator_syn_3/eqn[4] prbs_generator_syn_3/eqn[4]
+ prbs_generator_syn_3/eqn[4] prbs_generator_syn_3/eqn[1] prbs_generator_syn_3/eqn[4]
+ prbs_generator_syn_9/inj_err prbs_generator_syn_7/eqn[9] prbs_generator_syn_3/eqn[31]
+ prbs_generator_syn_3/out DVSS: DVDD: prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_1/a_293_74#
+ prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_15/X prbs_generator_syn_3/sky130_fd_sc_hs__nand2_1_35/B
+ prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_51/Y prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_9/A
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_9/CLK prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_47/a_27_74#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_37/a_1226_296# prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_3/B
+ prbs_generator_syn_3/sky130_fd_sc_hs__nor2b_1_7/a_27_112# prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_29/B
+ prbs_generator_syn_3/sky130_fd_sc_hs__sdlclkp_2_1/a_580_74# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_1/a_1141_508#
+ prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_5/Y prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_41/a_230_79#
+ prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_61/a_138_385# prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_43/a_132_392#
+ prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_3/a_222_392# prbs_generator_syn_3/sky130_fd_sc_hs__nor2b_1_9/a_27_112#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_61/a_27_74# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_35/a_206_368#
+ prbs_generator_syn_3/sky130_fd_sc_hs__nand2_2_3/Y prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_25/B
+ prbs_generator_syn_3/sky130_fd_sc_hs__nand2_1_11/a_117_74# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_67/a_651_503#
+ prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_45/X prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_39/a_696_458#
+ prbs_generator_syn_3/sky130_fd_sc_hs__sdlclkp_2_1/a_1198_74# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_45/a_1034_424#
+ prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_17/a_222_392# prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_55/a_222_392#
+ prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_53/Y prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_35/A
+ prbs_generator_syn_3/m3_13600_1651# prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_59/a_52_123#
+ prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_5/a_293_74# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_35/a_1226_296#
+ prbs_generator_syn_3/sky130_fd_sc_hs__nand2_1_51/B prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_5/a_651_503#
+ prbs_generator_syn_3/sky130_fd_sc_hs__nand2_1_21/B prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_8/a_27_74#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_15/a_27_74# prbs_generator_syn_3/sky130_fd_sc_hs__and2b_2_1/X
+ prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_13/X prbs_generator_syn_3/sky130_fd_sc_hs__nand2_2_3/a_27_74#
+ prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_50/a_138_385# prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_33/a_132_392#
+ prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_1/a_376_368# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_25/a_206_368#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_35/a_437_503# prbs_generator_syn_3/sky130_fd_sc_hs__sdlclkp_2_1/a_708_451#
+ prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_45/a_230_79# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_29/a_696_458#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_32/a_27_74# prbs_generator_syn_3/sky130_fd_sc_hs__nor2b_1_4/Y
+ prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_59/a_293_74# prbs_generator_syn_3/sky130_fd_sc_hs__nand2_1_47/a_117_74#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_73/a_735_102# prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_21/a_112_119#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_23/a_1141_508# prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_25/a_293_74#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_7/Q prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_3/a_112_119#
+ prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_35/B prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_51/X
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_53/a_1178_124# prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_23/a_132_392#
+ prbs_generator_syn_3/sky130_fd_sc_hs__nand2_1_3/B prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_15/a_206_368#
+ prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_63/a_132_392# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_55/a_27_74#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_25/a_437_503# prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_41/a_52_123#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_47/a_651_503# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_73/a_1141_508#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_19/a_696_458# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_57/a_696_458#
+ prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_7/X prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_43/a_1034_424#
+ prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_55/A prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_11/a_112_119#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_21/a_1141_508# prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_35/a_222_392#
+ prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_49/a_230_79# prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_67/Y
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_71/a_27_74# prbs_generator_syn_3/sky130_fd_sc_hs__nand2_1_33/B
+ prbs_generator_syn_3/sky130_fd_sc_hs__conb_1_1/LO prbs_generator_syn_3/sky130_fd_sc_hs__nand2_1_19/a_117_74#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_51/a_1178_124# prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_33/X
+ prbs_generator_syn_3/sky130_fd_sc_hs__nand2_1_29/B prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_41/Y
+ prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_53/a_132_392# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_45/a_206_368#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_15/a_437_503# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_37/a_651_503#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_39/a_544_485# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_53/a_735_102#
+ prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_45/a_52_123# prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_1/B
+ prbs_generator_syn_3/sky130_fd_sc_hs__nand2_2_3/B prbs_generator_syn_3/sky130_fd_sc_hs__clkbuf_16_1/A
+ prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_21/X prbs_generator_syn_3/sky130_fd_sc_hs__nand2_1_25/B
+ prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_39/a_376_368# prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_63/X
+ prbs_generator_syn_3/m3_13600_3481# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_69/a_1178_124#
+ prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_21/a_138_385# prbs_generator_syn_3/sky130_fd_sc_hs__nor2b_1_8/Y
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_19/a_1178_124# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_49/a_27_74#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_45/a_437_503# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_27/a_651_503#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_71/a_1141_508# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_65/a_651_503#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_29/a_544_485# prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_3/a_138_385#
+ prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_55/X prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_43/a_735_102#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_41/a_1034_424# prbs_generator_syn_3/sky130_fd_sc_hs__nand2_1_9/B
+ prbs_generator_syn_3/sky130_fd_sc_hs__nor2b_1_9/Y prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_59/a_1034_424#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_39/a_1141_508# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_33/a_1226_296#
+ prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_49/a_52_123# prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_47/Y
+ prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_43/Y prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_4/a_651_503#
+ prbs_generator_syn_3/sky130_fd_sc_hs__nand2_1_49/B prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_19/A
+ prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_11/a_138_385# prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_5/X
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_63/a_206_368# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_17/a_651_503#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_19/a_544_485# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_55/a_651_503#
+ prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_9/Y prbs_generator_syn_3/sky130_fd_sc_hs__nand2_1_17/B
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_57/a_544_485# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_67/a_696_458#
+ prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_35/X prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_19/a_27_74#
+ prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_45/a_222_392# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_32/a_1226_296#
+ prbs_generator_syn_3/sky130_fd_sc_hs__nand2_1_43/B prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_25/A
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_1/a_206_368# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_49/a_1226_296#
+ prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_1/a_112_119# prbs_generator_syn_3/sky130_fd_sc_hs__or2_1_1/X
+ prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_59/a_376_368# prbs_generator_syn_3/sky130_fd_sc_hs__nand2_1_19/B
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_5/a_696_458# prbs_generator_syn_3/sky130_fd_sc_hs__nor2b_1_1/Y
+ prbs_generator_syn_3/sky130_fd_sc_hs__nor2b_1_5/a_278_368# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_17/a_1178_124#
+ prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_39/X prbs_generator_syn_3/m3_13600_5433#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_63/a_437_503# prbs_generator_syn_3/sky130_fd_sc_hs__nand2_2_5/B
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_23/a_735_102# prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_53/A
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_61/a_735_102# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_57/a_1034_424#
+ prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_63/B prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_37/a_1141_508#
+ prbs_generator_syn_3/sky130_fd_sc_hs__nand2_1_47/B prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_29/X
+ prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_65/Y prbs_generator_syn_3/m3_13600_4701#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_1/a_437_503# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_67/a_1178_124#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_9/a_735_102# prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_13/a_132_392#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_15/a_1178_124# prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_15/A
+ prbs_generator_syn_3/sky130_fd_sc_hs__nand2_1_1/B prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_43/B
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_35/a_651_503# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_8/D
+ prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_29/A prbs_generator_syn_3/sky130_fd_sc_hs__nand2_1_7/B
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_13/a_735_102# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_47/a_696_458#
+ prbs_generator_syn_3/sky130_fd_sc_hs__nand2_1_31/B prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_51/a_735_102#
+ prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_59/X prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_35/a_1141_508#
+ prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_25/a_222_392# prbs_generator_syn_3/sky130_fd_sc_hs__sdlclkp_2_1/a_288_48#
+ prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_55/B prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_17/B
+ prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_43/A prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_7/A
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_65/a_1178_124# prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_59/Y
+ prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_41/X prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_21/a_230_79#
+ prbs_generator_syn_3/sky130_fd_sc_hs__nand2_1_57/a_117_74# prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_1/a_222_392#
+ prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_19/B prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_35/a_293_74#
+ prbs_generator_syn_3/sky130_fd_sc_hs__nand2_1_23/a_117_74# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_73/a_206_368#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_25/a_651_503# prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_1/a_138_385#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_37/a_696_458# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_67/a_544_485#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_43/a_27_74# prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_9/X
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_55/a_1034_424# prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_39/a_112_119#
+ prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_15/a_222_392# prbs_generator_syn_3/sky130_fd_sc_hs__conb_1_1/HI
+ prbs_generator_syn_3/sky130_fd_sc_hs__nand2_1_23/B prbs_generator_syn_3/sky130_fd_sc_hs__nand2_1_53/B
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_9/a_1178_124# prbs_generator_syn_3/sky130_fd_sc_hs__nor2b_1_4/A
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_47/a_1226_296# prbs_generator_syn_3/m3_13600_11045#
+ prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_17/X prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_29/a_376_368#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_5/a_544_485# prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_3/X
+ prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_31/a_132_392# prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_61/A
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_15/a_651_503# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_73/a_437_503#
+ prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_25/a_230_79# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_27/a_696_458#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_65/a_696_458# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_33/a_735_102#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_71/a_735_102# prbs_generator_syn_3/m3_13600_7263#
+ prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_43/a_222_392# prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_50/Y
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_8/a_1178_124# prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_53/B
+ prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_19/a_376_368# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_63/a_1178_124#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_4/a_696_458# prbs_generator_syn_3/sky130_fd_sc_hs__nor2b_1_4/a_278_368#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_13/a_1178_124# prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_61/a_132_392#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_53/a_206_368# prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_21/a_52_123#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_45/a_651_503# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_17/a_696_458#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_47/a_544_485# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_55/a_696_458#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_21/a_735_102# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_37/a_27_74#
+ prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_61/B prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_61/X
+ prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_59/a_112_119# prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_31/A
+ prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_33/a_222_392# prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_29/a_230_79#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_45/a_1226_296# prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_9/a_132_392#
+ prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_5/A prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_57/Y
+ prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_31/X prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_51/a_27_74#
+ prbs_generator_syn_3/sky130_fd_sc_hs__nor2b_1_8/a_27_112# prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_47/a_376_368#
+ prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_53/a_293_74# prbs_generator_syn_3/sky130_fd_sc_hs__nand2_1_43/a_117_74#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_8/a_735_102# prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_21/a_293_74#
+ prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_39/a_138_385# prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_63/Y
+ prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_51/a_132_392# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_43/a_206_368#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_53/a_437_503# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_37/a_544_485#
+ prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_57/X prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_53/a_1034_424#
+ prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_25/a_52_123# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_33/a_1141_508#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_63/Q prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_23/a_222_392#
+ prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_63/a_222_392# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_7/a_1178_124#
+ prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_53/X prbs_generator_syn_3/sky130_fd_sc_hs__nand2_2_5/Y
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_61/a_1178_124# prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_1/a_230_79#
+ prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_43/a_230_79# prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_11/a_230_79#
+ prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_41/a_132_392# prbs_generator_syn_3/sky130_fd_sc_hs__nand2_1_13/a_117_74#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_43/a_437_503# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_27/a_544_485#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_63/a_651_503# prbs_generator_syn_3/sky130_fd_sc_hs__nand2_1_7/a_117_74#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_35/a_696_458# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_65/a_544_485#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_51/a_1034_424# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_41/a_735_102#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_32/a_1141_508# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_49/a_1141_508#
+ prbs_generator_syn_3/sky130_fd_sc_hs__nand2_1_55/B prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_53/a_222_392#
+ prbs_generator_syn_3/sky130_fd_sc_hs__sdlclkp_2_1/a_114_112# prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_9/a_293_74#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_43/a_1226_296# prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_29/a_52_123#
+ prbs_generator_syn_3/sky130_fd_sc_hs__nand2_1_37/B prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_1/a_651_503#
+ prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_27/a_376_368# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_4/a_544_485#
+ prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_67/a_376_368# prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_27/X
+ prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_1/X prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_59/a_138_385#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_29/a_1178_124# prbs_generator_syn_3/m3_13600_2871#
+ prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_5/a_230_79# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_23/a_206_368#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_61/a_206_368# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_17/a_544_485#
+ prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_15/a_230_79# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_25/a_696_458#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_55/a_544_485# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_32/a_735_102#
+ prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_29/a_293_74# prbs_generator_syn_3/sky130_fd_sc_hs__nand2_1_17/a_117_74#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_69/a_1034_424# prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_29/a_112_119#
+ prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_37/X prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_31/B
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_19/a_1034_424# prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_33/A
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_9/a_206_368# prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_57/a_376_368#
+ prbs_generator_syn_3/sky130_fd_sc_hs__sdlclkp_2_1/a_706_317# prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_11/B
+ prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_1/a_52_123# prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_39/B
+ prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_21/a_132_392# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_13/a_206_368#
+ prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_43/a_52_123# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_51/a_206_368#
+ prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_47/X prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_23/a_437_503#
+ prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_11/a_52_123# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_61/a_437_503#
+ prbs_generator_syn_3/sky130_fd_sc_hs__nor2b_1_7/Y prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_51/A
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_15/a_696_458# prbs_generator_syn_3/sky130_fd_sc_hs__nor2b_1_5/Y
+ prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_9/a_230_79# prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_25/X
+ prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_19/a_112_119# prbs_generator_syn_3/sky130_fd_sc_hs__nand2_1_45/B
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_5/a_1178_124# prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_19/a_230_79#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_41/a_1226_296# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_59/a_1226_296#
+ prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_63/a_230_79# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_51/Q
+ prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_7/a_132_392# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_9/a_437_503#
+ prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_46/a_376_368# prbs_generator_syn_3/sky130_fd_sc_hs__nand2_1_33/a_117_74#
+ prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_11/a_293_74# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_27/a_1178_124#
+ prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_11/a_132_392# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_13/a_437_503#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_51/a_437_503# prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_5/a_52_123#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_35/a_544_485# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_73/a_651_503#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_45/a_696_458# prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_15/a_52_123#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_47/a_1141_508# prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_47/a_112_119#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_4/a_1178_124# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_17/a_1034_424#
+ prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_23/B prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_37/a_376_368#
+ prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_15/B prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_7/Y
+ prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_29/a_138_385# prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_33/a_230_79#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_25/a_1178_124# prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_47/a_293_74#
+ prbs_generator_syn_3/sky130_fd_sc_hs__nand2_1_37/a_117_74# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_33/a_206_368#
+ prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_15/a_293_74# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_71/a_206_368#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_25/a_544_485# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_67/a_1034_424#
+ prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_13/a_222_392# prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_9/a_52_123#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_15/a_1034_424# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_57/a_1226_296#
+ prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_19/a_52_123# prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_23/X
+ prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_63/a_52_123# prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_19/a_138_385#
+ prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_9/a_376_368# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_21/a_206_368#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_33/a_437_503# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_71/a_437_503#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_53/a_651_503# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_15/a_544_485#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_63/a_696_458# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_65/a_1034_424#
+ prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_19/a_293_74# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_45/a_1141_508#
+ prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_27/a_112_119# prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_67/a_112_119#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_1/a_1178_124# prbs_generator_syn_3/sky130_fd_sc_hs__conb_1_1/a_21_290#
+ prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_63/a_293_74# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_8/a_206_368#
+ prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_17/a_376_368# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_63/a_27_74#
+ prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_21/A prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_55/a_376_368#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_1/a_696_458# prbs_generator_syn_3/sky130_fd_sc_hs__nor2b_1_1/a_278_368#
+ prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_47/a_138_385# prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_33/a_52_123#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_9/a_1034_424# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_21/a_437_503#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_1/a_27_74# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_43/a_651_503#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_1/Q prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_45/a_544_485#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_69/a_735_102# prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_57/a_112_119#
+ prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_31/a_222_392# prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_13/A
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_55/a_1226_296# prbs_generator_syn_3/sky130_fd_sc_hs__nand2_2_5/a_27_74#
+ prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_53/a_230_79# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_8/a_437_503#
+ prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_67/a_293_74# prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_33/a_293_74#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_7/a_735_102# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_23/a_1178_124#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_41/a_206_368# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_8/a_1034_424#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_63/a_1034_424# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_59/a_735_102#
+ prbs_generator_syn_3/sky130_fd_sc_hs__nand2_1_5/B prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_43/a_1141_508#
+ prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_46/a_112_119# prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_61/a_222_392#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_13/a_1034_424# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_73/a_1178_124#
+ prbs_generator_syn_3/sky130_fd_sc_hs__nand2_1_27/B prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_13/B
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_57/a_27_74# prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_57/a_230_79#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_21/a_1178_124# prbs_generator_syn_3/sky130_fd_sc_hs__nor2b_1_1/a_27_112#
+ prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_27/a_138_385# prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_23/a_230_79#
+ prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_67/a_138_385# prbs_generator_syn_3/sky130_fd_sc_hs__nand2_1_41/B
+ prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_9/a_222_392# prbs_generator_syn_3/sky130_fd_sc_hs__nand2_1_27/a_117_74#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_32/a_206_368# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_23/a_651_503#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_41/a_437_503# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_73/a_27_74#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_61/a_651_503# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_63/a_544_485#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_49/a_735_102# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_73/a_696_458#
+ prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_37/a_112_119# prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_51/a_222_392#
+ prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_43/X prbs_generator_syn_3/sky130_fd_sc_hs__nand2_2_1/B
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_9/a_651_503# prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_53/a_52_123#
+ prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_49/X prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_25/a_376_368#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_1/a_544_485# prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_65/a_376_368#
+ prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_57/a_138_385# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_27/a_27_74#
+ prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_39/a_132_392# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_7/a_1034_424#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_13/a_651_503# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_32/a_437_503#
+ prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_27/a_230_79# prbs_generator_syn_3/m3_13600_12265#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_51/a_651_503# prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_59/B
+ prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_47/A prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_61/a_1034_424#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_41/a_1141_508# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_59/a_1141_508#
+ prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_41/a_222_392# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_53/a_1226_296#
+ prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_3/A prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_71/a_1178_124#
+ prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_9/a_112_119# prbs_generator_syn_3/sky130_fd_sc_hs__nand2_1_3/a_117_74#
+ prbs_generator_syn_3/m3_13600_8483# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_39/a_1178_124#
+ prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_57/a_52_123# prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_46/a_138_385#
+ prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_23/a_52_123# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_67/a_27_74#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_53/a_696_458# prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_17/a_112_119#
+ prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_11/A prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_55/a_112_119#
+ prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_1/A prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_51/a_1226_296#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_29/a_1034_424# prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_59/A
+ prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_23/A prbs_generator_syn_3/sky130_fd_sc_hs__nand2_1_39/B
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_5/a_27_74# prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_57/a_293_74#
+ prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_37/a_138_385# prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_59/a_132_392#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_33/a_651_503# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_71/a_651_503#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_43/a_696_458# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_73/a_544_485#
+ prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_27/a_52_123# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_57/a_1141_508#
+ prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_21/a_222_392# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_35/a_27_74#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_69/a_1226_296# prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_37/B
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_19/a_1226_296# prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_35/a_376_368#
+ prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_47/a_230_79# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_37/a_1178_124#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_5/a_1034_424# prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_49/a_132_392#
+ prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_7/a_222_392# prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_27/a_293_74#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_21/a_651_503# prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_9/a_138_385#
+ prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_11/a_222_392# prbs_generator_syn_3/m3_13600_14095#
+ prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_50/A prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_27/a_1034_424#
+ prbs_generator_syn_3/sky130_fd_sc_hs__nand2_1_13/B prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_8/a_651_503#
+ prbs_generator_syn_3/m3_13600_9703# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_35/a_1178_124#
+ prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_17/a_138_385# prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_55/a_138_385#
+ prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_7/a_230_79# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_4/a_1034_424#
+ prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_7/a_376_368# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_69/a_206_368#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_23/a_696_458# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_53/a_544_485#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_39/a_735_102# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_61/a_696_458#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_55/a_1141_508# prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_25/a_112_119#
+ prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_65/a_112_119# prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_43/a_293_74#
+ prbs_generator_syn_3/sky130_fd_sc_hs__nand2_1_57/B prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_25/a_1034_424#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_7/a_206_368# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_17/a_1226_296#
+ prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_15/a_376_368# prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_53/a_376_368#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_9/a_696_458# prbs_generator_syn_3/m3_13600_431#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_45/a_27_74# prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_47/a_52_123#
+ prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_29/a_132_392# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_59/a_206_368#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_69/a_437_503# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_41/a_651_503#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_43/a_544_485# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_13/a_696_458#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_29/a_735_102# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_51/a_696_458#
+ prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_61/Y prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_67/a_1226_296#
+ prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_5/a_132_392# prbs_generator_syn_3/sky130_fd_sc_hs__and2b_2_1/a_198_48#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_7/a_437_503# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_15/a_1226_296#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_69/a_27_74# prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_46/a_293_74#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_1/a_1034_424# prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_19/a_132_392#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_49/a_206_368# prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_7/a_52_123#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_59/a_437_503# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_32/a_651_503#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_7/a_27_74# prbs_generator_syn_3/sky130_fd_sc_hs__nand2_2_1/a_27_74#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_19/a_735_102# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_57/a_735_102#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_65/a_1226_296# prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_37/A
+ prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_33/a_376_368# prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_37/a_230_79#
+ prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_25/a_138_385# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_39/a_27_74#
+ prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_65/a_138_385# prbs_generator_syn_3/sky130_fd_sc_hs__nor2b_1_9/a_278_368#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_49/a_437_503# prbs_generator_syn_3/sky130_fd_sc_hs__and2b_2_1/a_505_74#
+ prbs_generator_syn_3/sky130_fd_sc_hs__nand2_1_51/a_117_74# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_23/a_544_485#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_33/a_696_458# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_61/a_544_485#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_9/a_1226_296# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_53/a_1141_508#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_71/a_696_458# prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_35/a_112_119#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_23/a_1034_424# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_9/a_544_485#
+ prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_63/a_376_368# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_33/a_1178_124#
+ prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_5/a_376_368# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_13/a_544_485#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_73/a_1034_424# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_21/a_696_458#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_51/a_544_485# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_8/a_1226_296#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_51/a_1141_508# prbs_generator_syn_3/sky130_fd_sc_hs__nand2_1_55/a_117_74#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_21/a_1034_424# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_63/a_1226_296#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_23/a_27_74# prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_7/a_112_119#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_13/a_1226_296# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_8/a_696_458#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_32/a_1178_124# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_49/a_1178_124#
+ prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_37/a_52_123# prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_27/a_132_392#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_71/Q prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_67/a_735_102#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_69/a_1141_508# prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_15/a_112_119#
+ prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_53/a_112_119# prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_39/a_222_392#
+ prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_55/a_230_79# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_19/a_1141_508#
+ prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_37/a_293_74# prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_43/a_376_368#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_5/a_735_102# prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_35/a_138_385#
+ prbs_generator_syn_3/sky130_fd_sc_hs__sdlclkp_2_1/a_114_424# prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_57/a_132_392#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_71/a_1034_424# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_7/a_1226_296#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_33/a_544_485# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_41/a_696_458#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_71/a_544_485# prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_21/B
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_61/a_1226_296# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_39/a_1034_424#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_17/a_27_74# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_9/a_27_74#
+ prbs_generator_syn_3/sky130_fd_sc_hs__nor2b_1_5/a_27_112# prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_47/a_132_392#
+ prbs_generator_syn_3/sky130_fd_sc_hs__nor2b_1_8/a_278_368# prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_9/B
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_39/a_206_368# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_33/a_27_74#
+ prbs_generator_syn_3/sky130_fd_sc_hs__nand2_1_41/a_117_74# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_69/a_651_503#
+ prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_51/a_293_74# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_21/a_544_485#
+ prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_7/a_138_385# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_32/a_696_458#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_47/a_735_102# prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_33/a_112_119#
+ prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_59/a_222_392# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_17/a_1141_508#
+ prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_55/a_52_123# prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_3/a_293_74#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_7/a_651_503# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_29/a_1226_296#
+ prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_23/a_376_368# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_8/a_544_485#
+ prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_47/B prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_47/a_1178_124#
+ prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_15/a_138_385# prbs_generator_syn_3/sky130_fd_sc_hs__sdlclkp_2_1/a_1195_374#
+ prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_53/a_138_385# prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_37/a_132_392#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_29/a_206_368# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_39/a_437_503#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_59/a_651_503# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_37/a_735_102#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_67/a_1141_508# prbs_generator_syn_3/sky130_fd_sc_hs__and2b_2_1/a_27_74#
+ prbs_generator_syn_3/sky130_fd_sc_hs__conb_1_1/a_165_290# prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_55/a_293_74#
+ prbs_generator_syn_3/sky130_fd_sc_hs__nand2_1_45/a_117_74# prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_63/a_112_119#
+ prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_49/a_222_392# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_37/a_1034_424#
+ prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_23/a_293_74# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_15/a_1141_508#
+ prbs_generator_syn_3/sky130_fd_sc_hs__nand2_1_5/a_117_74# prbs_generator_syn_3/m3_13600_13485#
+ prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_5/a_112_119# prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_13/a_376_368#
+ prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_51/a_376_368# prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_7/a_293_74#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_19/a_206_368# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_57/a_206_368#
+ prbs_generator_syn_3/sky130_fd_sc_hs__sdlclkp_2_1/a_318_74# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_29/a_437_503#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_49/a_651_503# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_25/a_27_74#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_5/a_1226_296# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_41/a_544_485#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_27/a_735_102# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_65/a_1141_508#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_65/a_735_102# prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_3/a_230_79#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_35/a_1034_424# prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_13/a_230_79#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_41/a_27_74# prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_3/a_132_392#
+ prbs_generator_syn_3/sky130_fd_sc_hs__nand2_1_49/a_117_74# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_27/a_1226_296#
+ prbs_generator_syn_3/sky130_fd_sc_hs__nand2_1_15/a_117_74# prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_41/a_376_368#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_45/a_1178_124# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_4/a_735_102#
+ prbs_generator_syn_3/sky130_fd_sc_hs__nand2_1_9/a_117_74# prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_33/a_138_385#
+ prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_17/a_132_392# prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_55/a_132_392#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_9/a_1141_508# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_19/a_437_503#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_57/a_437_503# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_4/a_1226_296#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_32/a_544_485# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_17/a_735_102#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_55/a_735_102# prbs_generator_syn_3/m3_13600_2261#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_65/a_27_74# prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_29/a_222_392#
+ prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_43/a_112_119# prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_19/X
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_25/a_1226_296# prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_31/a_376_368#
+ prbs_generator_syn_3/sky130_fd_sc_hs__or2_1_1/a_63_368# prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_17/a_230_79#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_4/a_27_74# prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_61/a_230_79#
+ prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_63/a_138_385# prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_5/a_222_392#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_8/a_1141_508# prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_41/a_293_74#
+ prbs_generator_syn_3/sky130_fd_sc_hs__nand2_1_31/a_117_74# prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_5/a_138_385#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_63/a_1141_508# prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_19/a_222_392#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_13/a_1141_508# prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_3/a_52_123#
+ prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_13/a_52_123# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_43/a_1178_124#
+ prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_61/a_376_368# prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_35/a_132_392#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_67/a_206_368# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_1/a_1226_296#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_69/a_696_458# prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_31/a_230_79#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_35/a_735_102# prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_23/a_112_119#
+ prbs_generator_syn_3/sky130_fd_sc_hs__nand2_1_35/a_117_74# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_59/a_27_74#
+ prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_13/a_293_74# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_5/a_206_368#
+ prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_50/a_376_368# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_7/a_696_458#
+ prbs_generator_syn_3/sky130_fd_sc_hs__nor2b_1_7/a_278_368# prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_17/a_52_123#
+ prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_43/a_138_385# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_7/a_1141_508#
+ prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_61/a_52_123# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_67/a_437_503#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_61/a_1141_508# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_25/a_735_102#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_59/a_696_458# prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_13/a_112_119#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_33/a_1034_424# prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_51/a_112_119#
+ prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_35/a_230_79# prbs_generator_syn_3/m3_13600_4091#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_23/a_1226_296# prbs_generator_syn_3/sky130_fd_sc_hs__nand2_1_39/a_117_74#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_29/a_27_74# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_5/a_437_503#
+ prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_17/a_293_74# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_41/a_1178_124#
+ prbs_generator_syn_3/sky130_fd_sc_hs__or2_1_1/a_152_368# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_59/a_1178_124#
+ prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_61/a_293_74# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_47/a_206_368#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_39/a_651_503# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_49/a_696_458#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_15/a_735_102# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_32/a_1034_424#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_73/a_1226_296# prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_27/a_222_392#
+ prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_41/a_112_119# prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_31/a_52_123#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_49/a_1034_424# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_29/a_1141_508#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_21/a_1226_296# prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_39/a_230_79#
+ prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_23/a_138_385# prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_51/a_230_79#
+ prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_45/a_132_392# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_37/a_206_368#
+ prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_65/a_293_74# prbs_generator_syn_3/sky130_fd_sc_hs__nand2_1_53/a_117_74#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_47/a_437_503# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_29/a_651_503#
+ prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_31/a_293_74# prbs_generator_syn_3/sky130_fd_sc_hs__nand2_1_21/a_117_74#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_69/a_544_485# prbs_generator_syn_3/sky130_fd_sc_hs__clkbuf_16_1/a_114_74#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_45/a_735_102# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_13/a_27_74#
+ prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_31/a_112_119# prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_57/a_222_392#
+ prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_35/a_52_123# prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_21/a_376_368#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_7/a_544_485# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_57/a_1178_124#
+ prbs_generator_syn_3/m3_13600_6043# prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_13/a_138_385#
+ prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_51/a_138_385# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_5/a_1141_508#
+ prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_3/a_376_368# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_27/a_206_368#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_65/a_206_368# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_37/a_437_503#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_19/a_651_503# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_57/a_651_503#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_59/a_544_485# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_71/a_1226_296#
+ prbs_generator_syn_3/sky130_fd_sc_hs__nand2_1_25/a_117_74# prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_61/a_112_119#
+ prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_47/a_222_392# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_27/a_1141_508#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_53/a_27_74# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_4/a_206_368#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_39/a_1226_296# prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_11/a_376_368#
+ prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_39/a_52_123# prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_41/a_138_385#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_4/a_1141_508# prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_25/a_132_392#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_17/a_206_368# prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_41/A
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_55/a_206_368# prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_51/a_52_123#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_27/a_437_503# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_65/a_437_503#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_49/a_544_485# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_63/a_735_102#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_47/a_1034_424# prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_50/a_112_119#
+ prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_37/a_222_392# prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_59/a_230_79#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_25/a_1141_508# prbs_generator_syn_3/sky130_fd_sc_hs__nor2b_1_4/a_27_112#
+ prbs_generator_syn_3/sky130_fd_sc_hs__sdlclkp_2_1/a_685_81# prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_1/a_132_392#
+ prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_39/a_293_74# prbs_generator_syn_3/sky130_fd_sc_hs__nand2_1_29/a_117_74#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_4/a_437_503# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_55/a_1178_124#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_21/a_27_74# prbs_generator_syn_3/m3_13600_12875#
+ prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_50/a_293_74# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_1/a_735_102#
+ prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_31/a_138_385# prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_15/a_132_392#
+ prbs_generator_syn_3/sky130_fd_sc_hs__nand2_1_1/a_117_74# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_17/a_437_503#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_55/a_437_503# prbs_generator_syn
Xsky130_fd_sc_hs__clkdlyinv5sd2_1_1 DVSS: DVDD: DVSS: DVDD: dout_p sky130_fd_sc_hs__nand2_2_1/B
+ sky130_fd_sc_hs__clkdlyinv5sd2_1_1/a_28_74# sky130_fd_sc_hs__clkdlyinv5sd2_1_1/a_682_74#
+ sky130_fd_sc_hs__clkdlyinv5sd2_1_1/a_549_74# sky130_fd_sc_hs__clkdlyinv5sd2_1_1/a_288_74#
+ sky130_fd_sc_hs__clkdlyinv5sd2_1
Xsky130_fd_sc_hs__o21bai_2_9 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__nand2_2_7/A
+ sky130_fd_sc_hs__o21bai_4_7/A1 sky130_fd_sc_hs__dlrtp_1_65/D sky130_fd_sc_hs__buf_2_57/A
+ sky130_fd_sc_hs__o21bai_2_9/a_27_74# sky130_fd_sc_hs__o21bai_2_9/a_225_74# sky130_fd_sc_hs__o21bai_2_9/a_507_368#
+ sky130_fd_sc_hs__o21bai_2
Xsky130_fd_sc_hs__o21ai_2_14 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__inv_4_17/Y sky130_fd_sc_hs__o21ai_2_55/A1
+ sky130_fd_sc_hs__nand2_2_7/A sky130_fd_sc_hs__o21ai_2_15/Y sky130_fd_sc_hs__o21ai_2_15/a_116_368#
+ sky130_fd_sc_hs__o21ai_2_15/a_27_74# sky130_fd_sc_hs__o21ai_2
Xsky130_fd_sc_hs__o21ai_2_25 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__inv_4_15/Y sky130_fd_sc_hs__nand2_2_11/B
+ sky130_fd_sc_hs__o21ai_2_55/A1 sky130_fd_sc_hs__o21ai_2_25/Y sky130_fd_sc_hs__o21ai_2_25/a_116_368#
+ sky130_fd_sc_hs__o21ai_2_25/a_27_74# sky130_fd_sc_hs__o21ai_2
Xsky130_fd_sc_hs__o21ai_2_36 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__inv_4_23/Y sky130_fd_sc_hs__or2b_4_1/A
+ sky130_fd_sc_hs__nand2_2_15/B sky130_fd_sc_hs__o21ai_2_37/Y sky130_fd_sc_hs__o21ai_2_37/a_116_368#
+ sky130_fd_sc_hs__o21ai_2_37/a_27_74# sky130_fd_sc_hs__o21ai_2
Xsky130_fd_sc_hs__o21ai_2_47 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__nand2_2_27/B
+ sky130_fd_sc_hs__nand2_2_21/B sky130_fd_sc_hs__clkinv_4_7/Y sky130_fd_sc_hs__o21ai_2_47/Y
+ sky130_fd_sc_hs__o21ai_2_47/a_116_368# sky130_fd_sc_hs__o21ai_2_47/a_27_74# sky130_fd_sc_hs__o21ai_2
Xsky130_fd_sc_hs__clkinv_4_17 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__nor2_4_3/B
+ sky130_fd_sc_hs__nand2_2_7/A sky130_fd_sc_hs__clkinv_4
Xprbs_generator_syn_19 prbs_generator_syn_19/clk prbs_generator_syn_19/rst prbs_generator_syn_19/cke
+ sky130_fd_sc_hs__conb_1_209/LO sky130_fd_sc_hs__conb_1_209/LO sky130_fd_sc_hs__conb_1_209/HI
+ sky130_fd_sc_hs__conb_1_209/HI sky130_fd_sc_hs__conb_1_209/LO sky130_fd_sc_hs__conb_1_209/LO
+ sky130_fd_sc_hs__conb_1_209/LO sky130_fd_sc_hs__conb_1_209/HI sky130_fd_sc_hs__conb_1_209/HI
+ sky130_fd_sc_hs__conb_1_209/HI sky130_fd_sc_hs__conb_1_209/HI prbs_generator_syn_19/cke
+ prbs_generator_syn_19/eqn[31] prbs_generator_syn_19/cke prbs_generator_syn_19/eqn[31]
+ prbs_generator_syn_19/eqn[31] prbs_generator_syn_19/eqn[31] prbs_generator_syn_19/eqn[31]
+ prbs_generator_syn_19/eqn[2] prbs_generator_syn_19/eqn[2] prbs_generator_syn_19/eqn[2]
+ prbs_generator_syn_19/eqn[2] prbs_generator_syn_19/eqn[2] prbs_generator_syn_19/eqn[1]
+ sky130_fd_sc_hs__conb_1_203/HI sky130_fd_sc_hs__conb_1_203/HI sky130_fd_sc_hs__conb_1_203/HI
+ sky130_fd_sc_hs__conb_1_203/HI sky130_fd_sc_hs__conb_1_203/LO sky130_fd_sc_hs__conb_1_203/LO
+ sky130_fd_sc_hs__conb_1_203/HI sky130_fd_sc_hs__conb_1_203/HI prbs_generator_syn_19/eqn[31]
+ prbs_generator_syn_19/eqn[30] prbs_generator_syn_19/eqn[30] prbs_generator_syn_19/eqn[30]
+ prbs_generator_syn_19/eqn[30] prbs_generator_syn_19/eqn[30] prbs_generator_syn_19/eqn[30]
+ prbs_generator_syn_19/eqn[30] prbs_generator_syn_19/eqn[30] prbs_generator_syn_19/eqn[22]
+ prbs_generator_syn_19/eqn[22] prbs_generator_syn_19/eqn[20] prbs_generator_syn_19/eqn[22]
+ prbs_generator_syn_19/eqn[22] prbs_generator_syn_19/eqn[22] prbs_generator_syn_19/eqn[22]
+ prbs_generator_syn_19/eqn[22] prbs_generator_syn_19/eqn[22] prbs_generator_syn_19/eqn[13]
+ prbs_generator_syn_19/eqn[13] prbs_generator_syn_19/eqn[13] prbs_generator_syn_19/eqn[9]
+ prbs_generator_syn_19/eqn[9] prbs_generator_syn_19/eqn[9] prbs_generator_syn_19/eqn[9]
+ prbs_generator_syn_19/eqn[9] prbs_generator_syn_19/eqn[9] prbs_generator_syn_19/eqn[9]
+ prbs_generator_syn_19/eqn[9] prbs_generator_syn_19/eqn[2] prbs_generator_syn_19/eqn[1]
+ prbs_generator_syn_19/eqn[2] prbs_generator_syn_19/inj_err prbs_generator_syn_19/eqn[31]
+ prbs_generator_syn_19/eqn[31] prbs_generator_syn_19/out DVSS: DVDD: prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_1/a_293_74#
+ prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_15/X prbs_generator_syn_19/sky130_fd_sc_hs__nand2_1_35/B
+ prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_51/Y prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_9/A
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_9/CLK prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_47/a_27_74#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_37/a_1226_296# prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_3/B
+ prbs_generator_syn_19/sky130_fd_sc_hs__nor2b_1_7/a_27_112# prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_29/B
+ prbs_generator_syn_19/sky130_fd_sc_hs__sdlclkp_2_1/a_580_74# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_1/a_1141_508#
+ prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_5/Y prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_41/a_230_79#
+ prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_61/a_138_385# prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_43/a_132_392#
+ prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_3/a_222_392# prbs_generator_syn_19/sky130_fd_sc_hs__nor2b_1_9/a_27_112#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_61/a_27_74# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_35/a_206_368#
+ prbs_generator_syn_19/sky130_fd_sc_hs__nand2_2_3/Y prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_25/B
+ prbs_generator_syn_19/sky130_fd_sc_hs__nand2_1_11/a_117_74# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_67/a_651_503#
+ prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_45/X prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_39/a_696_458#
+ prbs_generator_syn_19/sky130_fd_sc_hs__sdlclkp_2_1/a_1198_74# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_45/a_1034_424#
+ prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_17/a_222_392# prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_55/a_222_392#
+ prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_53/Y prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_35/A
+ prbs_generator_syn_19/m3_13600_1651# prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_59/a_52_123#
+ prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_5/a_293_74# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_35/a_1226_296#
+ prbs_generator_syn_19/sky130_fd_sc_hs__nand2_1_51/B prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_5/a_651_503#
+ prbs_generator_syn_19/sky130_fd_sc_hs__nand2_1_21/B prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_8/a_27_74#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_15/a_27_74# prbs_generator_syn_19/sky130_fd_sc_hs__and2b_2_1/X
+ prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_13/X prbs_generator_syn_19/sky130_fd_sc_hs__nand2_2_3/a_27_74#
+ prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_50/a_138_385# prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_33/a_132_392#
+ prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_1/a_376_368# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_25/a_206_368#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_35/a_437_503# prbs_generator_syn_19/sky130_fd_sc_hs__sdlclkp_2_1/a_708_451#
+ prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_45/a_230_79# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_29/a_696_458#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_32/a_27_74# prbs_generator_syn_19/sky130_fd_sc_hs__nor2b_1_4/Y
+ prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_59/a_293_74# prbs_generator_syn_19/sky130_fd_sc_hs__nand2_1_47/a_117_74#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_73/a_735_102# prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_21/a_112_119#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_23/a_1141_508# prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_25/a_293_74#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_7/Q prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_3/a_112_119#
+ prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_35/B prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_51/X
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_53/a_1178_124# prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_23/a_132_392#
+ prbs_generator_syn_19/sky130_fd_sc_hs__nand2_1_3/B prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_15/a_206_368#
+ prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_63/a_132_392# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_55/a_27_74#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_25/a_437_503# prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_41/a_52_123#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_47/a_651_503# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_73/a_1141_508#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_19/a_696_458# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_57/a_696_458#
+ prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_7/X prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_43/a_1034_424#
+ prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_55/A prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_11/a_112_119#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_21/a_1141_508# prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_35/a_222_392#
+ prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_49/a_230_79# prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_67/Y
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_71/a_27_74# prbs_generator_syn_19/sky130_fd_sc_hs__nand2_1_33/B
+ prbs_generator_syn_19/sky130_fd_sc_hs__conb_1_1/LO prbs_generator_syn_19/sky130_fd_sc_hs__nand2_1_19/a_117_74#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_51/a_1178_124# prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_33/X
+ prbs_generator_syn_19/sky130_fd_sc_hs__nand2_1_29/B prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_41/Y
+ prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_53/a_132_392# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_45/a_206_368#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_15/a_437_503# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_37/a_651_503#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_39/a_544_485# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_53/a_735_102#
+ prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_45/a_52_123# prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_1/B
+ prbs_generator_syn_19/sky130_fd_sc_hs__nand2_2_3/B prbs_generator_syn_19/sky130_fd_sc_hs__clkbuf_16_1/A
+ prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_21/X prbs_generator_syn_19/sky130_fd_sc_hs__nand2_1_25/B
+ prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_39/a_376_368# prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_63/X
+ prbs_generator_syn_19/m3_13600_3481# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_69/a_1178_124#
+ prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_21/a_138_385# prbs_generator_syn_19/sky130_fd_sc_hs__nor2b_1_8/Y
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_19/a_1178_124# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_49/a_27_74#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_45/a_437_503# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_27/a_651_503#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_71/a_1141_508# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_65/a_651_503#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_29/a_544_485# prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_3/a_138_385#
+ prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_55/X prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_43/a_735_102#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_41/a_1034_424# prbs_generator_syn_19/sky130_fd_sc_hs__nand2_1_9/B
+ prbs_generator_syn_19/sky130_fd_sc_hs__nor2b_1_9/Y prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_59/a_1034_424#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_39/a_1141_508# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_33/a_1226_296#
+ prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_49/a_52_123# prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_47/Y
+ prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_43/Y prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_4/a_651_503#
+ prbs_generator_syn_19/sky130_fd_sc_hs__nand2_1_49/B prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_19/A
+ prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_11/a_138_385# prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_5/X
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_63/a_206_368# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_17/a_651_503#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_19/a_544_485# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_55/a_651_503#
+ prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_9/Y prbs_generator_syn_19/sky130_fd_sc_hs__nand2_1_17/B
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_57/a_544_485# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_67/a_696_458#
+ prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_35/X prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_19/a_27_74#
+ prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_45/a_222_392# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_32/a_1226_296#
+ prbs_generator_syn_19/sky130_fd_sc_hs__nand2_1_43/B prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_25/A
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_1/a_206_368# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_49/a_1226_296#
+ prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_1/a_112_119# prbs_generator_syn_19/sky130_fd_sc_hs__or2_1_1/X
+ prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_59/a_376_368# prbs_generator_syn_19/sky130_fd_sc_hs__nand2_1_19/B
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_5/a_696_458# prbs_generator_syn_19/sky130_fd_sc_hs__nor2b_1_1/Y
+ prbs_generator_syn_19/sky130_fd_sc_hs__nor2b_1_5/a_278_368# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_17/a_1178_124#
+ prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_39/X prbs_generator_syn_19/m3_13600_5433#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_63/a_437_503# prbs_generator_syn_19/sky130_fd_sc_hs__nand2_2_5/B
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_23/a_735_102# prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_53/A
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_61/a_735_102# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_57/a_1034_424#
+ prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_63/B prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_37/a_1141_508#
+ prbs_generator_syn_19/sky130_fd_sc_hs__nand2_1_47/B prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_29/X
+ prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_65/Y prbs_generator_syn_19/m3_13600_4701#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_1/a_437_503# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_67/a_1178_124#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_9/a_735_102# prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_13/a_132_392#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_15/a_1178_124# prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_15/A
+ prbs_generator_syn_19/sky130_fd_sc_hs__nand2_1_1/B prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_43/B
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_35/a_651_503# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_8/D
+ prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_29/A prbs_generator_syn_19/sky130_fd_sc_hs__nand2_1_7/B
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_13/a_735_102# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_47/a_696_458#
+ prbs_generator_syn_19/sky130_fd_sc_hs__nand2_1_31/B prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_51/a_735_102#
+ prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_59/X prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_35/a_1141_508#
+ prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_25/a_222_392# prbs_generator_syn_19/sky130_fd_sc_hs__sdlclkp_2_1/a_288_48#
+ prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_55/B prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_17/B
+ prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_43/A prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_7/A
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_65/a_1178_124# prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_59/Y
+ prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_41/X prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_21/a_230_79#
+ prbs_generator_syn_19/sky130_fd_sc_hs__nand2_1_57/a_117_74# prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_1/a_222_392#
+ prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_19/B prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_35/a_293_74#
+ prbs_generator_syn_19/sky130_fd_sc_hs__nand2_1_23/a_117_74# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_73/a_206_368#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_25/a_651_503# prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_1/a_138_385#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_37/a_696_458# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_67/a_544_485#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_43/a_27_74# prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_9/X
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_55/a_1034_424# prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_39/a_112_119#
+ prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_15/a_222_392# prbs_generator_syn_19/sky130_fd_sc_hs__conb_1_1/HI
+ prbs_generator_syn_19/sky130_fd_sc_hs__nand2_1_23/B prbs_generator_syn_19/sky130_fd_sc_hs__nand2_1_53/B
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_9/a_1178_124# prbs_generator_syn_19/sky130_fd_sc_hs__nor2b_1_4/A
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_47/a_1226_296# prbs_generator_syn_19/m3_13600_11045#
+ prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_17/X prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_29/a_376_368#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_5/a_544_485# prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_3/X
+ prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_31/a_132_392# prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_61/A
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_15/a_651_503# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_73/a_437_503#
+ prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_25/a_230_79# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_27/a_696_458#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_65/a_696_458# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_33/a_735_102#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_71/a_735_102# prbs_generator_syn_19/m3_13600_7263#
+ prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_43/a_222_392# prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_50/Y
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_8/a_1178_124# prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_53/B
+ prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_19/a_376_368# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_63/a_1178_124#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_4/a_696_458# prbs_generator_syn_19/sky130_fd_sc_hs__nor2b_1_4/a_278_368#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_13/a_1178_124# prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_61/a_132_392#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_53/a_206_368# prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_21/a_52_123#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_45/a_651_503# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_17/a_696_458#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_47/a_544_485# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_55/a_696_458#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_21/a_735_102# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_37/a_27_74#
+ prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_61/B prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_61/X
+ prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_59/a_112_119# prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_31/A
+ prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_33/a_222_392# prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_29/a_230_79#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_45/a_1226_296# prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_9/a_132_392#
+ prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_5/A prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_57/Y
+ prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_31/X prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_51/a_27_74#
+ prbs_generator_syn_19/sky130_fd_sc_hs__nor2b_1_8/a_27_112# prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_47/a_376_368#
+ prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_53/a_293_74# prbs_generator_syn_19/sky130_fd_sc_hs__nand2_1_43/a_117_74#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_8/a_735_102# prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_21/a_293_74#
+ prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_39/a_138_385# prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_63/Y
+ prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_51/a_132_392# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_43/a_206_368#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_53/a_437_503# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_37/a_544_485#
+ prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_57/X prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_53/a_1034_424#
+ prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_25/a_52_123# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_33/a_1141_508#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_63/Q prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_23/a_222_392#
+ prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_63/a_222_392# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_7/a_1178_124#
+ prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_53/X prbs_generator_syn_19/sky130_fd_sc_hs__nand2_2_5/Y
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_61/a_1178_124# prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_1/a_230_79#
+ prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_43/a_230_79# prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_11/a_230_79#
+ prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_41/a_132_392# prbs_generator_syn_19/sky130_fd_sc_hs__nand2_1_13/a_117_74#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_43/a_437_503# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_27/a_544_485#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_63/a_651_503# prbs_generator_syn_19/sky130_fd_sc_hs__nand2_1_7/a_117_74#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_35/a_696_458# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_65/a_544_485#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_51/a_1034_424# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_41/a_735_102#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_32/a_1141_508# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_49/a_1141_508#
+ prbs_generator_syn_19/sky130_fd_sc_hs__nand2_1_55/B prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_53/a_222_392#
+ prbs_generator_syn_19/sky130_fd_sc_hs__sdlclkp_2_1/a_114_112# prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_9/a_293_74#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_43/a_1226_296# prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_29/a_52_123#
+ prbs_generator_syn_19/sky130_fd_sc_hs__nand2_1_37/B prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_1/a_651_503#
+ prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_27/a_376_368# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_4/a_544_485#
+ prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_67/a_376_368# prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_27/X
+ prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_1/X prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_59/a_138_385#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_29/a_1178_124# prbs_generator_syn_19/m3_13600_2871#
+ prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_5/a_230_79# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_23/a_206_368#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_61/a_206_368# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_17/a_544_485#
+ prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_15/a_230_79# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_25/a_696_458#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_55/a_544_485# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_32/a_735_102#
+ prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_29/a_293_74# prbs_generator_syn_19/sky130_fd_sc_hs__nand2_1_17/a_117_74#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_69/a_1034_424# prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_29/a_112_119#
+ prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_37/X prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_31/B
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_19/a_1034_424# prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_33/A
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_9/a_206_368# prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_57/a_376_368#
+ prbs_generator_syn_19/sky130_fd_sc_hs__sdlclkp_2_1/a_706_317# prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_11/B
+ prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_1/a_52_123# prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_39/B
+ prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_21/a_132_392# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_13/a_206_368#
+ prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_43/a_52_123# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_51/a_206_368#
+ prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_47/X prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_23/a_437_503#
+ prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_11/a_52_123# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_61/a_437_503#
+ prbs_generator_syn_19/sky130_fd_sc_hs__nor2b_1_7/Y prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_51/A
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_15/a_696_458# prbs_generator_syn_19/sky130_fd_sc_hs__nor2b_1_5/Y
+ prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_9/a_230_79# prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_25/X
+ prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_19/a_112_119# prbs_generator_syn_19/sky130_fd_sc_hs__nand2_1_45/B
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_5/a_1178_124# prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_19/a_230_79#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_41/a_1226_296# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_59/a_1226_296#
+ prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_63/a_230_79# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_51/Q
+ prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_7/a_132_392# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_9/a_437_503#
+ prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_46/a_376_368# prbs_generator_syn_19/sky130_fd_sc_hs__nand2_1_33/a_117_74#
+ prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_11/a_293_74# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_27/a_1178_124#
+ prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_11/a_132_392# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_13/a_437_503#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_51/a_437_503# prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_5/a_52_123#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_35/a_544_485# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_73/a_651_503#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_45/a_696_458# prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_15/a_52_123#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_47/a_1141_508# prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_47/a_112_119#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_4/a_1178_124# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_17/a_1034_424#
+ prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_23/B prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_37/a_376_368#
+ prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_15/B prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_7/Y
+ prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_29/a_138_385# prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_33/a_230_79#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_25/a_1178_124# prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_47/a_293_74#
+ prbs_generator_syn_19/sky130_fd_sc_hs__nand2_1_37/a_117_74# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_33/a_206_368#
+ prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_15/a_293_74# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_71/a_206_368#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_25/a_544_485# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_67/a_1034_424#
+ prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_13/a_222_392# prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_9/a_52_123#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_15/a_1034_424# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_57/a_1226_296#
+ prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_19/a_52_123# prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_23/X
+ prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_63/a_52_123# prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_19/a_138_385#
+ prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_9/a_376_368# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_21/a_206_368#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_33/a_437_503# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_71/a_437_503#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_53/a_651_503# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_15/a_544_485#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_63/a_696_458# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_65/a_1034_424#
+ prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_19/a_293_74# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_45/a_1141_508#
+ prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_27/a_112_119# prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_67/a_112_119#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_1/a_1178_124# prbs_generator_syn_19/sky130_fd_sc_hs__conb_1_1/a_21_290#
+ prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_63/a_293_74# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_8/a_206_368#
+ prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_17/a_376_368# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_63/a_27_74#
+ prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_21/A prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_55/a_376_368#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_1/a_696_458# prbs_generator_syn_19/sky130_fd_sc_hs__nor2b_1_1/a_278_368#
+ prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_47/a_138_385# prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_33/a_52_123#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_9/a_1034_424# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_21/a_437_503#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_1/a_27_74# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_43/a_651_503#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_1/Q prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_45/a_544_485#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_69/a_735_102# prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_57/a_112_119#
+ prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_31/a_222_392# prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_13/A
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_55/a_1226_296# prbs_generator_syn_19/sky130_fd_sc_hs__nand2_2_5/a_27_74#
+ prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_53/a_230_79# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_8/a_437_503#
+ prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_67/a_293_74# prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_33/a_293_74#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_7/a_735_102# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_23/a_1178_124#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_41/a_206_368# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_8/a_1034_424#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_63/a_1034_424# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_59/a_735_102#
+ prbs_generator_syn_19/sky130_fd_sc_hs__nand2_1_5/B prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_43/a_1141_508#
+ prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_46/a_112_119# prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_61/a_222_392#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_13/a_1034_424# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_73/a_1178_124#
+ prbs_generator_syn_19/sky130_fd_sc_hs__nand2_1_27/B prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_13/B
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_57/a_27_74# prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_57/a_230_79#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_21/a_1178_124# prbs_generator_syn_19/sky130_fd_sc_hs__nor2b_1_1/a_27_112#
+ prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_27/a_138_385# prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_23/a_230_79#
+ prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_67/a_138_385# prbs_generator_syn_19/sky130_fd_sc_hs__nand2_1_41/B
+ prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_9/a_222_392# prbs_generator_syn_19/sky130_fd_sc_hs__nand2_1_27/a_117_74#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_32/a_206_368# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_23/a_651_503#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_41/a_437_503# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_73/a_27_74#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_61/a_651_503# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_63/a_544_485#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_49/a_735_102# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_73/a_696_458#
+ prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_37/a_112_119# prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_51/a_222_392#
+ prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_43/X prbs_generator_syn_19/sky130_fd_sc_hs__nand2_2_1/B
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_9/a_651_503# prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_53/a_52_123#
+ prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_49/X prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_25/a_376_368#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_1/a_544_485# prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_65/a_376_368#
+ prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_57/a_138_385# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_27/a_27_74#
+ prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_39/a_132_392# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_7/a_1034_424#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_13/a_651_503# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_32/a_437_503#
+ prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_27/a_230_79# prbs_generator_syn_19/m3_13600_12265#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_51/a_651_503# prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_59/B
+ prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_47/A prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_61/a_1034_424#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_41/a_1141_508# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_59/a_1141_508#
+ prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_41/a_222_392# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_53/a_1226_296#
+ prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_3/A prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_71/a_1178_124#
+ prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_9/a_112_119# prbs_generator_syn_19/sky130_fd_sc_hs__nand2_1_3/a_117_74#
+ prbs_generator_syn_19/m3_13600_8483# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_39/a_1178_124#
+ prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_57/a_52_123# prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_46/a_138_385#
+ prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_23/a_52_123# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_67/a_27_74#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_53/a_696_458# prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_17/a_112_119#
+ prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_11/A prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_55/a_112_119#
+ prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_1/A prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_51/a_1226_296#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_29/a_1034_424# prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_59/A
+ prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_23/A prbs_generator_syn_19/sky130_fd_sc_hs__nand2_1_39/B
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_5/a_27_74# prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_57/a_293_74#
+ prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_37/a_138_385# prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_59/a_132_392#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_33/a_651_503# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_71/a_651_503#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_43/a_696_458# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_73/a_544_485#
+ prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_27/a_52_123# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_57/a_1141_508#
+ prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_21/a_222_392# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_35/a_27_74#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_69/a_1226_296# prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_37/B
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_19/a_1226_296# prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_35/a_376_368#
+ prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_47/a_230_79# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_37/a_1178_124#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_5/a_1034_424# prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_49/a_132_392#
+ prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_7/a_222_392# prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_27/a_293_74#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_21/a_651_503# prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_9/a_138_385#
+ prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_11/a_222_392# prbs_generator_syn_19/m3_13600_14095#
+ prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_50/A prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_27/a_1034_424#
+ prbs_generator_syn_19/sky130_fd_sc_hs__nand2_1_13/B prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_8/a_651_503#
+ prbs_generator_syn_19/m3_13600_9703# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_35/a_1178_124#
+ prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_17/a_138_385# prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_55/a_138_385#
+ prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_7/a_230_79# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_4/a_1034_424#
+ prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_7/a_376_368# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_69/a_206_368#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_23/a_696_458# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_53/a_544_485#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_39/a_735_102# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_61/a_696_458#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_55/a_1141_508# prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_25/a_112_119#
+ prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_65/a_112_119# prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_43/a_293_74#
+ prbs_generator_syn_19/sky130_fd_sc_hs__nand2_1_57/B prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_25/a_1034_424#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_7/a_206_368# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_17/a_1226_296#
+ prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_15/a_376_368# prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_53/a_376_368#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_9/a_696_458# prbs_generator_syn_19/m3_13600_431#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_45/a_27_74# prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_47/a_52_123#
+ prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_29/a_132_392# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_59/a_206_368#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_69/a_437_503# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_41/a_651_503#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_43/a_544_485# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_13/a_696_458#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_29/a_735_102# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_51/a_696_458#
+ prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_61/Y prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_67/a_1226_296#
+ prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_5/a_132_392# prbs_generator_syn_19/sky130_fd_sc_hs__and2b_2_1/a_198_48#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_7/a_437_503# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_15/a_1226_296#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_69/a_27_74# prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_46/a_293_74#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_1/a_1034_424# prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_19/a_132_392#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_49/a_206_368# prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_7/a_52_123#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_59/a_437_503# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_32/a_651_503#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_7/a_27_74# prbs_generator_syn_19/sky130_fd_sc_hs__nand2_2_1/a_27_74#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_19/a_735_102# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_57/a_735_102#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_65/a_1226_296# prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_37/A
+ prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_33/a_376_368# prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_37/a_230_79#
+ prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_25/a_138_385# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_39/a_27_74#
+ prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_65/a_138_385# prbs_generator_syn_19/sky130_fd_sc_hs__nor2b_1_9/a_278_368#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_49/a_437_503# prbs_generator_syn_19/sky130_fd_sc_hs__and2b_2_1/a_505_74#
+ prbs_generator_syn_19/sky130_fd_sc_hs__nand2_1_51/a_117_74# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_23/a_544_485#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_33/a_696_458# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_61/a_544_485#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_9/a_1226_296# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_53/a_1141_508#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_71/a_696_458# prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_35/a_112_119#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_23/a_1034_424# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_9/a_544_485#
+ prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_63/a_376_368# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_33/a_1178_124#
+ prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_5/a_376_368# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_13/a_544_485#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_73/a_1034_424# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_21/a_696_458#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_51/a_544_485# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_8/a_1226_296#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_51/a_1141_508# prbs_generator_syn_19/sky130_fd_sc_hs__nand2_1_55/a_117_74#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_21/a_1034_424# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_63/a_1226_296#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_23/a_27_74# prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_7/a_112_119#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_13/a_1226_296# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_8/a_696_458#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_32/a_1178_124# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_49/a_1178_124#
+ prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_37/a_52_123# prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_27/a_132_392#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_71/Q prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_67/a_735_102#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_69/a_1141_508# prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_15/a_112_119#
+ prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_53/a_112_119# prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_39/a_222_392#
+ prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_55/a_230_79# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_19/a_1141_508#
+ prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_37/a_293_74# prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_43/a_376_368#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_5/a_735_102# prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_35/a_138_385#
+ prbs_generator_syn_19/sky130_fd_sc_hs__sdlclkp_2_1/a_114_424# prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_57/a_132_392#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_71/a_1034_424# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_7/a_1226_296#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_33/a_544_485# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_41/a_696_458#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_71/a_544_485# prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_21/B
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_61/a_1226_296# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_39/a_1034_424#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_17/a_27_74# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_9/a_27_74#
+ prbs_generator_syn_19/sky130_fd_sc_hs__nor2b_1_5/a_27_112# prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_47/a_132_392#
+ prbs_generator_syn_19/sky130_fd_sc_hs__nor2b_1_8/a_278_368# prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_9/B
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_39/a_206_368# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_33/a_27_74#
+ prbs_generator_syn_19/sky130_fd_sc_hs__nand2_1_41/a_117_74# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_69/a_651_503#
+ prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_51/a_293_74# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_21/a_544_485#
+ prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_7/a_138_385# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_32/a_696_458#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_47/a_735_102# prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_33/a_112_119#
+ prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_59/a_222_392# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_17/a_1141_508#
+ prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_55/a_52_123# prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_3/a_293_74#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_7/a_651_503# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_29/a_1226_296#
+ prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_23/a_376_368# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_8/a_544_485#
+ prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_47/B prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_47/a_1178_124#
+ prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_15/a_138_385# prbs_generator_syn_19/sky130_fd_sc_hs__sdlclkp_2_1/a_1195_374#
+ prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_53/a_138_385# prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_37/a_132_392#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_29/a_206_368# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_39/a_437_503#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_59/a_651_503# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_37/a_735_102#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_67/a_1141_508# prbs_generator_syn_19/sky130_fd_sc_hs__and2b_2_1/a_27_74#
+ prbs_generator_syn_19/sky130_fd_sc_hs__conb_1_1/a_165_290# prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_55/a_293_74#
+ prbs_generator_syn_19/sky130_fd_sc_hs__nand2_1_45/a_117_74# prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_63/a_112_119#
+ prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_49/a_222_392# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_37/a_1034_424#
+ prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_23/a_293_74# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_15/a_1141_508#
+ prbs_generator_syn_19/sky130_fd_sc_hs__nand2_1_5/a_117_74# prbs_generator_syn_19/m3_13600_13485#
+ prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_5/a_112_119# prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_13/a_376_368#
+ prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_51/a_376_368# prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_7/a_293_74#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_19/a_206_368# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_57/a_206_368#
+ prbs_generator_syn_19/sky130_fd_sc_hs__sdlclkp_2_1/a_318_74# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_29/a_437_503#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_49/a_651_503# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_25/a_27_74#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_5/a_1226_296# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_41/a_544_485#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_27/a_735_102# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_65/a_1141_508#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_65/a_735_102# prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_3/a_230_79#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_35/a_1034_424# prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_13/a_230_79#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_41/a_27_74# prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_3/a_132_392#
+ prbs_generator_syn_19/sky130_fd_sc_hs__nand2_1_49/a_117_74# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_27/a_1226_296#
+ prbs_generator_syn_19/sky130_fd_sc_hs__nand2_1_15/a_117_74# prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_41/a_376_368#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_45/a_1178_124# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_4/a_735_102#
+ prbs_generator_syn_19/sky130_fd_sc_hs__nand2_1_9/a_117_74# prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_33/a_138_385#
+ prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_17/a_132_392# prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_55/a_132_392#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_9/a_1141_508# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_19/a_437_503#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_57/a_437_503# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_4/a_1226_296#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_32/a_544_485# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_17/a_735_102#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_55/a_735_102# prbs_generator_syn_19/m3_13600_2261#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_65/a_27_74# prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_29/a_222_392#
+ prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_43/a_112_119# prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_19/X
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_25/a_1226_296# prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_31/a_376_368#
+ prbs_generator_syn_19/sky130_fd_sc_hs__or2_1_1/a_63_368# prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_17/a_230_79#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_4/a_27_74# prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_61/a_230_79#
+ prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_63/a_138_385# prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_5/a_222_392#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_8/a_1141_508# prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_41/a_293_74#
+ prbs_generator_syn_19/sky130_fd_sc_hs__nand2_1_31/a_117_74# prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_5/a_138_385#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_63/a_1141_508# prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_19/a_222_392#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_13/a_1141_508# prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_3/a_52_123#
+ prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_13/a_52_123# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_43/a_1178_124#
+ prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_61/a_376_368# prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_35/a_132_392#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_67/a_206_368# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_1/a_1226_296#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_69/a_696_458# prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_31/a_230_79#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_35/a_735_102# prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_23/a_112_119#
+ prbs_generator_syn_19/sky130_fd_sc_hs__nand2_1_35/a_117_74# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_59/a_27_74#
+ prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_13/a_293_74# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_5/a_206_368#
+ prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_50/a_376_368# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_7/a_696_458#
+ prbs_generator_syn_19/sky130_fd_sc_hs__nor2b_1_7/a_278_368# prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_17/a_52_123#
+ prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_43/a_138_385# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_7/a_1141_508#
+ prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_61/a_52_123# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_67/a_437_503#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_61/a_1141_508# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_25/a_735_102#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_59/a_696_458# prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_13/a_112_119#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_33/a_1034_424# prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_51/a_112_119#
+ prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_35/a_230_79# prbs_generator_syn_19/m3_13600_4091#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_23/a_1226_296# prbs_generator_syn_19/sky130_fd_sc_hs__nand2_1_39/a_117_74#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_29/a_27_74# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_5/a_437_503#
+ prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_17/a_293_74# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_41/a_1178_124#
+ prbs_generator_syn_19/sky130_fd_sc_hs__or2_1_1/a_152_368# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_59/a_1178_124#
+ prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_61/a_293_74# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_47/a_206_368#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_39/a_651_503# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_49/a_696_458#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_15/a_735_102# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_32/a_1034_424#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_73/a_1226_296# prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_27/a_222_392#
+ prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_41/a_112_119# prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_31/a_52_123#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_49/a_1034_424# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_29/a_1141_508#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_21/a_1226_296# prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_39/a_230_79#
+ prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_23/a_138_385# prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_51/a_230_79#
+ prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_45/a_132_392# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_37/a_206_368#
+ prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_65/a_293_74# prbs_generator_syn_19/sky130_fd_sc_hs__nand2_1_53/a_117_74#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_47/a_437_503# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_29/a_651_503#
+ prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_31/a_293_74# prbs_generator_syn_19/sky130_fd_sc_hs__nand2_1_21/a_117_74#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_69/a_544_485# prbs_generator_syn_19/sky130_fd_sc_hs__clkbuf_16_1/a_114_74#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_45/a_735_102# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_13/a_27_74#
+ prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_31/a_112_119# prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_57/a_222_392#
+ prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_35/a_52_123# prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_21/a_376_368#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_7/a_544_485# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_57/a_1178_124#
+ prbs_generator_syn_19/m3_13600_6043# prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_13/a_138_385#
+ prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_51/a_138_385# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_5/a_1141_508#
+ prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_3/a_376_368# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_27/a_206_368#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_65/a_206_368# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_37/a_437_503#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_19/a_651_503# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_57/a_651_503#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_59/a_544_485# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_71/a_1226_296#
+ prbs_generator_syn_19/sky130_fd_sc_hs__nand2_1_25/a_117_74# prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_61/a_112_119#
+ prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_47/a_222_392# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_27/a_1141_508#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_53/a_27_74# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_4/a_206_368#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_39/a_1226_296# prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_11/a_376_368#
+ prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_39/a_52_123# prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_41/a_138_385#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_4/a_1141_508# prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_25/a_132_392#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_17/a_206_368# prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_41/A
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_55/a_206_368# prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_51/a_52_123#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_27/a_437_503# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_65/a_437_503#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_49/a_544_485# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_63/a_735_102#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_47/a_1034_424# prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_50/a_112_119#
+ prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_37/a_222_392# prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_59/a_230_79#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_25/a_1141_508# prbs_generator_syn_19/sky130_fd_sc_hs__nor2b_1_4/a_27_112#
+ prbs_generator_syn_19/sky130_fd_sc_hs__sdlclkp_2_1/a_685_81# prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_1/a_132_392#
+ prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_39/a_293_74# prbs_generator_syn_19/sky130_fd_sc_hs__nand2_1_29/a_117_74#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_4/a_437_503# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_55/a_1178_124#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_21/a_27_74# prbs_generator_syn_19/m3_13600_12875#
+ prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_50/a_293_74# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_1/a_735_102#
+ prbs_generator_syn_19/sky130_fd_sc_hs__xnor2_1_31/a_138_385# prbs_generator_syn_19/sky130_fd_sc_hs__a22o_1_15/a_132_392#
+ prbs_generator_syn_19/sky130_fd_sc_hs__nand2_1_1/a_117_74# prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_17/a_437_503#
+ prbs_generator_syn_19/sky130_fd_sc_hs__dfxtp_4_55/a_437_503# prbs_generator_syn
Xsky130_fd_sc_hs__buf_2_106 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__buf_2_111/X sky130_fd_sc_hs__buf_2_107/X
+ sky130_fd_sc_hs__buf_2_107/a_21_260# sky130_fd_sc_hs__buf_2
Xsky130_fd_sc_hs__buf_2_117 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__buf_2_117/A sky130_fd_sc_hs__buf_2_117/X
+ sky130_fd_sc_hs__buf_2_117/a_21_260# sky130_fd_sc_hs__buf_2
Xsky130_fd_sc_hs__buf_2_128 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__buf_2_129/A sky130_fd_sc_hs__buf_2_129/X
+ sky130_fd_sc_hs__buf_2_129/a_21_260# sky130_fd_sc_hs__buf_2
Xsky130_fd_sc_hs__buf_2_139 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__buf_2_139/A sky130_fd_sc_hs__buf_2_139/X
+ sky130_fd_sc_hs__buf_2_139/a_21_260# sky130_fd_sc_hs__buf_2
Xsky130_fd_sc_hs__einvp_2_18 DVSS: DVDD: DVDD: DVSS: dout_n sky130_fd_sc_hs__einvp_2_9/A
+ sky130_fd_sc_hs__dlrtp_1_1/Q sky130_fd_sc_hs__einvp_2_19/a_263_323# sky130_fd_sc_hs__einvp_2_19/a_36_74#
+ sky130_fd_sc_hs__einvp_2_19/a_27_368# sky130_fd_sc_hs__einvp_2
Xsky130_fd_sc_hs__einvp_2_29 DVSS: DVDD: DVDD: DVSS: dout_n sky130_fd_sc_hs__buf_8_1/A
+ sky130_fd_sc_hs__dlrtp_1_25/Q sky130_fd_sc_hs__einvp_2_29/a_263_323# sky130_fd_sc_hs__einvp_2_29/a_36_74#
+ sky130_fd_sc_hs__einvp_2_29/a_27_368# sky130_fd_sc_hs__einvp_2
Xsky130_fd_sc_hs__conb_1_17 DVSS: DVDD: DVDD: DVSS: prbs_generator_syn_3/eqn[22] prbs_generator_syn_3/eqn[20]
+ sky130_fd_sc_hs__conb_1_17/a_165_290# sky130_fd_sc_hs__conb_1_17/a_21_290# sky130_fd_sc_hs__conb_1
Xsky130_fd_sc_hs__conb_1_28 DVSS: DVDD: DVDD: DVSS: prbs_generator_syn_5/eqn[9] sky130_fd_sc_hs__conb_1_29/HI
+ sky130_fd_sc_hs__conb_1_29/a_165_290# sky130_fd_sc_hs__conb_1_29/a_21_290# sky130_fd_sc_hs__conb_1
Xsky130_fd_sc_hs__conb_1_39 DVSS: DVDD: DVDD: DVSS: prbs_generator_syn_9/eqn[28] sky130_fd_sc_hs__conb_1_39/HI
+ sky130_fd_sc_hs__conb_1_39/a_165_290# sky130_fd_sc_hs__conb_1_39/a_21_290# sky130_fd_sc_hs__conb_1
Xsky130_fd_sc_hs__inv_4_13 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__inv_4_13/Y sky130_fd_sc_hs__inv_4_13/A
+ sky130_fd_sc_hs__inv_4
Xsky130_fd_sc_hs__inv_4_24 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__inv_4_25/Y sky130_fd_sc_hs__inv_4_25/A
+ sky130_fd_sc_hs__inv_4
Xsky130_fd_sc_hs__inv_4_35 DVSS: DVDD: DVDD: DVSS: osc_core_1/pi1_r[0] osc_core_1/pi1_l[0]
+ sky130_fd_sc_hs__inv_4
Xsky130_fd_sc_hs__inv_4_46 DVSS: DVDD: DVDD: DVSS: osc_core_1/pi2_r[0] osc_core_1/pi2_l[0]
+ sky130_fd_sc_hs__inv_4
Xsky130_fd_sc_hs__inv_4_57 DVSS: DVDD: DVDD: DVSS: osc_core_1/pi3_r[0] osc_core_1/pi3_l[0]
+ sky130_fd_sc_hs__inv_4
Xsky130_fd_sc_hs__inv_4_68 DVSS: DVDD: DVDD: DVSS: osc_core_1/pi5_r[3] osc_core_1/pi5_l[3]
+ sky130_fd_sc_hs__inv_4
Xsky130_fd_sc_hs__inv_4_79 DVSS: DVDD: DVDD: DVSS: hr_16t4_mux_top_3/din[12] prbs_generator_syn_21/out
+ sky130_fd_sc_hs__inv_4
Xsky130_fd_sc_hs__conb_1_190 DVSS: DVDD: DVDD: DVSS: prbs_generator_syn_29/eqn[28]
+ sky130_fd_sc_hs__conb_1_191/HI sky130_fd_sc_hs__conb_1_191/a_165_290# sky130_fd_sc_hs__conb_1_191/a_21_290#
+ sky130_fd_sc_hs__conb_1
Xsky130_fd_sc_hs__dlrtp_1_19 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__dlrtp_1_19/Q
+ sky130_fd_sc_hs__dlrtp_1_9/GATE sky130_fd_sc_hs__conb_1_121/HI sky130_fd_sc_hs__dlrtp_1_19/D
+ sky130_fd_sc_hs__dlrtp_1_19/a_216_424# sky130_fd_sc_hs__dlrtp_1_19/a_759_508# sky130_fd_sc_hs__dlrtp_1_19/a_565_74#
+ sky130_fd_sc_hs__dlrtp_1_19/a_27_424# sky130_fd_sc_hs__dlrtp_1_19/a_1045_74# sky130_fd_sc_hs__dlrtp_1_19/a_643_74#
+ sky130_fd_sc_hs__dlrtp_1_19/a_817_48# sky130_fd_sc_hs__dlrtp_1_19/a_568_392# sky130_fd_sc_hs__dlrtp_1_19/a_363_74#
+ sky130_fd_sc_hs__dlrtp_1_19/a_769_74# sky130_fd_sc_hs__dlrtp_1
Xsky130_fd_sc_hs__clkbuf_16_40 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__einvp_2_9/A
+ sky130_fd_sc_hs__buf_8_1/A sky130_fd_sc_hs__clkbuf_16_41/a_114_74# sky130_fd_sc_hs__clkbuf_16
Xsky130_fd_sc_hs__clkbuf_16_51 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__clkbuf_16_53/A
+ sky130_fd_sc_hs__nand2_2_7/Y sky130_fd_sc_hs__clkbuf_16_51/a_114_74# sky130_fd_sc_hs__clkbuf_16
Xsky130_fd_sc_hs__clkbuf_16_62 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__nor4_2_1/C
+ sky130_fd_sc_hs__clkbuf_16_63/A sky130_fd_sc_hs__clkbuf_16_63/a_114_74# sky130_fd_sc_hs__clkbuf_16
Xsky130_fd_sc_hs__clkbuf_16_73 DVSS: DVDD: DVDD: DVSS: prbs_generator_syn_19/clk sky130_fd_sc_hs__clkbuf_16_75/X
+ sky130_fd_sc_hs__clkbuf_16_73/a_114_74# sky130_fd_sc_hs__clkbuf_16
Xsky130_fd_sc_hs__clkbuf_16_84 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__nand2_2_7/A
+ sky130_fd_sc_hs__clkbuf_16_99/X sky130_fd_sc_hs__clkbuf_16_85/a_114_74# sky130_fd_sc_hs__clkbuf_16
Xsky130_fd_sc_hs__clkbuf_16_95 DVSS: DVDD: DVDD: DVSS: osc_core_1/glob_en osc_en sky130_fd_sc_hs__clkbuf_16_95/a_114_74#
+ sky130_fd_sc_hs__clkbuf_16
Xsky130_fd_sc_hs__o21ai_4_0 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__o21ai_4_1/Y sky130_fd_sc_hs__o21ai_4_1/A1
+ sky130_fd_sc_hs__or2b_4_1/A sky130_fd_sc_hs__inv_4_19/Y sky130_fd_sc_hs__o21ai_4_1/a_116_368#
+ sky130_fd_sc_hs__o21ai_4_1/a_27_74# sky130_fd_sc_hs__o21ai_4
Xsky130_fd_sc_hs__nand2_2_14 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__nand2_2_15/Y
+ sky130_fd_sc_hs__nand2_2_15/B sky130_fd_sc_hs__inv_4_23/Y sky130_fd_sc_hs__nand2_2_15/a_27_74#
+ sky130_fd_sc_hs__nand2_2
Xsky130_fd_sc_hs__nand2_2_25 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__nand2_2_25/Y
+ sky130_fd_sc_hs__nor4_2_1/B sky130_fd_sc_hs__nor4_2_1/A sky130_fd_sc_hs__nand2_2_25/a_27_74#
+ sky130_fd_sc_hs__nand2_2
Xprbs_generator_syn_3 prbs_generator_syn_9/clk prbs_generator_syn_9/rst prbs_generator_syn_3/cke
+ sky130_fd_sc_hs__conb_1_49/LO sky130_fd_sc_hs__conb_1_49/LO sky130_fd_sc_hs__conb_1_49/LO
+ prbs_generator_syn_7/eqn[1] prbs_generator_syn_7/eqn[1] prbs_generator_syn_7/eqn[1]
+ prbs_generator_syn_7/eqn[1] prbs_generator_syn_7/eqn[1] sky130_fd_sc_hs__conb_1_49/HI
+ sky130_fd_sc_hs__conb_1_49/HI sky130_fd_sc_hs__conb_1_49/HI prbs_generator_syn_3/cke
+ prbs_generator_syn_3/cke prbs_generator_syn_3/cke prbs_generator_syn_7/eqn[9] sky130_fd_sc_hs__conb_1_51/HI
+ prbs_generator_syn_7/eqn[9] sky130_fd_sc_hs__conb_1_51/HI prbs_generator_syn_9/eqn[16]
+ prbs_generator_syn_9/eqn[16] prbs_generator_syn_9/eqn[22] prbs_generator_syn_9/eqn[22]
+ prbs_generator_syn_9/eqn[22] prbs_generator_syn_9/eqn[28] sky130_fd_sc_hs__conb_1_39/HI
+ sky130_fd_sc_hs__conb_1_39/HI prbs_generator_syn_9/eqn[28] prbs_generator_syn_9/eqn[30]
+ sky130_fd_sc_hs__conb_1_55/HI sky130_fd_sc_hs__conb_1_55/HI prbs_generator_syn_9/eqn[30]
+ prbs_generator_syn_9/eqn[30] prbs_generator_syn_3/eqn[31] prbs_generator_syn_3/eqn[30]
+ prbs_generator_syn_3/eqn[30] prbs_generator_syn_3/eqn[28] prbs_generator_syn_3/eqn[28]
+ prbs_generator_syn_3/eqn[28] prbs_generator_syn_3/eqn[28] prbs_generator_syn_3/eqn[28]
+ prbs_generator_syn_3/eqn[28] prbs_generator_syn_3/eqn[22] prbs_generator_syn_3/eqn[22]
+ prbs_generator_syn_3/eqn[20] prbs_generator_syn_3/eqn[22] prbs_generator_syn_3/eqn[22]
+ prbs_generator_syn_3/eqn[22] prbs_generator_syn_3/eqn[22] prbs_generator_syn_3/eqn[22]
+ prbs_generator_syn_3/eqn[9] prbs_generator_syn_3/eqn[9] prbs_generator_syn_3/eqn[9]
+ prbs_generator_syn_3/eqn[9] prbs_generator_syn_3/eqn[9] prbs_generator_syn_3/eqn[9]
+ prbs_generator_syn_3/eqn[8] prbs_generator_syn_3/eqn[8] prbs_generator_syn_3/eqn[8]
+ prbs_generator_syn_3/eqn[8] prbs_generator_syn_3/eqn[4] prbs_generator_syn_3/eqn[4]
+ prbs_generator_syn_3/eqn[4] prbs_generator_syn_3/eqn[1] prbs_generator_syn_3/eqn[4]
+ prbs_generator_syn_9/inj_err prbs_generator_syn_7/eqn[9] prbs_generator_syn_3/eqn[31]
+ prbs_generator_syn_3/out DVSS: DVDD: prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_1/a_293_74#
+ prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_15/X prbs_generator_syn_3/sky130_fd_sc_hs__nand2_1_35/B
+ prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_51/Y prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_9/A
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_9/CLK prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_47/a_27_74#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_37/a_1226_296# prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_3/B
+ prbs_generator_syn_3/sky130_fd_sc_hs__nor2b_1_7/a_27_112# prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_29/B
+ prbs_generator_syn_3/sky130_fd_sc_hs__sdlclkp_2_1/a_580_74# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_1/a_1141_508#
+ prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_5/Y prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_41/a_230_79#
+ prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_61/a_138_385# prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_43/a_132_392#
+ prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_3/a_222_392# prbs_generator_syn_3/sky130_fd_sc_hs__nor2b_1_9/a_27_112#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_61/a_27_74# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_35/a_206_368#
+ prbs_generator_syn_3/sky130_fd_sc_hs__nand2_2_3/Y prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_25/B
+ prbs_generator_syn_3/sky130_fd_sc_hs__nand2_1_11/a_117_74# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_67/a_651_503#
+ prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_45/X prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_39/a_696_458#
+ prbs_generator_syn_3/sky130_fd_sc_hs__sdlclkp_2_1/a_1198_74# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_45/a_1034_424#
+ prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_17/a_222_392# prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_55/a_222_392#
+ prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_53/Y prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_35/A
+ prbs_generator_syn_3/m3_13600_1651# prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_59/a_52_123#
+ prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_5/a_293_74# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_35/a_1226_296#
+ prbs_generator_syn_3/sky130_fd_sc_hs__nand2_1_51/B prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_5/a_651_503#
+ prbs_generator_syn_3/sky130_fd_sc_hs__nand2_1_21/B prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_8/a_27_74#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_15/a_27_74# prbs_generator_syn_3/sky130_fd_sc_hs__and2b_2_1/X
+ prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_13/X prbs_generator_syn_3/sky130_fd_sc_hs__nand2_2_3/a_27_74#
+ prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_50/a_138_385# prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_33/a_132_392#
+ prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_1/a_376_368# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_25/a_206_368#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_35/a_437_503# prbs_generator_syn_3/sky130_fd_sc_hs__sdlclkp_2_1/a_708_451#
+ prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_45/a_230_79# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_29/a_696_458#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_32/a_27_74# prbs_generator_syn_3/sky130_fd_sc_hs__nor2b_1_4/Y
+ prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_59/a_293_74# prbs_generator_syn_3/sky130_fd_sc_hs__nand2_1_47/a_117_74#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_73/a_735_102# prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_21/a_112_119#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_23/a_1141_508# prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_25/a_293_74#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_7/Q prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_3/a_112_119#
+ prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_35/B prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_51/X
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_53/a_1178_124# prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_23/a_132_392#
+ prbs_generator_syn_3/sky130_fd_sc_hs__nand2_1_3/B prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_15/a_206_368#
+ prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_63/a_132_392# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_55/a_27_74#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_25/a_437_503# prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_41/a_52_123#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_47/a_651_503# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_73/a_1141_508#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_19/a_696_458# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_57/a_696_458#
+ prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_7/X prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_43/a_1034_424#
+ prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_55/A prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_11/a_112_119#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_21/a_1141_508# prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_35/a_222_392#
+ prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_49/a_230_79# prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_67/Y
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_71/a_27_74# prbs_generator_syn_3/sky130_fd_sc_hs__nand2_1_33/B
+ prbs_generator_syn_3/sky130_fd_sc_hs__conb_1_1/LO prbs_generator_syn_3/sky130_fd_sc_hs__nand2_1_19/a_117_74#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_51/a_1178_124# prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_33/X
+ prbs_generator_syn_3/sky130_fd_sc_hs__nand2_1_29/B prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_41/Y
+ prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_53/a_132_392# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_45/a_206_368#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_15/a_437_503# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_37/a_651_503#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_39/a_544_485# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_53/a_735_102#
+ prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_45/a_52_123# prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_1/B
+ prbs_generator_syn_3/sky130_fd_sc_hs__nand2_2_3/B prbs_generator_syn_3/sky130_fd_sc_hs__clkbuf_16_1/A
+ prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_21/X prbs_generator_syn_3/sky130_fd_sc_hs__nand2_1_25/B
+ prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_39/a_376_368# prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_63/X
+ prbs_generator_syn_3/m3_13600_3481# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_69/a_1178_124#
+ prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_21/a_138_385# prbs_generator_syn_3/sky130_fd_sc_hs__nor2b_1_8/Y
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_19/a_1178_124# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_49/a_27_74#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_45/a_437_503# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_27/a_651_503#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_71/a_1141_508# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_65/a_651_503#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_29/a_544_485# prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_3/a_138_385#
+ prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_55/X prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_43/a_735_102#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_41/a_1034_424# prbs_generator_syn_3/sky130_fd_sc_hs__nand2_1_9/B
+ prbs_generator_syn_3/sky130_fd_sc_hs__nor2b_1_9/Y prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_59/a_1034_424#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_39/a_1141_508# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_33/a_1226_296#
+ prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_49/a_52_123# prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_47/Y
+ prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_43/Y prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_4/a_651_503#
+ prbs_generator_syn_3/sky130_fd_sc_hs__nand2_1_49/B prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_19/A
+ prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_11/a_138_385# prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_5/X
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_63/a_206_368# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_17/a_651_503#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_19/a_544_485# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_55/a_651_503#
+ prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_9/Y prbs_generator_syn_3/sky130_fd_sc_hs__nand2_1_17/B
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_57/a_544_485# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_67/a_696_458#
+ prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_35/X prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_19/a_27_74#
+ prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_45/a_222_392# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_32/a_1226_296#
+ prbs_generator_syn_3/sky130_fd_sc_hs__nand2_1_43/B prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_25/A
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_1/a_206_368# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_49/a_1226_296#
+ prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_1/a_112_119# prbs_generator_syn_3/sky130_fd_sc_hs__or2_1_1/X
+ prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_59/a_376_368# prbs_generator_syn_3/sky130_fd_sc_hs__nand2_1_19/B
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_5/a_696_458# prbs_generator_syn_3/sky130_fd_sc_hs__nor2b_1_1/Y
+ prbs_generator_syn_3/sky130_fd_sc_hs__nor2b_1_5/a_278_368# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_17/a_1178_124#
+ prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_39/X prbs_generator_syn_3/m3_13600_5433#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_63/a_437_503# prbs_generator_syn_3/sky130_fd_sc_hs__nand2_2_5/B
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_23/a_735_102# prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_53/A
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_61/a_735_102# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_57/a_1034_424#
+ prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_63/B prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_37/a_1141_508#
+ prbs_generator_syn_3/sky130_fd_sc_hs__nand2_1_47/B prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_29/X
+ prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_65/Y prbs_generator_syn_3/m3_13600_4701#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_1/a_437_503# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_67/a_1178_124#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_9/a_735_102# prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_13/a_132_392#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_15/a_1178_124# prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_15/A
+ prbs_generator_syn_3/sky130_fd_sc_hs__nand2_1_1/B prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_43/B
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_35/a_651_503# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_8/D
+ prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_29/A prbs_generator_syn_3/sky130_fd_sc_hs__nand2_1_7/B
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_13/a_735_102# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_47/a_696_458#
+ prbs_generator_syn_3/sky130_fd_sc_hs__nand2_1_31/B prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_51/a_735_102#
+ prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_59/X prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_35/a_1141_508#
+ prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_25/a_222_392# prbs_generator_syn_3/sky130_fd_sc_hs__sdlclkp_2_1/a_288_48#
+ prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_55/B prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_17/B
+ prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_43/A prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_7/A
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_65/a_1178_124# prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_59/Y
+ prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_41/X prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_21/a_230_79#
+ prbs_generator_syn_3/sky130_fd_sc_hs__nand2_1_57/a_117_74# prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_1/a_222_392#
+ prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_19/B prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_35/a_293_74#
+ prbs_generator_syn_3/sky130_fd_sc_hs__nand2_1_23/a_117_74# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_73/a_206_368#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_25/a_651_503# prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_1/a_138_385#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_37/a_696_458# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_67/a_544_485#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_43/a_27_74# prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_9/X
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_55/a_1034_424# prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_39/a_112_119#
+ prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_15/a_222_392# prbs_generator_syn_3/sky130_fd_sc_hs__conb_1_1/HI
+ prbs_generator_syn_3/sky130_fd_sc_hs__nand2_1_23/B prbs_generator_syn_3/sky130_fd_sc_hs__nand2_1_53/B
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_9/a_1178_124# prbs_generator_syn_3/sky130_fd_sc_hs__nor2b_1_4/A
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_47/a_1226_296# prbs_generator_syn_3/m3_13600_11045#
+ prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_17/X prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_29/a_376_368#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_5/a_544_485# prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_3/X
+ prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_31/a_132_392# prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_61/A
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_15/a_651_503# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_73/a_437_503#
+ prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_25/a_230_79# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_27/a_696_458#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_65/a_696_458# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_33/a_735_102#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_71/a_735_102# prbs_generator_syn_3/m3_13600_7263#
+ prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_43/a_222_392# prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_50/Y
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_8/a_1178_124# prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_53/B
+ prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_19/a_376_368# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_63/a_1178_124#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_4/a_696_458# prbs_generator_syn_3/sky130_fd_sc_hs__nor2b_1_4/a_278_368#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_13/a_1178_124# prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_61/a_132_392#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_53/a_206_368# prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_21/a_52_123#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_45/a_651_503# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_17/a_696_458#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_47/a_544_485# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_55/a_696_458#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_21/a_735_102# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_37/a_27_74#
+ prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_61/B prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_61/X
+ prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_59/a_112_119# prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_31/A
+ prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_33/a_222_392# prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_29/a_230_79#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_45/a_1226_296# prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_9/a_132_392#
+ prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_5/A prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_57/Y
+ prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_31/X prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_51/a_27_74#
+ prbs_generator_syn_3/sky130_fd_sc_hs__nor2b_1_8/a_27_112# prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_47/a_376_368#
+ prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_53/a_293_74# prbs_generator_syn_3/sky130_fd_sc_hs__nand2_1_43/a_117_74#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_8/a_735_102# prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_21/a_293_74#
+ prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_39/a_138_385# prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_63/Y
+ prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_51/a_132_392# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_43/a_206_368#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_53/a_437_503# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_37/a_544_485#
+ prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_57/X prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_53/a_1034_424#
+ prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_25/a_52_123# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_33/a_1141_508#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_63/Q prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_23/a_222_392#
+ prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_63/a_222_392# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_7/a_1178_124#
+ prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_53/X prbs_generator_syn_3/sky130_fd_sc_hs__nand2_2_5/Y
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_61/a_1178_124# prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_1/a_230_79#
+ prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_43/a_230_79# prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_11/a_230_79#
+ prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_41/a_132_392# prbs_generator_syn_3/sky130_fd_sc_hs__nand2_1_13/a_117_74#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_43/a_437_503# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_27/a_544_485#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_63/a_651_503# prbs_generator_syn_3/sky130_fd_sc_hs__nand2_1_7/a_117_74#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_35/a_696_458# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_65/a_544_485#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_51/a_1034_424# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_41/a_735_102#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_32/a_1141_508# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_49/a_1141_508#
+ prbs_generator_syn_3/sky130_fd_sc_hs__nand2_1_55/B prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_53/a_222_392#
+ prbs_generator_syn_3/sky130_fd_sc_hs__sdlclkp_2_1/a_114_112# prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_9/a_293_74#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_43/a_1226_296# prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_29/a_52_123#
+ prbs_generator_syn_3/sky130_fd_sc_hs__nand2_1_37/B prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_1/a_651_503#
+ prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_27/a_376_368# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_4/a_544_485#
+ prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_67/a_376_368# prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_27/X
+ prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_1/X prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_59/a_138_385#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_29/a_1178_124# prbs_generator_syn_3/m3_13600_2871#
+ prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_5/a_230_79# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_23/a_206_368#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_61/a_206_368# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_17/a_544_485#
+ prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_15/a_230_79# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_25/a_696_458#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_55/a_544_485# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_32/a_735_102#
+ prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_29/a_293_74# prbs_generator_syn_3/sky130_fd_sc_hs__nand2_1_17/a_117_74#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_69/a_1034_424# prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_29/a_112_119#
+ prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_37/X prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_31/B
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_19/a_1034_424# prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_33/A
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_9/a_206_368# prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_57/a_376_368#
+ prbs_generator_syn_3/sky130_fd_sc_hs__sdlclkp_2_1/a_706_317# prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_11/B
+ prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_1/a_52_123# prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_39/B
+ prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_21/a_132_392# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_13/a_206_368#
+ prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_43/a_52_123# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_51/a_206_368#
+ prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_47/X prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_23/a_437_503#
+ prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_11/a_52_123# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_61/a_437_503#
+ prbs_generator_syn_3/sky130_fd_sc_hs__nor2b_1_7/Y prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_51/A
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_15/a_696_458# prbs_generator_syn_3/sky130_fd_sc_hs__nor2b_1_5/Y
+ prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_9/a_230_79# prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_25/X
+ prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_19/a_112_119# prbs_generator_syn_3/sky130_fd_sc_hs__nand2_1_45/B
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_5/a_1178_124# prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_19/a_230_79#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_41/a_1226_296# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_59/a_1226_296#
+ prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_63/a_230_79# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_51/Q
+ prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_7/a_132_392# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_9/a_437_503#
+ prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_46/a_376_368# prbs_generator_syn_3/sky130_fd_sc_hs__nand2_1_33/a_117_74#
+ prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_11/a_293_74# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_27/a_1178_124#
+ prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_11/a_132_392# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_13/a_437_503#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_51/a_437_503# prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_5/a_52_123#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_35/a_544_485# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_73/a_651_503#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_45/a_696_458# prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_15/a_52_123#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_47/a_1141_508# prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_47/a_112_119#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_4/a_1178_124# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_17/a_1034_424#
+ prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_23/B prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_37/a_376_368#
+ prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_15/B prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_7/Y
+ prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_29/a_138_385# prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_33/a_230_79#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_25/a_1178_124# prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_47/a_293_74#
+ prbs_generator_syn_3/sky130_fd_sc_hs__nand2_1_37/a_117_74# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_33/a_206_368#
+ prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_15/a_293_74# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_71/a_206_368#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_25/a_544_485# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_67/a_1034_424#
+ prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_13/a_222_392# prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_9/a_52_123#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_15/a_1034_424# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_57/a_1226_296#
+ prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_19/a_52_123# prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_23/X
+ prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_63/a_52_123# prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_19/a_138_385#
+ prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_9/a_376_368# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_21/a_206_368#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_33/a_437_503# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_71/a_437_503#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_53/a_651_503# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_15/a_544_485#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_63/a_696_458# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_65/a_1034_424#
+ prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_19/a_293_74# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_45/a_1141_508#
+ prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_27/a_112_119# prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_67/a_112_119#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_1/a_1178_124# prbs_generator_syn_3/sky130_fd_sc_hs__conb_1_1/a_21_290#
+ prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_63/a_293_74# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_8/a_206_368#
+ prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_17/a_376_368# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_63/a_27_74#
+ prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_21/A prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_55/a_376_368#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_1/a_696_458# prbs_generator_syn_3/sky130_fd_sc_hs__nor2b_1_1/a_278_368#
+ prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_47/a_138_385# prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_33/a_52_123#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_9/a_1034_424# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_21/a_437_503#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_1/a_27_74# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_43/a_651_503#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_1/Q prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_45/a_544_485#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_69/a_735_102# prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_57/a_112_119#
+ prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_31/a_222_392# prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_13/A
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_55/a_1226_296# prbs_generator_syn_3/sky130_fd_sc_hs__nand2_2_5/a_27_74#
+ prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_53/a_230_79# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_8/a_437_503#
+ prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_67/a_293_74# prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_33/a_293_74#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_7/a_735_102# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_23/a_1178_124#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_41/a_206_368# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_8/a_1034_424#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_63/a_1034_424# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_59/a_735_102#
+ prbs_generator_syn_3/sky130_fd_sc_hs__nand2_1_5/B prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_43/a_1141_508#
+ prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_46/a_112_119# prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_61/a_222_392#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_13/a_1034_424# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_73/a_1178_124#
+ prbs_generator_syn_3/sky130_fd_sc_hs__nand2_1_27/B prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_13/B
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_57/a_27_74# prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_57/a_230_79#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_21/a_1178_124# prbs_generator_syn_3/sky130_fd_sc_hs__nor2b_1_1/a_27_112#
+ prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_27/a_138_385# prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_23/a_230_79#
+ prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_67/a_138_385# prbs_generator_syn_3/sky130_fd_sc_hs__nand2_1_41/B
+ prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_9/a_222_392# prbs_generator_syn_3/sky130_fd_sc_hs__nand2_1_27/a_117_74#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_32/a_206_368# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_23/a_651_503#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_41/a_437_503# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_73/a_27_74#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_61/a_651_503# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_63/a_544_485#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_49/a_735_102# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_73/a_696_458#
+ prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_37/a_112_119# prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_51/a_222_392#
+ prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_43/X prbs_generator_syn_3/sky130_fd_sc_hs__nand2_2_1/B
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_9/a_651_503# prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_53/a_52_123#
+ prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_49/X prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_25/a_376_368#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_1/a_544_485# prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_65/a_376_368#
+ prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_57/a_138_385# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_27/a_27_74#
+ prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_39/a_132_392# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_7/a_1034_424#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_13/a_651_503# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_32/a_437_503#
+ prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_27/a_230_79# prbs_generator_syn_3/m3_13600_12265#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_51/a_651_503# prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_59/B
+ prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_47/A prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_61/a_1034_424#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_41/a_1141_508# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_59/a_1141_508#
+ prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_41/a_222_392# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_53/a_1226_296#
+ prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_3/A prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_71/a_1178_124#
+ prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_9/a_112_119# prbs_generator_syn_3/sky130_fd_sc_hs__nand2_1_3/a_117_74#
+ prbs_generator_syn_3/m3_13600_8483# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_39/a_1178_124#
+ prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_57/a_52_123# prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_46/a_138_385#
+ prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_23/a_52_123# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_67/a_27_74#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_53/a_696_458# prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_17/a_112_119#
+ prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_11/A prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_55/a_112_119#
+ prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_1/A prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_51/a_1226_296#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_29/a_1034_424# prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_59/A
+ prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_23/A prbs_generator_syn_3/sky130_fd_sc_hs__nand2_1_39/B
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_5/a_27_74# prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_57/a_293_74#
+ prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_37/a_138_385# prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_59/a_132_392#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_33/a_651_503# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_71/a_651_503#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_43/a_696_458# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_73/a_544_485#
+ prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_27/a_52_123# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_57/a_1141_508#
+ prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_21/a_222_392# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_35/a_27_74#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_69/a_1226_296# prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_37/B
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_19/a_1226_296# prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_35/a_376_368#
+ prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_47/a_230_79# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_37/a_1178_124#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_5/a_1034_424# prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_49/a_132_392#
+ prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_7/a_222_392# prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_27/a_293_74#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_21/a_651_503# prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_9/a_138_385#
+ prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_11/a_222_392# prbs_generator_syn_3/m3_13600_14095#
+ prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_50/A prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_27/a_1034_424#
+ prbs_generator_syn_3/sky130_fd_sc_hs__nand2_1_13/B prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_8/a_651_503#
+ prbs_generator_syn_3/m3_13600_9703# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_35/a_1178_124#
+ prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_17/a_138_385# prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_55/a_138_385#
+ prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_7/a_230_79# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_4/a_1034_424#
+ prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_7/a_376_368# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_69/a_206_368#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_23/a_696_458# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_53/a_544_485#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_39/a_735_102# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_61/a_696_458#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_55/a_1141_508# prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_25/a_112_119#
+ prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_65/a_112_119# prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_43/a_293_74#
+ prbs_generator_syn_3/sky130_fd_sc_hs__nand2_1_57/B prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_25/a_1034_424#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_7/a_206_368# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_17/a_1226_296#
+ prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_15/a_376_368# prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_53/a_376_368#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_9/a_696_458# prbs_generator_syn_3/m3_13600_431#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_45/a_27_74# prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_47/a_52_123#
+ prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_29/a_132_392# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_59/a_206_368#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_69/a_437_503# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_41/a_651_503#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_43/a_544_485# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_13/a_696_458#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_29/a_735_102# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_51/a_696_458#
+ prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_61/Y prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_67/a_1226_296#
+ prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_5/a_132_392# prbs_generator_syn_3/sky130_fd_sc_hs__and2b_2_1/a_198_48#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_7/a_437_503# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_15/a_1226_296#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_69/a_27_74# prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_46/a_293_74#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_1/a_1034_424# prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_19/a_132_392#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_49/a_206_368# prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_7/a_52_123#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_59/a_437_503# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_32/a_651_503#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_7/a_27_74# prbs_generator_syn_3/sky130_fd_sc_hs__nand2_2_1/a_27_74#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_19/a_735_102# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_57/a_735_102#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_65/a_1226_296# prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_37/A
+ prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_33/a_376_368# prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_37/a_230_79#
+ prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_25/a_138_385# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_39/a_27_74#
+ prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_65/a_138_385# prbs_generator_syn_3/sky130_fd_sc_hs__nor2b_1_9/a_278_368#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_49/a_437_503# prbs_generator_syn_3/sky130_fd_sc_hs__and2b_2_1/a_505_74#
+ prbs_generator_syn_3/sky130_fd_sc_hs__nand2_1_51/a_117_74# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_23/a_544_485#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_33/a_696_458# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_61/a_544_485#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_9/a_1226_296# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_53/a_1141_508#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_71/a_696_458# prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_35/a_112_119#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_23/a_1034_424# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_9/a_544_485#
+ prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_63/a_376_368# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_33/a_1178_124#
+ prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_5/a_376_368# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_13/a_544_485#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_73/a_1034_424# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_21/a_696_458#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_51/a_544_485# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_8/a_1226_296#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_51/a_1141_508# prbs_generator_syn_3/sky130_fd_sc_hs__nand2_1_55/a_117_74#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_21/a_1034_424# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_63/a_1226_296#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_23/a_27_74# prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_7/a_112_119#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_13/a_1226_296# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_8/a_696_458#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_32/a_1178_124# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_49/a_1178_124#
+ prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_37/a_52_123# prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_27/a_132_392#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_71/Q prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_67/a_735_102#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_69/a_1141_508# prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_15/a_112_119#
+ prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_53/a_112_119# prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_39/a_222_392#
+ prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_55/a_230_79# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_19/a_1141_508#
+ prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_37/a_293_74# prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_43/a_376_368#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_5/a_735_102# prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_35/a_138_385#
+ prbs_generator_syn_3/sky130_fd_sc_hs__sdlclkp_2_1/a_114_424# prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_57/a_132_392#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_71/a_1034_424# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_7/a_1226_296#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_33/a_544_485# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_41/a_696_458#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_71/a_544_485# prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_21/B
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_61/a_1226_296# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_39/a_1034_424#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_17/a_27_74# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_9/a_27_74#
+ prbs_generator_syn_3/sky130_fd_sc_hs__nor2b_1_5/a_27_112# prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_47/a_132_392#
+ prbs_generator_syn_3/sky130_fd_sc_hs__nor2b_1_8/a_278_368# prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_9/B
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_39/a_206_368# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_33/a_27_74#
+ prbs_generator_syn_3/sky130_fd_sc_hs__nand2_1_41/a_117_74# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_69/a_651_503#
+ prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_51/a_293_74# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_21/a_544_485#
+ prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_7/a_138_385# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_32/a_696_458#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_47/a_735_102# prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_33/a_112_119#
+ prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_59/a_222_392# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_17/a_1141_508#
+ prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_55/a_52_123# prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_3/a_293_74#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_7/a_651_503# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_29/a_1226_296#
+ prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_23/a_376_368# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_8/a_544_485#
+ prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_47/B prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_47/a_1178_124#
+ prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_15/a_138_385# prbs_generator_syn_3/sky130_fd_sc_hs__sdlclkp_2_1/a_1195_374#
+ prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_53/a_138_385# prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_37/a_132_392#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_29/a_206_368# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_39/a_437_503#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_59/a_651_503# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_37/a_735_102#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_67/a_1141_508# prbs_generator_syn_3/sky130_fd_sc_hs__and2b_2_1/a_27_74#
+ prbs_generator_syn_3/sky130_fd_sc_hs__conb_1_1/a_165_290# prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_55/a_293_74#
+ prbs_generator_syn_3/sky130_fd_sc_hs__nand2_1_45/a_117_74# prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_63/a_112_119#
+ prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_49/a_222_392# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_37/a_1034_424#
+ prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_23/a_293_74# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_15/a_1141_508#
+ prbs_generator_syn_3/sky130_fd_sc_hs__nand2_1_5/a_117_74# prbs_generator_syn_3/m3_13600_13485#
+ prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_5/a_112_119# prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_13/a_376_368#
+ prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_51/a_376_368# prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_7/a_293_74#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_19/a_206_368# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_57/a_206_368#
+ prbs_generator_syn_3/sky130_fd_sc_hs__sdlclkp_2_1/a_318_74# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_29/a_437_503#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_49/a_651_503# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_25/a_27_74#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_5/a_1226_296# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_41/a_544_485#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_27/a_735_102# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_65/a_1141_508#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_65/a_735_102# prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_3/a_230_79#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_35/a_1034_424# prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_13/a_230_79#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_41/a_27_74# prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_3/a_132_392#
+ prbs_generator_syn_3/sky130_fd_sc_hs__nand2_1_49/a_117_74# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_27/a_1226_296#
+ prbs_generator_syn_3/sky130_fd_sc_hs__nand2_1_15/a_117_74# prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_41/a_376_368#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_45/a_1178_124# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_4/a_735_102#
+ prbs_generator_syn_3/sky130_fd_sc_hs__nand2_1_9/a_117_74# prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_33/a_138_385#
+ prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_17/a_132_392# prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_55/a_132_392#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_9/a_1141_508# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_19/a_437_503#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_57/a_437_503# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_4/a_1226_296#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_32/a_544_485# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_17/a_735_102#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_55/a_735_102# prbs_generator_syn_3/m3_13600_2261#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_65/a_27_74# prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_29/a_222_392#
+ prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_43/a_112_119# prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_19/X
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_25/a_1226_296# prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_31/a_376_368#
+ prbs_generator_syn_3/sky130_fd_sc_hs__or2_1_1/a_63_368# prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_17/a_230_79#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_4/a_27_74# prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_61/a_230_79#
+ prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_63/a_138_385# prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_5/a_222_392#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_8/a_1141_508# prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_41/a_293_74#
+ prbs_generator_syn_3/sky130_fd_sc_hs__nand2_1_31/a_117_74# prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_5/a_138_385#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_63/a_1141_508# prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_19/a_222_392#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_13/a_1141_508# prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_3/a_52_123#
+ prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_13/a_52_123# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_43/a_1178_124#
+ prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_61/a_376_368# prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_35/a_132_392#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_67/a_206_368# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_1/a_1226_296#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_69/a_696_458# prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_31/a_230_79#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_35/a_735_102# prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_23/a_112_119#
+ prbs_generator_syn_3/sky130_fd_sc_hs__nand2_1_35/a_117_74# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_59/a_27_74#
+ prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_13/a_293_74# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_5/a_206_368#
+ prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_50/a_376_368# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_7/a_696_458#
+ prbs_generator_syn_3/sky130_fd_sc_hs__nor2b_1_7/a_278_368# prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_17/a_52_123#
+ prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_43/a_138_385# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_7/a_1141_508#
+ prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_61/a_52_123# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_67/a_437_503#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_61/a_1141_508# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_25/a_735_102#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_59/a_696_458# prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_13/a_112_119#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_33/a_1034_424# prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_51/a_112_119#
+ prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_35/a_230_79# prbs_generator_syn_3/m3_13600_4091#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_23/a_1226_296# prbs_generator_syn_3/sky130_fd_sc_hs__nand2_1_39/a_117_74#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_29/a_27_74# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_5/a_437_503#
+ prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_17/a_293_74# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_41/a_1178_124#
+ prbs_generator_syn_3/sky130_fd_sc_hs__or2_1_1/a_152_368# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_59/a_1178_124#
+ prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_61/a_293_74# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_47/a_206_368#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_39/a_651_503# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_49/a_696_458#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_15/a_735_102# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_32/a_1034_424#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_73/a_1226_296# prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_27/a_222_392#
+ prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_41/a_112_119# prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_31/a_52_123#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_49/a_1034_424# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_29/a_1141_508#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_21/a_1226_296# prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_39/a_230_79#
+ prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_23/a_138_385# prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_51/a_230_79#
+ prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_45/a_132_392# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_37/a_206_368#
+ prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_65/a_293_74# prbs_generator_syn_3/sky130_fd_sc_hs__nand2_1_53/a_117_74#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_47/a_437_503# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_29/a_651_503#
+ prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_31/a_293_74# prbs_generator_syn_3/sky130_fd_sc_hs__nand2_1_21/a_117_74#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_69/a_544_485# prbs_generator_syn_3/sky130_fd_sc_hs__clkbuf_16_1/a_114_74#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_45/a_735_102# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_13/a_27_74#
+ prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_31/a_112_119# prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_57/a_222_392#
+ prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_35/a_52_123# prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_21/a_376_368#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_7/a_544_485# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_57/a_1178_124#
+ prbs_generator_syn_3/m3_13600_6043# prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_13/a_138_385#
+ prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_51/a_138_385# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_5/a_1141_508#
+ prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_3/a_376_368# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_27/a_206_368#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_65/a_206_368# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_37/a_437_503#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_19/a_651_503# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_57/a_651_503#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_59/a_544_485# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_71/a_1226_296#
+ prbs_generator_syn_3/sky130_fd_sc_hs__nand2_1_25/a_117_74# prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_61/a_112_119#
+ prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_47/a_222_392# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_27/a_1141_508#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_53/a_27_74# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_4/a_206_368#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_39/a_1226_296# prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_11/a_376_368#
+ prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_39/a_52_123# prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_41/a_138_385#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_4/a_1141_508# prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_25/a_132_392#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_17/a_206_368# prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_41/A
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_55/a_206_368# prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_51/a_52_123#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_27/a_437_503# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_65/a_437_503#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_49/a_544_485# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_63/a_735_102#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_47/a_1034_424# prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_50/a_112_119#
+ prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_37/a_222_392# prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_59/a_230_79#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_25/a_1141_508# prbs_generator_syn_3/sky130_fd_sc_hs__nor2b_1_4/a_27_112#
+ prbs_generator_syn_3/sky130_fd_sc_hs__sdlclkp_2_1/a_685_81# prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_1/a_132_392#
+ prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_39/a_293_74# prbs_generator_syn_3/sky130_fd_sc_hs__nand2_1_29/a_117_74#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_4/a_437_503# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_55/a_1178_124#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_21/a_27_74# prbs_generator_syn_3/m3_13600_12875#
+ prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_50/a_293_74# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_1/a_735_102#
+ prbs_generator_syn_3/sky130_fd_sc_hs__xnor2_1_31/a_138_385# prbs_generator_syn_3/sky130_fd_sc_hs__a22o_1_15/a_132_392#
+ prbs_generator_syn_3/sky130_fd_sc_hs__nand2_1_1/a_117_74# prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_17/a_437_503#
+ prbs_generator_syn_3/sky130_fd_sc_hs__dfxtp_4_55/a_437_503# prbs_generator_syn
Xsky130_fd_sc_hs__clkdlyinv5sd2_1_2 DVSS: DVDD: DVSS: DVDD: dout_p sky130_fd_sc_hs__nand2_2_1/A
+ sky130_fd_sc_hs__clkdlyinv5sd2_1_3/a_28_74# sky130_fd_sc_hs__clkdlyinv5sd2_1_3/a_682_74#
+ sky130_fd_sc_hs__clkdlyinv5sd2_1_3/a_549_74# sky130_fd_sc_hs__clkdlyinv5sd2_1_3/a_288_74#
+ sky130_fd_sc_hs__clkdlyinv5sd2_1
Xsky130_fd_sc_hs__nor4_2_0 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__nor4_2_1/C sky130_fd_sc_hs__nor4_2_1/A
+ sky130_fd_sc_hs__nor4_2_1/B sky130_fd_sc_hs__nor4_2_1/D sky130_fd_sc_hs__nor4_2_1/Y
+ sky130_fd_sc_hs__nor4_2_1/a_116_368# sky130_fd_sc_hs__nor4_2_1/a_490_368# sky130_fd_sc_hs__nor4_2_1/a_27_368#
+ sky130_fd_sc_hs__nor4_2
Xsky130_fd_sc_hs__clkbuf_4_90 DVSS: DVDD: DVDD: DVSS: div_ratio_half[4] sky130_fd_sc_hs__clkbuf_4_91/X
+ sky130_fd_sc_hs__clkbuf_4_91/a_83_270# sky130_fd_sc_hs__clkbuf_4
Xsky130_fd_sc_hs__einvn_8_0 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__inv_4_27/Y sky130_fd_sc_hs__clkinv_8_15/Y
+ sky130_fd_sc_hs__einvn_8_1/Z sky130_fd_sc_hs__einvn_8_1/a_126_74# sky130_fd_sc_hs__einvn_8_1/a_239_368#
+ sky130_fd_sc_hs__einvn_8_1/a_293_74# sky130_fd_sc_hs__einvn_8
Xsky130_fd_sc_hs__o21ai_2_15 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__inv_4_17/Y sky130_fd_sc_hs__o21ai_2_55/A1
+ sky130_fd_sc_hs__nand2_2_7/A sky130_fd_sc_hs__o21ai_2_15/Y sky130_fd_sc_hs__o21ai_2_15/a_116_368#
+ sky130_fd_sc_hs__o21ai_2_15/a_27_74# sky130_fd_sc_hs__o21ai_2
Xsky130_fd_sc_hs__o21ai_2_26 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__inv_4_21/Y sky130_fd_sc_hs__o21ai_2_31/A2
+ sky130_fd_sc_hs__buf_8_3/X sky130_fd_sc_hs__buf_2_85/A sky130_fd_sc_hs__o21ai_2_27/a_116_368#
+ sky130_fd_sc_hs__o21ai_2_27/a_27_74# sky130_fd_sc_hs__o21ai_2
Xsky130_fd_sc_hs__o21ai_2_37 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__inv_4_23/Y sky130_fd_sc_hs__or2b_4_1/A
+ sky130_fd_sc_hs__nand2_2_15/B sky130_fd_sc_hs__o21ai_2_37/Y sky130_fd_sc_hs__o21ai_2_37/a_116_368#
+ sky130_fd_sc_hs__o21ai_2_37/a_27_74# sky130_fd_sc_hs__o21ai_2
Xsky130_fd_sc_hs__o21ai_2_48 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__inv_4_25/Y sky130_fd_sc_hs__or2b_4_1/X
+ sky130_fd_sc_hs__o21ai_2_51/A1 sky130_fd_sc_hs__buf_2_135/A sky130_fd_sc_hs__o21ai_2_49/a_116_368#
+ sky130_fd_sc_hs__o21ai_2_49/a_27_74# sky130_fd_sc_hs__o21ai_2
Xsky130_fd_sc_hs__buf_2_107 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__buf_2_111/X sky130_fd_sc_hs__buf_2_107/X
+ sky130_fd_sc_hs__buf_2_107/a_21_260# sky130_fd_sc_hs__buf_2
Xsky130_fd_sc_hs__buf_2_118 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__buf_2_119/A sky130_fd_sc_hs__buf_2_119/X
+ sky130_fd_sc_hs__buf_2_119/a_21_260# sky130_fd_sc_hs__buf_2
Xsky130_fd_sc_hs__buf_2_129 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__buf_2_129/A sky130_fd_sc_hs__buf_2_129/X
+ sky130_fd_sc_hs__buf_2_129/a_21_260# sky130_fd_sc_hs__buf_2
Xsky130_fd_sc_hs__einvp_2_19 DVSS: DVDD: DVDD: DVSS: dout_n sky130_fd_sc_hs__einvp_2_9/A
+ sky130_fd_sc_hs__dlrtp_1_1/Q sky130_fd_sc_hs__einvp_2_19/a_263_323# sky130_fd_sc_hs__einvp_2_19/a_36_74#
+ sky130_fd_sc_hs__einvp_2_19/a_27_368# sky130_fd_sc_hs__einvp_2
Xsky130_fd_sc_hs__conb_1_18 DVSS: DVDD: DVDD: DVSS: prbs_generator_syn_9/eqn[22] prbs_generator_syn_9/eqn[20]
+ sky130_fd_sc_hs__conb_1_19/a_165_290# sky130_fd_sc_hs__conb_1_19/a_21_290# sky130_fd_sc_hs__conb_1
Xsky130_fd_sc_hs__conb_1_29 DVSS: DVDD: DVDD: DVSS: prbs_generator_syn_5/eqn[9] sky130_fd_sc_hs__conb_1_29/HI
+ sky130_fd_sc_hs__conb_1_29/a_165_290# sky130_fd_sc_hs__conb_1_29/a_21_290# sky130_fd_sc_hs__conb_1
Xsky130_fd_sc_hs__inv_4_14 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__inv_4_15/Y sky130_fd_sc_hs__inv_4_15/A
+ sky130_fd_sc_hs__inv_4
Xsky130_fd_sc_hs__inv_4_25 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__inv_4_25/Y sky130_fd_sc_hs__inv_4_25/A
+ sky130_fd_sc_hs__inv_4
Xsky130_fd_sc_hs__inv_4_36 DVSS: DVDD: DVDD: DVSS: osc_core_1/pi1_r[2] osc_core_1/pi1_l[2]
+ sky130_fd_sc_hs__inv_4
Xsky130_fd_sc_hs__inv_4_47 DVSS: DVDD: DVDD: DVSS: osc_core_1/pi2_r[0] osc_core_1/pi2_l[0]
+ sky130_fd_sc_hs__inv_4
Xsky130_fd_sc_hs__inv_4_58 DVSS: DVDD: DVDD: DVSS: osc_core_1/pi4_r[2] osc_core_1/pi4_l[2]
+ sky130_fd_sc_hs__inv_4
Xsky130_fd_sc_hs__inv_4_69 DVSS: DVDD: DVDD: DVSS: osc_core_1/pi5_r[3] osc_core_1/pi5_l[3]
+ sky130_fd_sc_hs__inv_4
Xsky130_fd_sc_hs__conb_1_180 DVSS: DVDD: DVDD: DVSS: prbs_generator_syn_23/eqn[28]
+ sky130_fd_sc_hs__conb_1_181/HI sky130_fd_sc_hs__conb_1_181/a_165_290# sky130_fd_sc_hs__conb_1_181/a_21_290#
+ sky130_fd_sc_hs__conb_1
Xsky130_fd_sc_hs__conb_1_191 DVSS: DVDD: DVDD: DVSS: prbs_generator_syn_29/eqn[28]
+ sky130_fd_sc_hs__conb_1_191/HI sky130_fd_sc_hs__conb_1_191/a_165_290# sky130_fd_sc_hs__conb_1_191/a_21_290#
+ sky130_fd_sc_hs__conb_1
Xsky130_fd_sc_hs__clkbuf_16_30 DVSS: DVDD: DVDD: DVSS: osc_core_1/pi2_l[3] sky130_fd_sc_hs__clkbuf_8_1/X
+ sky130_fd_sc_hs__clkbuf_16_31/a_114_74# sky130_fd_sc_hs__clkbuf_16
Xsky130_fd_sc_hs__clkbuf_16_41 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__einvp_2_9/A
+ sky130_fd_sc_hs__buf_8_1/A sky130_fd_sc_hs__clkbuf_16_41/a_114_74# sky130_fd_sc_hs__clkbuf_16
Xsky130_fd_sc_hs__clkbuf_16_52 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__clkbuf_16_53/X
+ sky130_fd_sc_hs__clkbuf_16_53/A sky130_fd_sc_hs__clkbuf_16_53/a_114_74# sky130_fd_sc_hs__clkbuf_16
Xsky130_fd_sc_hs__clkbuf_16_63 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__nor4_2_1/C
+ sky130_fd_sc_hs__clkbuf_16_63/A sky130_fd_sc_hs__clkbuf_16_63/a_114_74# sky130_fd_sc_hs__clkbuf_16
Xsky130_fd_sc_hs__clkbuf_16_74 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__clkbuf_16_75/X
+ sky130_fd_sc_hs__and2_4_1/X sky130_fd_sc_hs__clkbuf_16_75/a_114_74# sky130_fd_sc_hs__clkbuf_16
Xsky130_fd_sc_hs__clkbuf_16_85 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__nand2_2_7/A
+ sky130_fd_sc_hs__clkbuf_16_99/X sky130_fd_sc_hs__clkbuf_16_85/a_114_74# sky130_fd_sc_hs__clkbuf_16
Xsky130_fd_sc_hs__clkbuf_16_96 DVSS: DVDD: DVDD: DVSS: prbs_generator_syn_19/rst prbs_generator_syn_31/rst
+ sky130_fd_sc_hs__clkbuf_16_97/a_114_74# sky130_fd_sc_hs__clkbuf_16
Xsky130_fd_sc_hs__o21ai_4_1 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__o21ai_4_1/Y sky130_fd_sc_hs__o21ai_4_1/A1
+ sky130_fd_sc_hs__or2b_4_1/A sky130_fd_sc_hs__inv_4_19/Y sky130_fd_sc_hs__o21ai_4_1/a_116_368#
+ sky130_fd_sc_hs__o21ai_4_1/a_27_74# sky130_fd_sc_hs__o21ai_4
Xsky130_fd_sc_hs__nand2_2_15 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__nand2_2_15/Y
+ sky130_fd_sc_hs__nand2_2_15/B sky130_fd_sc_hs__inv_4_23/Y sky130_fd_sc_hs__nand2_2_15/a_27_74#
+ sky130_fd_sc_hs__nand2_2
Xsky130_fd_sc_hs__nand2_2_26 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__nand2_2_27/Y
+ sky130_fd_sc_hs__nand2_2_27/B sky130_fd_sc_hs__o21ai_4_1/A1 sky130_fd_sc_hs__nand2_2_27/a_27_74#
+ sky130_fd_sc_hs__nand2_2
Xprbs_generator_syn_4 prbs_generator_syn_9/clk prbs_generator_syn_9/rst prbs_generator_syn_5/cke
+ sky130_fd_sc_hs__conb_1_67/LO sky130_fd_sc_hs__conb_1_67/LO sky130_fd_sc_hs__conb_1_67/LO
+ sky130_fd_sc_hs__conb_1_67/LO sky130_fd_sc_hs__conb_1_67/LO sky130_fd_sc_hs__conb_1_67/LO
+ sky130_fd_sc_hs__conb_1_67/LO sky130_fd_sc_hs__conb_1_67/LO sky130_fd_sc_hs__conb_1_35/LO
+ sky130_fd_sc_hs__conb_1_35/LO sky130_fd_sc_hs__conb_1_35/LO sky130_fd_sc_hs__conb_1_35/HI
+ sky130_fd_sc_hs__conb_1_35/HI sky130_fd_sc_hs__conb_1_35/HI sky130_fd_sc_hs__conb_1_35/HI
+ sky130_fd_sc_hs__conb_1_35/HI sky130_fd_sc_hs__conb_1_35/HI sky130_fd_sc_hs__conb_1_35/HI
+ prbs_generator_syn_7/eqn[20] prbs_generator_syn_7/eqn[20] prbs_generator_syn_7/eqn[20]
+ prbs_generator_syn_7/eqn[20] prbs_generator_syn_7/eqn[20] sky130_fd_sc_hs__conb_1_69/HI
+ sky130_fd_sc_hs__conb_1_69/HI sky130_fd_sc_hs__conb_1_69/HI sky130_fd_sc_hs__conb_1_69/HI
+ prbs_generator_syn_7/cke prbs_generator_syn_7/cke prbs_generator_syn_7/cke prbs_generator_syn_7/cke
+ prbs_generator_syn_7/cke prbs_generator_syn_5/eqn[31] prbs_generator_syn_5/eqn[31]
+ prbs_generator_syn_5/eqn[31] prbs_generator_syn_5/eqn[31] prbs_generator_syn_5/eqn[31]
+ prbs_generator_syn_5/eqn[31] prbs_generator_syn_5/eqn[31] prbs_generator_syn_5/eqn[31]
+ prbs_generator_syn_5/eqn[23] prbs_generator_syn_5/eqn[23] prbs_generator_syn_5/eqn[23]
+ prbs_generator_syn_5/eqn[20] prbs_generator_syn_5/eqn[23] prbs_generator_syn_5/eqn[23]
+ prbs_generator_syn_5/eqn[23] prbs_generator_syn_5/eqn[23] prbs_generator_syn_5/eqn[23]
+ prbs_generator_syn_5/eqn[9] prbs_generator_syn_5/eqn[13] prbs_generator_syn_5/eqn[9]
+ prbs_generator_syn_5/eqn[9] prbs_generator_syn_5/eqn[9] prbs_generator_syn_5/eqn[9]
+ prbs_generator_syn_5/eqn[9] prbs_generator_syn_5/eqn[9] prbs_generator_syn_5/eqn[9]
+ prbs_generator_syn_5/eqn[5] prbs_generator_syn_5/eqn[5] prbs_generator_syn_5/eqn[5]
+ prbs_generator_syn_5/eqn[5] prbs_generator_syn_5/eqn[1] prbs_generator_syn_7/eqn[9]
+ prbs_generator_syn_9/inj_err sky130_fd_sc_hs__conb_1_35/LO sky130_fd_sc_hs__conb_1_35/LO
+ prbs_generator_syn_5/out DVSS: DVDD: prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_1/a_293_74#
+ prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_15/X prbs_generator_syn_5/sky130_fd_sc_hs__nand2_1_35/B
+ prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_51/Y prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_9/A
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_9/CLK prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_47/a_27_74#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_37/a_1226_296# prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_3/B
+ prbs_generator_syn_5/sky130_fd_sc_hs__nor2b_1_7/a_27_112# prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_29/B
+ prbs_generator_syn_5/sky130_fd_sc_hs__sdlclkp_2_1/a_580_74# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_1/a_1141_508#
+ prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_5/Y prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_41/a_230_79#
+ prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_61/a_138_385# prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_43/a_132_392#
+ prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_3/a_222_392# prbs_generator_syn_5/sky130_fd_sc_hs__nor2b_1_9/a_27_112#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_61/a_27_74# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_35/a_206_368#
+ prbs_generator_syn_5/sky130_fd_sc_hs__nand2_2_3/Y prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_25/B
+ prbs_generator_syn_5/sky130_fd_sc_hs__nand2_1_11/a_117_74# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_67/a_651_503#
+ prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_45/X prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_39/a_696_458#
+ prbs_generator_syn_5/sky130_fd_sc_hs__sdlclkp_2_1/a_1198_74# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_45/a_1034_424#
+ prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_17/a_222_392# prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_55/a_222_392#
+ prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_53/Y prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_35/A
+ prbs_generator_syn_5/m3_13600_1651# prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_59/a_52_123#
+ prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_5/a_293_74# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_35/a_1226_296#
+ prbs_generator_syn_5/sky130_fd_sc_hs__nand2_1_51/B prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_5/a_651_503#
+ prbs_generator_syn_5/sky130_fd_sc_hs__nand2_1_21/B prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_8/a_27_74#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_15/a_27_74# prbs_generator_syn_5/sky130_fd_sc_hs__and2b_2_1/X
+ prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_13/X prbs_generator_syn_5/sky130_fd_sc_hs__nand2_2_3/a_27_74#
+ prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_50/a_138_385# prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_33/a_132_392#
+ prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_1/a_376_368# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_25/a_206_368#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_35/a_437_503# prbs_generator_syn_5/sky130_fd_sc_hs__sdlclkp_2_1/a_708_451#
+ prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_45/a_230_79# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_29/a_696_458#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_32/a_27_74# prbs_generator_syn_5/sky130_fd_sc_hs__nor2b_1_4/Y
+ prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_59/a_293_74# prbs_generator_syn_5/sky130_fd_sc_hs__nand2_1_47/a_117_74#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_73/a_735_102# prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_21/a_112_119#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_23/a_1141_508# prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_25/a_293_74#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_7/Q prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_3/a_112_119#
+ prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_35/B prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_51/X
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_53/a_1178_124# prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_23/a_132_392#
+ prbs_generator_syn_5/sky130_fd_sc_hs__nand2_1_3/B prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_15/a_206_368#
+ prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_63/a_132_392# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_55/a_27_74#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_25/a_437_503# prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_41/a_52_123#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_47/a_651_503# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_73/a_1141_508#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_19/a_696_458# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_57/a_696_458#
+ prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_7/X prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_43/a_1034_424#
+ prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_55/A prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_11/a_112_119#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_21/a_1141_508# prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_35/a_222_392#
+ prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_49/a_230_79# prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_67/Y
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_71/a_27_74# prbs_generator_syn_5/sky130_fd_sc_hs__nand2_1_33/B
+ prbs_generator_syn_5/sky130_fd_sc_hs__conb_1_1/LO prbs_generator_syn_5/sky130_fd_sc_hs__nand2_1_19/a_117_74#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_51/a_1178_124# prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_33/X
+ prbs_generator_syn_5/sky130_fd_sc_hs__nand2_1_29/B prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_41/Y
+ prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_53/a_132_392# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_45/a_206_368#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_15/a_437_503# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_37/a_651_503#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_39/a_544_485# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_53/a_735_102#
+ prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_45/a_52_123# prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_1/B
+ prbs_generator_syn_5/sky130_fd_sc_hs__nand2_2_3/B prbs_generator_syn_5/sky130_fd_sc_hs__clkbuf_16_1/A
+ prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_21/X prbs_generator_syn_5/sky130_fd_sc_hs__nand2_1_25/B
+ prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_39/a_376_368# prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_63/X
+ prbs_generator_syn_5/m3_13600_3481# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_69/a_1178_124#
+ prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_21/a_138_385# prbs_generator_syn_5/sky130_fd_sc_hs__nor2b_1_8/Y
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_19/a_1178_124# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_49/a_27_74#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_45/a_437_503# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_27/a_651_503#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_71/a_1141_508# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_65/a_651_503#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_29/a_544_485# prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_3/a_138_385#
+ prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_55/X prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_43/a_735_102#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_41/a_1034_424# prbs_generator_syn_5/sky130_fd_sc_hs__nand2_1_9/B
+ prbs_generator_syn_5/sky130_fd_sc_hs__nor2b_1_9/Y prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_59/a_1034_424#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_39/a_1141_508# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_33/a_1226_296#
+ prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_49/a_52_123# prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_47/Y
+ prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_43/Y prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_4/a_651_503#
+ prbs_generator_syn_5/sky130_fd_sc_hs__nand2_1_49/B prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_19/A
+ prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_11/a_138_385# prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_5/X
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_63/a_206_368# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_17/a_651_503#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_19/a_544_485# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_55/a_651_503#
+ prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_9/Y prbs_generator_syn_5/sky130_fd_sc_hs__nand2_1_17/B
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_57/a_544_485# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_67/a_696_458#
+ prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_35/X prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_19/a_27_74#
+ prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_45/a_222_392# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_32/a_1226_296#
+ prbs_generator_syn_5/sky130_fd_sc_hs__nand2_1_43/B prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_25/A
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_1/a_206_368# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_49/a_1226_296#
+ prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_1/a_112_119# prbs_generator_syn_5/sky130_fd_sc_hs__or2_1_1/X
+ prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_59/a_376_368# prbs_generator_syn_5/sky130_fd_sc_hs__nand2_1_19/B
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_5/a_696_458# prbs_generator_syn_5/sky130_fd_sc_hs__nor2b_1_1/Y
+ prbs_generator_syn_5/sky130_fd_sc_hs__nor2b_1_5/a_278_368# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_17/a_1178_124#
+ prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_39/X prbs_generator_syn_5/m3_13600_5433#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_63/a_437_503# prbs_generator_syn_5/sky130_fd_sc_hs__nand2_2_5/B
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_23/a_735_102# prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_53/A
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_61/a_735_102# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_57/a_1034_424#
+ prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_63/B prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_37/a_1141_508#
+ prbs_generator_syn_5/sky130_fd_sc_hs__nand2_1_47/B prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_29/X
+ prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_65/Y prbs_generator_syn_5/m3_13600_4701#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_1/a_437_503# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_67/a_1178_124#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_9/a_735_102# prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_13/a_132_392#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_15/a_1178_124# prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_15/A
+ prbs_generator_syn_5/sky130_fd_sc_hs__nand2_1_1/B prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_43/B
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_35/a_651_503# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_8/D
+ prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_29/A prbs_generator_syn_5/sky130_fd_sc_hs__nand2_1_7/B
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_13/a_735_102# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_47/a_696_458#
+ prbs_generator_syn_5/sky130_fd_sc_hs__nand2_1_31/B prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_51/a_735_102#
+ prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_59/X prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_35/a_1141_508#
+ prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_25/a_222_392# prbs_generator_syn_5/sky130_fd_sc_hs__sdlclkp_2_1/a_288_48#
+ prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_55/B prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_17/B
+ prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_43/A prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_7/A
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_65/a_1178_124# prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_59/Y
+ prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_41/X prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_21/a_230_79#
+ prbs_generator_syn_5/sky130_fd_sc_hs__nand2_1_57/a_117_74# prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_1/a_222_392#
+ prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_19/B prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_35/a_293_74#
+ prbs_generator_syn_5/sky130_fd_sc_hs__nand2_1_23/a_117_74# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_73/a_206_368#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_25/a_651_503# prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_1/a_138_385#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_37/a_696_458# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_67/a_544_485#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_43/a_27_74# prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_9/X
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_55/a_1034_424# prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_39/a_112_119#
+ prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_15/a_222_392# prbs_generator_syn_5/sky130_fd_sc_hs__conb_1_1/HI
+ prbs_generator_syn_5/sky130_fd_sc_hs__nand2_1_23/B prbs_generator_syn_5/sky130_fd_sc_hs__nand2_1_53/B
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_9/a_1178_124# prbs_generator_syn_5/sky130_fd_sc_hs__nor2b_1_4/A
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_47/a_1226_296# prbs_generator_syn_5/m3_13600_11045#
+ prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_17/X prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_29/a_376_368#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_5/a_544_485# prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_3/X
+ prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_31/a_132_392# prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_61/A
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_15/a_651_503# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_73/a_437_503#
+ prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_25/a_230_79# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_27/a_696_458#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_65/a_696_458# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_33/a_735_102#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_71/a_735_102# prbs_generator_syn_5/m3_13600_7263#
+ prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_43/a_222_392# prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_50/Y
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_8/a_1178_124# prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_53/B
+ prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_19/a_376_368# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_63/a_1178_124#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_4/a_696_458# prbs_generator_syn_5/sky130_fd_sc_hs__nor2b_1_4/a_278_368#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_13/a_1178_124# prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_61/a_132_392#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_53/a_206_368# prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_21/a_52_123#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_45/a_651_503# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_17/a_696_458#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_47/a_544_485# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_55/a_696_458#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_21/a_735_102# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_37/a_27_74#
+ prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_61/B prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_61/X
+ prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_59/a_112_119# prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_31/A
+ prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_33/a_222_392# prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_29/a_230_79#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_45/a_1226_296# prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_9/a_132_392#
+ prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_5/A prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_57/Y
+ prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_31/X prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_51/a_27_74#
+ prbs_generator_syn_5/sky130_fd_sc_hs__nor2b_1_8/a_27_112# prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_47/a_376_368#
+ prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_53/a_293_74# prbs_generator_syn_5/sky130_fd_sc_hs__nand2_1_43/a_117_74#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_8/a_735_102# prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_21/a_293_74#
+ prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_39/a_138_385# prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_63/Y
+ prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_51/a_132_392# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_43/a_206_368#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_53/a_437_503# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_37/a_544_485#
+ prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_57/X prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_53/a_1034_424#
+ prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_25/a_52_123# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_33/a_1141_508#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_63/Q prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_23/a_222_392#
+ prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_63/a_222_392# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_7/a_1178_124#
+ prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_53/X prbs_generator_syn_5/sky130_fd_sc_hs__nand2_2_5/Y
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_61/a_1178_124# prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_1/a_230_79#
+ prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_43/a_230_79# prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_11/a_230_79#
+ prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_41/a_132_392# prbs_generator_syn_5/sky130_fd_sc_hs__nand2_1_13/a_117_74#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_43/a_437_503# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_27/a_544_485#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_63/a_651_503# prbs_generator_syn_5/sky130_fd_sc_hs__nand2_1_7/a_117_74#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_35/a_696_458# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_65/a_544_485#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_51/a_1034_424# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_41/a_735_102#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_32/a_1141_508# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_49/a_1141_508#
+ prbs_generator_syn_5/sky130_fd_sc_hs__nand2_1_55/B prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_53/a_222_392#
+ prbs_generator_syn_5/sky130_fd_sc_hs__sdlclkp_2_1/a_114_112# prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_9/a_293_74#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_43/a_1226_296# prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_29/a_52_123#
+ prbs_generator_syn_5/sky130_fd_sc_hs__nand2_1_37/B prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_1/a_651_503#
+ prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_27/a_376_368# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_4/a_544_485#
+ prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_67/a_376_368# prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_27/X
+ prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_1/X prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_59/a_138_385#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_29/a_1178_124# prbs_generator_syn_5/m3_13600_2871#
+ prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_5/a_230_79# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_23/a_206_368#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_61/a_206_368# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_17/a_544_485#
+ prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_15/a_230_79# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_25/a_696_458#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_55/a_544_485# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_32/a_735_102#
+ prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_29/a_293_74# prbs_generator_syn_5/sky130_fd_sc_hs__nand2_1_17/a_117_74#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_69/a_1034_424# prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_29/a_112_119#
+ prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_37/X prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_31/B
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_19/a_1034_424# prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_33/A
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_9/a_206_368# prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_57/a_376_368#
+ prbs_generator_syn_5/sky130_fd_sc_hs__sdlclkp_2_1/a_706_317# prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_11/B
+ prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_1/a_52_123# prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_39/B
+ prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_21/a_132_392# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_13/a_206_368#
+ prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_43/a_52_123# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_51/a_206_368#
+ prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_47/X prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_23/a_437_503#
+ prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_11/a_52_123# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_61/a_437_503#
+ prbs_generator_syn_5/sky130_fd_sc_hs__nor2b_1_7/Y prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_51/A
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_15/a_696_458# prbs_generator_syn_5/sky130_fd_sc_hs__nor2b_1_5/Y
+ prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_9/a_230_79# prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_25/X
+ prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_19/a_112_119# prbs_generator_syn_5/sky130_fd_sc_hs__nand2_1_45/B
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_5/a_1178_124# prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_19/a_230_79#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_41/a_1226_296# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_59/a_1226_296#
+ prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_63/a_230_79# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_51/Q
+ prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_7/a_132_392# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_9/a_437_503#
+ prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_46/a_376_368# prbs_generator_syn_5/sky130_fd_sc_hs__nand2_1_33/a_117_74#
+ prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_11/a_293_74# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_27/a_1178_124#
+ prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_11/a_132_392# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_13/a_437_503#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_51/a_437_503# prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_5/a_52_123#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_35/a_544_485# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_73/a_651_503#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_45/a_696_458# prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_15/a_52_123#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_47/a_1141_508# prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_47/a_112_119#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_4/a_1178_124# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_17/a_1034_424#
+ prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_23/B prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_37/a_376_368#
+ prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_15/B prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_7/Y
+ prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_29/a_138_385# prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_33/a_230_79#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_25/a_1178_124# prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_47/a_293_74#
+ prbs_generator_syn_5/sky130_fd_sc_hs__nand2_1_37/a_117_74# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_33/a_206_368#
+ prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_15/a_293_74# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_71/a_206_368#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_25/a_544_485# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_67/a_1034_424#
+ prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_13/a_222_392# prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_9/a_52_123#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_15/a_1034_424# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_57/a_1226_296#
+ prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_19/a_52_123# prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_23/X
+ prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_63/a_52_123# prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_19/a_138_385#
+ prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_9/a_376_368# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_21/a_206_368#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_33/a_437_503# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_71/a_437_503#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_53/a_651_503# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_15/a_544_485#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_63/a_696_458# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_65/a_1034_424#
+ prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_19/a_293_74# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_45/a_1141_508#
+ prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_27/a_112_119# prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_67/a_112_119#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_1/a_1178_124# prbs_generator_syn_5/sky130_fd_sc_hs__conb_1_1/a_21_290#
+ prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_63/a_293_74# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_8/a_206_368#
+ prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_17/a_376_368# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_63/a_27_74#
+ prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_21/A prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_55/a_376_368#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_1/a_696_458# prbs_generator_syn_5/sky130_fd_sc_hs__nor2b_1_1/a_278_368#
+ prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_47/a_138_385# prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_33/a_52_123#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_9/a_1034_424# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_21/a_437_503#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_1/a_27_74# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_43/a_651_503#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_1/Q prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_45/a_544_485#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_69/a_735_102# prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_57/a_112_119#
+ prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_31/a_222_392# prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_13/A
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_55/a_1226_296# prbs_generator_syn_5/sky130_fd_sc_hs__nand2_2_5/a_27_74#
+ prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_53/a_230_79# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_8/a_437_503#
+ prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_67/a_293_74# prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_33/a_293_74#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_7/a_735_102# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_23/a_1178_124#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_41/a_206_368# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_8/a_1034_424#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_63/a_1034_424# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_59/a_735_102#
+ prbs_generator_syn_5/sky130_fd_sc_hs__nand2_1_5/B prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_43/a_1141_508#
+ prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_46/a_112_119# prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_61/a_222_392#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_13/a_1034_424# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_73/a_1178_124#
+ prbs_generator_syn_5/sky130_fd_sc_hs__nand2_1_27/B prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_13/B
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_57/a_27_74# prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_57/a_230_79#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_21/a_1178_124# prbs_generator_syn_5/sky130_fd_sc_hs__nor2b_1_1/a_27_112#
+ prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_27/a_138_385# prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_23/a_230_79#
+ prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_67/a_138_385# prbs_generator_syn_5/sky130_fd_sc_hs__nand2_1_41/B
+ prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_9/a_222_392# prbs_generator_syn_5/sky130_fd_sc_hs__nand2_1_27/a_117_74#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_32/a_206_368# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_23/a_651_503#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_41/a_437_503# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_73/a_27_74#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_61/a_651_503# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_63/a_544_485#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_49/a_735_102# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_73/a_696_458#
+ prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_37/a_112_119# prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_51/a_222_392#
+ prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_43/X prbs_generator_syn_5/sky130_fd_sc_hs__nand2_2_1/B
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_9/a_651_503# prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_53/a_52_123#
+ prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_49/X prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_25/a_376_368#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_1/a_544_485# prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_65/a_376_368#
+ prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_57/a_138_385# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_27/a_27_74#
+ prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_39/a_132_392# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_7/a_1034_424#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_13/a_651_503# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_32/a_437_503#
+ prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_27/a_230_79# prbs_generator_syn_5/m3_13600_12265#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_51/a_651_503# prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_59/B
+ prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_47/A prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_61/a_1034_424#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_41/a_1141_508# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_59/a_1141_508#
+ prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_41/a_222_392# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_53/a_1226_296#
+ prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_3/A prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_71/a_1178_124#
+ prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_9/a_112_119# prbs_generator_syn_5/sky130_fd_sc_hs__nand2_1_3/a_117_74#
+ prbs_generator_syn_5/m3_13600_8483# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_39/a_1178_124#
+ prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_57/a_52_123# prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_46/a_138_385#
+ prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_23/a_52_123# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_67/a_27_74#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_53/a_696_458# prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_17/a_112_119#
+ prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_11/A prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_55/a_112_119#
+ prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_1/A prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_51/a_1226_296#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_29/a_1034_424# prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_59/A
+ prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_23/A prbs_generator_syn_5/sky130_fd_sc_hs__nand2_1_39/B
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_5/a_27_74# prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_57/a_293_74#
+ prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_37/a_138_385# prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_59/a_132_392#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_33/a_651_503# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_71/a_651_503#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_43/a_696_458# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_73/a_544_485#
+ prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_27/a_52_123# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_57/a_1141_508#
+ prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_21/a_222_392# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_35/a_27_74#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_69/a_1226_296# prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_37/B
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_19/a_1226_296# prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_35/a_376_368#
+ prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_47/a_230_79# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_37/a_1178_124#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_5/a_1034_424# prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_49/a_132_392#
+ prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_7/a_222_392# prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_27/a_293_74#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_21/a_651_503# prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_9/a_138_385#
+ prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_11/a_222_392# prbs_generator_syn_5/m3_13600_14095#
+ prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_50/A prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_27/a_1034_424#
+ prbs_generator_syn_5/sky130_fd_sc_hs__nand2_1_13/B prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_8/a_651_503#
+ prbs_generator_syn_5/m3_13600_9703# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_35/a_1178_124#
+ prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_17/a_138_385# prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_55/a_138_385#
+ prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_7/a_230_79# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_4/a_1034_424#
+ prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_7/a_376_368# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_69/a_206_368#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_23/a_696_458# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_53/a_544_485#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_39/a_735_102# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_61/a_696_458#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_55/a_1141_508# prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_25/a_112_119#
+ prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_65/a_112_119# prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_43/a_293_74#
+ prbs_generator_syn_5/sky130_fd_sc_hs__nand2_1_57/B prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_25/a_1034_424#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_7/a_206_368# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_17/a_1226_296#
+ prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_15/a_376_368# prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_53/a_376_368#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_9/a_696_458# prbs_generator_syn_5/m3_13600_431#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_45/a_27_74# prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_47/a_52_123#
+ prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_29/a_132_392# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_59/a_206_368#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_69/a_437_503# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_41/a_651_503#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_43/a_544_485# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_13/a_696_458#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_29/a_735_102# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_51/a_696_458#
+ prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_61/Y prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_67/a_1226_296#
+ prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_5/a_132_392# prbs_generator_syn_5/sky130_fd_sc_hs__and2b_2_1/a_198_48#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_7/a_437_503# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_15/a_1226_296#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_69/a_27_74# prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_46/a_293_74#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_1/a_1034_424# prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_19/a_132_392#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_49/a_206_368# prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_7/a_52_123#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_59/a_437_503# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_32/a_651_503#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_7/a_27_74# prbs_generator_syn_5/sky130_fd_sc_hs__nand2_2_1/a_27_74#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_19/a_735_102# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_57/a_735_102#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_65/a_1226_296# prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_37/A
+ prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_33/a_376_368# prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_37/a_230_79#
+ prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_25/a_138_385# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_39/a_27_74#
+ prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_65/a_138_385# prbs_generator_syn_5/sky130_fd_sc_hs__nor2b_1_9/a_278_368#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_49/a_437_503# prbs_generator_syn_5/sky130_fd_sc_hs__and2b_2_1/a_505_74#
+ prbs_generator_syn_5/sky130_fd_sc_hs__nand2_1_51/a_117_74# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_23/a_544_485#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_33/a_696_458# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_61/a_544_485#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_9/a_1226_296# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_53/a_1141_508#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_71/a_696_458# prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_35/a_112_119#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_23/a_1034_424# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_9/a_544_485#
+ prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_63/a_376_368# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_33/a_1178_124#
+ prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_5/a_376_368# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_13/a_544_485#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_73/a_1034_424# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_21/a_696_458#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_51/a_544_485# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_8/a_1226_296#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_51/a_1141_508# prbs_generator_syn_5/sky130_fd_sc_hs__nand2_1_55/a_117_74#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_21/a_1034_424# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_63/a_1226_296#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_23/a_27_74# prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_7/a_112_119#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_13/a_1226_296# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_8/a_696_458#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_32/a_1178_124# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_49/a_1178_124#
+ prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_37/a_52_123# prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_27/a_132_392#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_71/Q prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_67/a_735_102#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_69/a_1141_508# prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_15/a_112_119#
+ prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_53/a_112_119# prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_39/a_222_392#
+ prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_55/a_230_79# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_19/a_1141_508#
+ prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_37/a_293_74# prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_43/a_376_368#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_5/a_735_102# prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_35/a_138_385#
+ prbs_generator_syn_5/sky130_fd_sc_hs__sdlclkp_2_1/a_114_424# prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_57/a_132_392#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_71/a_1034_424# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_7/a_1226_296#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_33/a_544_485# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_41/a_696_458#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_71/a_544_485# prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_21/B
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_61/a_1226_296# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_39/a_1034_424#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_17/a_27_74# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_9/a_27_74#
+ prbs_generator_syn_5/sky130_fd_sc_hs__nor2b_1_5/a_27_112# prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_47/a_132_392#
+ prbs_generator_syn_5/sky130_fd_sc_hs__nor2b_1_8/a_278_368# prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_9/B
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_39/a_206_368# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_33/a_27_74#
+ prbs_generator_syn_5/sky130_fd_sc_hs__nand2_1_41/a_117_74# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_69/a_651_503#
+ prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_51/a_293_74# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_21/a_544_485#
+ prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_7/a_138_385# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_32/a_696_458#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_47/a_735_102# prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_33/a_112_119#
+ prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_59/a_222_392# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_17/a_1141_508#
+ prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_55/a_52_123# prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_3/a_293_74#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_7/a_651_503# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_29/a_1226_296#
+ prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_23/a_376_368# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_8/a_544_485#
+ prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_47/B prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_47/a_1178_124#
+ prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_15/a_138_385# prbs_generator_syn_5/sky130_fd_sc_hs__sdlclkp_2_1/a_1195_374#
+ prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_53/a_138_385# prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_37/a_132_392#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_29/a_206_368# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_39/a_437_503#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_59/a_651_503# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_37/a_735_102#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_67/a_1141_508# prbs_generator_syn_5/sky130_fd_sc_hs__and2b_2_1/a_27_74#
+ prbs_generator_syn_5/sky130_fd_sc_hs__conb_1_1/a_165_290# prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_55/a_293_74#
+ prbs_generator_syn_5/sky130_fd_sc_hs__nand2_1_45/a_117_74# prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_63/a_112_119#
+ prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_49/a_222_392# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_37/a_1034_424#
+ prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_23/a_293_74# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_15/a_1141_508#
+ prbs_generator_syn_5/sky130_fd_sc_hs__nand2_1_5/a_117_74# prbs_generator_syn_5/m3_13600_13485#
+ prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_5/a_112_119# prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_13/a_376_368#
+ prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_51/a_376_368# prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_7/a_293_74#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_19/a_206_368# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_57/a_206_368#
+ prbs_generator_syn_5/sky130_fd_sc_hs__sdlclkp_2_1/a_318_74# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_29/a_437_503#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_49/a_651_503# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_25/a_27_74#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_5/a_1226_296# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_41/a_544_485#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_27/a_735_102# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_65/a_1141_508#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_65/a_735_102# prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_3/a_230_79#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_35/a_1034_424# prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_13/a_230_79#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_41/a_27_74# prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_3/a_132_392#
+ prbs_generator_syn_5/sky130_fd_sc_hs__nand2_1_49/a_117_74# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_27/a_1226_296#
+ prbs_generator_syn_5/sky130_fd_sc_hs__nand2_1_15/a_117_74# prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_41/a_376_368#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_45/a_1178_124# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_4/a_735_102#
+ prbs_generator_syn_5/sky130_fd_sc_hs__nand2_1_9/a_117_74# prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_33/a_138_385#
+ prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_17/a_132_392# prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_55/a_132_392#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_9/a_1141_508# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_19/a_437_503#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_57/a_437_503# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_4/a_1226_296#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_32/a_544_485# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_17/a_735_102#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_55/a_735_102# prbs_generator_syn_5/m3_13600_2261#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_65/a_27_74# prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_29/a_222_392#
+ prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_43/a_112_119# prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_19/X
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_25/a_1226_296# prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_31/a_376_368#
+ prbs_generator_syn_5/sky130_fd_sc_hs__or2_1_1/a_63_368# prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_17/a_230_79#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_4/a_27_74# prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_61/a_230_79#
+ prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_63/a_138_385# prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_5/a_222_392#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_8/a_1141_508# prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_41/a_293_74#
+ prbs_generator_syn_5/sky130_fd_sc_hs__nand2_1_31/a_117_74# prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_5/a_138_385#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_63/a_1141_508# prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_19/a_222_392#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_13/a_1141_508# prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_3/a_52_123#
+ prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_13/a_52_123# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_43/a_1178_124#
+ prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_61/a_376_368# prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_35/a_132_392#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_67/a_206_368# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_1/a_1226_296#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_69/a_696_458# prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_31/a_230_79#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_35/a_735_102# prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_23/a_112_119#
+ prbs_generator_syn_5/sky130_fd_sc_hs__nand2_1_35/a_117_74# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_59/a_27_74#
+ prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_13/a_293_74# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_5/a_206_368#
+ prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_50/a_376_368# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_7/a_696_458#
+ prbs_generator_syn_5/sky130_fd_sc_hs__nor2b_1_7/a_278_368# prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_17/a_52_123#
+ prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_43/a_138_385# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_7/a_1141_508#
+ prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_61/a_52_123# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_67/a_437_503#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_61/a_1141_508# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_25/a_735_102#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_59/a_696_458# prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_13/a_112_119#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_33/a_1034_424# prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_51/a_112_119#
+ prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_35/a_230_79# prbs_generator_syn_5/m3_13600_4091#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_23/a_1226_296# prbs_generator_syn_5/sky130_fd_sc_hs__nand2_1_39/a_117_74#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_29/a_27_74# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_5/a_437_503#
+ prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_17/a_293_74# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_41/a_1178_124#
+ prbs_generator_syn_5/sky130_fd_sc_hs__or2_1_1/a_152_368# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_59/a_1178_124#
+ prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_61/a_293_74# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_47/a_206_368#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_39/a_651_503# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_49/a_696_458#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_15/a_735_102# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_32/a_1034_424#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_73/a_1226_296# prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_27/a_222_392#
+ prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_41/a_112_119# prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_31/a_52_123#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_49/a_1034_424# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_29/a_1141_508#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_21/a_1226_296# prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_39/a_230_79#
+ prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_23/a_138_385# prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_51/a_230_79#
+ prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_45/a_132_392# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_37/a_206_368#
+ prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_65/a_293_74# prbs_generator_syn_5/sky130_fd_sc_hs__nand2_1_53/a_117_74#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_47/a_437_503# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_29/a_651_503#
+ prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_31/a_293_74# prbs_generator_syn_5/sky130_fd_sc_hs__nand2_1_21/a_117_74#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_69/a_544_485# prbs_generator_syn_5/sky130_fd_sc_hs__clkbuf_16_1/a_114_74#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_45/a_735_102# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_13/a_27_74#
+ prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_31/a_112_119# prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_57/a_222_392#
+ prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_35/a_52_123# prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_21/a_376_368#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_7/a_544_485# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_57/a_1178_124#
+ prbs_generator_syn_5/m3_13600_6043# prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_13/a_138_385#
+ prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_51/a_138_385# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_5/a_1141_508#
+ prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_3/a_376_368# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_27/a_206_368#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_65/a_206_368# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_37/a_437_503#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_19/a_651_503# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_57/a_651_503#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_59/a_544_485# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_71/a_1226_296#
+ prbs_generator_syn_5/sky130_fd_sc_hs__nand2_1_25/a_117_74# prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_61/a_112_119#
+ prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_47/a_222_392# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_27/a_1141_508#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_53/a_27_74# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_4/a_206_368#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_39/a_1226_296# prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_11/a_376_368#
+ prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_39/a_52_123# prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_41/a_138_385#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_4/a_1141_508# prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_25/a_132_392#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_17/a_206_368# prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_41/A
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_55/a_206_368# prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_51/a_52_123#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_27/a_437_503# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_65/a_437_503#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_49/a_544_485# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_63/a_735_102#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_47/a_1034_424# prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_50/a_112_119#
+ prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_37/a_222_392# prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_59/a_230_79#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_25/a_1141_508# prbs_generator_syn_5/sky130_fd_sc_hs__nor2b_1_4/a_27_112#
+ prbs_generator_syn_5/sky130_fd_sc_hs__sdlclkp_2_1/a_685_81# prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_1/a_132_392#
+ prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_39/a_293_74# prbs_generator_syn_5/sky130_fd_sc_hs__nand2_1_29/a_117_74#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_4/a_437_503# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_55/a_1178_124#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_21/a_27_74# prbs_generator_syn_5/m3_13600_12875#
+ prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_50/a_293_74# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_1/a_735_102#
+ prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_31/a_138_385# prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_15/a_132_392#
+ prbs_generator_syn_5/sky130_fd_sc_hs__nand2_1_1/a_117_74# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_17/a_437_503#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_55/a_437_503# prbs_generator_syn
Xsky130_fd_sc_hs__clkdlyinv5sd2_1_3 DVSS: DVDD: DVSS: DVDD: dout_p sky130_fd_sc_hs__nand2_2_1/A
+ sky130_fd_sc_hs__clkdlyinv5sd2_1_3/a_28_74# sky130_fd_sc_hs__clkdlyinv5sd2_1_3/a_682_74#
+ sky130_fd_sc_hs__clkdlyinv5sd2_1_3/a_549_74# sky130_fd_sc_hs__clkdlyinv5sd2_1_3/a_288_74#
+ sky130_fd_sc_hs__clkdlyinv5sd2_1
Xsky130_fd_sc_hs__nor4_2_1 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__nor4_2_1/C sky130_fd_sc_hs__nor4_2_1/A
+ sky130_fd_sc_hs__nor4_2_1/B sky130_fd_sc_hs__nor4_2_1/D sky130_fd_sc_hs__nor4_2_1/Y
+ sky130_fd_sc_hs__nor4_2_1/a_116_368# sky130_fd_sc_hs__nor4_2_1/a_490_368# sky130_fd_sc_hs__nor4_2_1/a_27_368#
+ sky130_fd_sc_hs__nor4_2
Xsky130_fd_sc_hs__clkbuf_4_80 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__nand2_8_1/Y
+ sky130_fd_sc_hs__clkbuf_4_81/X sky130_fd_sc_hs__clkbuf_4_81/a_83_270# sky130_fd_sc_hs__clkbuf_4
Xsky130_fd_sc_hs__clkbuf_4_91 DVSS: DVDD: DVDD: DVSS: div_ratio_half[4] sky130_fd_sc_hs__clkbuf_4_91/X
+ sky130_fd_sc_hs__clkbuf_4_91/a_83_270# sky130_fd_sc_hs__clkbuf_4
Xsky130_fd_sc_hs__einvn_8_1 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__inv_4_27/Y sky130_fd_sc_hs__clkinv_8_15/Y
+ sky130_fd_sc_hs__einvn_8_1/Z sky130_fd_sc_hs__einvn_8_1/a_126_74# sky130_fd_sc_hs__einvn_8_1/a_239_368#
+ sky130_fd_sc_hs__einvn_8_1/a_293_74# sky130_fd_sc_hs__einvn_8
Xsky130_fd_sc_hs__o21ai_2_16 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__inv_4_17/Y sky130_fd_sc_hs__or2b_4_5/X
+ sky130_fd_sc_hs__nand2_2_7/A sky130_fd_sc_hs__o21ai_2_17/Y sky130_fd_sc_hs__o21ai_2_17/a_116_368#
+ sky130_fd_sc_hs__o21ai_2_17/a_27_74# sky130_fd_sc_hs__o21ai_2
Xsky130_fd_sc_hs__o21ai_2_27 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__inv_4_21/Y sky130_fd_sc_hs__o21ai_2_31/A2
+ sky130_fd_sc_hs__buf_8_3/X sky130_fd_sc_hs__buf_2_85/A sky130_fd_sc_hs__o21ai_2_27/a_116_368#
+ sky130_fd_sc_hs__o21ai_2_27/a_27_74# sky130_fd_sc_hs__o21ai_2
Xsky130_fd_sc_hs__o21ai_2_38 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__inv_4_23/Y sky130_fd_sc_hs__or2b_4_1/X
+ sky130_fd_sc_hs__nand2_2_15/B sky130_fd_sc_hs__o21ai_2_39/Y sky130_fd_sc_hs__o21ai_2_39/a_116_368#
+ sky130_fd_sc_hs__o21ai_2_39/a_27_74# sky130_fd_sc_hs__o21ai_2
Xsky130_fd_sc_hs__o21ai_2_49 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__inv_4_25/Y sky130_fd_sc_hs__or2b_4_1/X
+ sky130_fd_sc_hs__o21ai_2_51/A1 sky130_fd_sc_hs__buf_2_135/A sky130_fd_sc_hs__o21ai_2_49/a_116_368#
+ sky130_fd_sc_hs__o21ai_2_49/a_27_74# sky130_fd_sc_hs__o21ai_2
Xsky130_fd_sc_hs__buf_2_108 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__buf_2_109/A sky130_fd_sc_hs__buf_2_109/X
+ sky130_fd_sc_hs__buf_2_109/a_21_260# sky130_fd_sc_hs__buf_2
Xsky130_fd_sc_hs__buf_2_119 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__buf_2_119/A sky130_fd_sc_hs__buf_2_119/X
+ sky130_fd_sc_hs__buf_2_119/a_21_260# sky130_fd_sc_hs__buf_2
Xsky130_fd_sc_hs__conb_1_19 DVSS: DVDD: DVDD: DVSS: prbs_generator_syn_9/eqn[22] prbs_generator_syn_9/eqn[20]
+ sky130_fd_sc_hs__conb_1_19/a_165_290# sky130_fd_sc_hs__conb_1_19/a_21_290# sky130_fd_sc_hs__conb_1
Xsky130_fd_sc_hs__inv_4_15 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__inv_4_15/Y sky130_fd_sc_hs__inv_4_15/A
+ sky130_fd_sc_hs__inv_4
Xsky130_fd_sc_hs__inv_4_26 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__inv_4_27/Y osc_core_1/p1
+ sky130_fd_sc_hs__inv_4
Xsky130_fd_sc_hs__inv_4_37 DVSS: DVDD: DVDD: DVSS: osc_core_1/pi1_r[2] osc_core_1/pi1_l[2]
+ sky130_fd_sc_hs__inv_4
Xsky130_fd_sc_hs__inv_4_48 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__inv_4_49/Y osc_core_1/p3
+ sky130_fd_sc_hs__inv_4
Xsky130_fd_sc_hs__inv_4_59 DVSS: DVDD: DVDD: DVSS: osc_core_1/pi4_r[2] osc_core_1/pi4_l[2]
+ sky130_fd_sc_hs__inv_4
Xsky130_fd_sc_hs__conb_1_170 DVSS: DVDD: DVDD: DVSS: qr_4t1_mux_top_3/din_3_dummy
+ sky130_fd_sc_hs__conb_1_171/HI sky130_fd_sc_hs__conb_1_171/a_165_290# sky130_fd_sc_hs__conb_1_171/a_21_290#
+ sky130_fd_sc_hs__conb_1
Xsky130_fd_sc_hs__conb_1_181 DVSS: DVDD: DVDD: DVSS: prbs_generator_syn_23/eqn[28]
+ sky130_fd_sc_hs__conb_1_181/HI sky130_fd_sc_hs__conb_1_181/a_165_290# sky130_fd_sc_hs__conb_1_181/a_21_290#
+ sky130_fd_sc_hs__conb_1
Xsky130_fd_sc_hs__conb_1_192 DVSS: DVDD: DVDD: DVSS: prbs_generator_syn_19/eqn[13]
+ sky130_fd_sc_hs__conb_1_193/HI sky130_fd_sc_hs__conb_1_193/a_165_290# sky130_fd_sc_hs__conb_1_193/a_21_290#
+ sky130_fd_sc_hs__conb_1
Xsky130_fd_sc_hs__nand2_1_0 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__or2b_2_1/A sky130_fd_sc_hs__nor4_2_1/D
+ sky130_fd_sc_hs__nor2_4_1/Y sky130_fd_sc_hs__nand2_1_1/a_117_74# sky130_fd_sc_hs__nand2_1
Xsky130_fd_sc_hs__clkbuf_16_20 DVSS: DVDD: DVDD: DVSS: osc_core_1/pi1_l[2] sky130_fd_sc_hs__clkbuf_4_21/X
+ sky130_fd_sc_hs__clkbuf_16_21/a_114_74# sky130_fd_sc_hs__clkbuf_16
Xsky130_fd_sc_hs__clkbuf_16_31 DVSS: DVDD: DVDD: DVSS: osc_core_1/pi2_l[3] sky130_fd_sc_hs__clkbuf_8_1/X
+ sky130_fd_sc_hs__clkbuf_16_31/a_114_74# sky130_fd_sc_hs__clkbuf_16
Xsky130_fd_sc_hs__clkbuf_16_42 DVSS: DVDD: DVDD: DVSS: test_mux_misc sky130_fd_sc_hs__inv_4_39/Y
+ sky130_fd_sc_hs__clkbuf_16_43/a_114_74# sky130_fd_sc_hs__clkbuf_16
Xsky130_fd_sc_hs__clkbuf_16_53 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__clkbuf_16_53/X
+ sky130_fd_sc_hs__clkbuf_16_53/A sky130_fd_sc_hs__clkbuf_16_53/a_114_74# sky130_fd_sc_hs__clkbuf_16
Xsky130_fd_sc_hs__clkbuf_16_64 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__nand2_2_3/B
+ sky130_fd_sc_hs__or2b_2_5/X sky130_fd_sc_hs__clkbuf_16_65/a_114_74# sky130_fd_sc_hs__clkbuf_16
Xsky130_fd_sc_hs__clkbuf_16_75 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__clkbuf_16_75/X
+ sky130_fd_sc_hs__and2_4_1/X sky130_fd_sc_hs__clkbuf_16_75/a_114_74# sky130_fd_sc_hs__clkbuf_16
Xsky130_fd_sc_hs__clkbuf_16_86 DVSS: DVDD: DVDD: DVSS: hr_16t4_mux_top_1/clk sky130_fd_sc_hs__buf_1_1/X
+ sky130_fd_sc_hs__clkbuf_16_87/a_114_74# sky130_fd_sc_hs__clkbuf_16
Xsky130_fd_sc_hs__clkbuf_16_97 DVSS: DVDD: DVDD: DVSS: prbs_generator_syn_19/rst prbs_generator_syn_31/rst
+ sky130_fd_sc_hs__clkbuf_16_97/a_114_74# sky130_fd_sc_hs__clkbuf_16
Xsky130_fd_sc_hs__clkbuf_16_130 DVSS: DVDD: DVDD: DVSS: osc_core_1/pi4_l[3] pi4_con[3]
+ sky130_fd_sc_hs__clkbuf_16_131/a_114_74# sky130_fd_sc_hs__clkbuf_16
Xsky130_fd_sc_hs__nand2_2_16 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__nand2_2_17/Y
+ sky130_fd_sc_hs__or2b_2_3/A sky130_fd_sc_hs__nand2_2_27/B sky130_fd_sc_hs__nand2_2_17/a_27_74#
+ sky130_fd_sc_hs__nand2_2
Xsky130_fd_sc_hs__nand2_2_27 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__nand2_2_27/Y
+ sky130_fd_sc_hs__nand2_2_27/B sky130_fd_sc_hs__o21ai_4_1/A1 sky130_fd_sc_hs__nand2_2_27/a_27_74#
+ sky130_fd_sc_hs__nand2_2
Xprbs_generator_syn_5 prbs_generator_syn_9/clk prbs_generator_syn_9/rst prbs_generator_syn_5/cke
+ sky130_fd_sc_hs__conb_1_67/LO sky130_fd_sc_hs__conb_1_67/LO sky130_fd_sc_hs__conb_1_67/LO
+ sky130_fd_sc_hs__conb_1_67/LO sky130_fd_sc_hs__conb_1_67/LO sky130_fd_sc_hs__conb_1_67/LO
+ sky130_fd_sc_hs__conb_1_67/LO sky130_fd_sc_hs__conb_1_67/LO sky130_fd_sc_hs__conb_1_35/LO
+ sky130_fd_sc_hs__conb_1_35/LO sky130_fd_sc_hs__conb_1_35/LO sky130_fd_sc_hs__conb_1_35/HI
+ sky130_fd_sc_hs__conb_1_35/HI sky130_fd_sc_hs__conb_1_35/HI sky130_fd_sc_hs__conb_1_35/HI
+ sky130_fd_sc_hs__conb_1_35/HI sky130_fd_sc_hs__conb_1_35/HI sky130_fd_sc_hs__conb_1_35/HI
+ prbs_generator_syn_7/eqn[20] prbs_generator_syn_7/eqn[20] prbs_generator_syn_7/eqn[20]
+ prbs_generator_syn_7/eqn[20] prbs_generator_syn_7/eqn[20] sky130_fd_sc_hs__conb_1_69/HI
+ sky130_fd_sc_hs__conb_1_69/HI sky130_fd_sc_hs__conb_1_69/HI sky130_fd_sc_hs__conb_1_69/HI
+ prbs_generator_syn_7/cke prbs_generator_syn_7/cke prbs_generator_syn_7/cke prbs_generator_syn_7/cke
+ prbs_generator_syn_7/cke prbs_generator_syn_5/eqn[31] prbs_generator_syn_5/eqn[31]
+ prbs_generator_syn_5/eqn[31] prbs_generator_syn_5/eqn[31] prbs_generator_syn_5/eqn[31]
+ prbs_generator_syn_5/eqn[31] prbs_generator_syn_5/eqn[31] prbs_generator_syn_5/eqn[31]
+ prbs_generator_syn_5/eqn[23] prbs_generator_syn_5/eqn[23] prbs_generator_syn_5/eqn[23]
+ prbs_generator_syn_5/eqn[20] prbs_generator_syn_5/eqn[23] prbs_generator_syn_5/eqn[23]
+ prbs_generator_syn_5/eqn[23] prbs_generator_syn_5/eqn[23] prbs_generator_syn_5/eqn[23]
+ prbs_generator_syn_5/eqn[9] prbs_generator_syn_5/eqn[13] prbs_generator_syn_5/eqn[9]
+ prbs_generator_syn_5/eqn[9] prbs_generator_syn_5/eqn[9] prbs_generator_syn_5/eqn[9]
+ prbs_generator_syn_5/eqn[9] prbs_generator_syn_5/eqn[9] prbs_generator_syn_5/eqn[9]
+ prbs_generator_syn_5/eqn[5] prbs_generator_syn_5/eqn[5] prbs_generator_syn_5/eqn[5]
+ prbs_generator_syn_5/eqn[5] prbs_generator_syn_5/eqn[1] prbs_generator_syn_7/eqn[9]
+ prbs_generator_syn_9/inj_err sky130_fd_sc_hs__conb_1_35/LO sky130_fd_sc_hs__conb_1_35/LO
+ prbs_generator_syn_5/out DVSS: DVDD: prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_1/a_293_74#
+ prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_15/X prbs_generator_syn_5/sky130_fd_sc_hs__nand2_1_35/B
+ prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_51/Y prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_9/A
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_9/CLK prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_47/a_27_74#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_37/a_1226_296# prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_3/B
+ prbs_generator_syn_5/sky130_fd_sc_hs__nor2b_1_7/a_27_112# prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_29/B
+ prbs_generator_syn_5/sky130_fd_sc_hs__sdlclkp_2_1/a_580_74# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_1/a_1141_508#
+ prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_5/Y prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_41/a_230_79#
+ prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_61/a_138_385# prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_43/a_132_392#
+ prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_3/a_222_392# prbs_generator_syn_5/sky130_fd_sc_hs__nor2b_1_9/a_27_112#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_61/a_27_74# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_35/a_206_368#
+ prbs_generator_syn_5/sky130_fd_sc_hs__nand2_2_3/Y prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_25/B
+ prbs_generator_syn_5/sky130_fd_sc_hs__nand2_1_11/a_117_74# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_67/a_651_503#
+ prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_45/X prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_39/a_696_458#
+ prbs_generator_syn_5/sky130_fd_sc_hs__sdlclkp_2_1/a_1198_74# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_45/a_1034_424#
+ prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_17/a_222_392# prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_55/a_222_392#
+ prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_53/Y prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_35/A
+ prbs_generator_syn_5/m3_13600_1651# prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_59/a_52_123#
+ prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_5/a_293_74# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_35/a_1226_296#
+ prbs_generator_syn_5/sky130_fd_sc_hs__nand2_1_51/B prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_5/a_651_503#
+ prbs_generator_syn_5/sky130_fd_sc_hs__nand2_1_21/B prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_8/a_27_74#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_15/a_27_74# prbs_generator_syn_5/sky130_fd_sc_hs__and2b_2_1/X
+ prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_13/X prbs_generator_syn_5/sky130_fd_sc_hs__nand2_2_3/a_27_74#
+ prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_50/a_138_385# prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_33/a_132_392#
+ prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_1/a_376_368# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_25/a_206_368#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_35/a_437_503# prbs_generator_syn_5/sky130_fd_sc_hs__sdlclkp_2_1/a_708_451#
+ prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_45/a_230_79# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_29/a_696_458#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_32/a_27_74# prbs_generator_syn_5/sky130_fd_sc_hs__nor2b_1_4/Y
+ prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_59/a_293_74# prbs_generator_syn_5/sky130_fd_sc_hs__nand2_1_47/a_117_74#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_73/a_735_102# prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_21/a_112_119#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_23/a_1141_508# prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_25/a_293_74#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_7/Q prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_3/a_112_119#
+ prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_35/B prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_51/X
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_53/a_1178_124# prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_23/a_132_392#
+ prbs_generator_syn_5/sky130_fd_sc_hs__nand2_1_3/B prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_15/a_206_368#
+ prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_63/a_132_392# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_55/a_27_74#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_25/a_437_503# prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_41/a_52_123#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_47/a_651_503# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_73/a_1141_508#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_19/a_696_458# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_57/a_696_458#
+ prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_7/X prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_43/a_1034_424#
+ prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_55/A prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_11/a_112_119#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_21/a_1141_508# prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_35/a_222_392#
+ prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_49/a_230_79# prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_67/Y
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_71/a_27_74# prbs_generator_syn_5/sky130_fd_sc_hs__nand2_1_33/B
+ prbs_generator_syn_5/sky130_fd_sc_hs__conb_1_1/LO prbs_generator_syn_5/sky130_fd_sc_hs__nand2_1_19/a_117_74#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_51/a_1178_124# prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_33/X
+ prbs_generator_syn_5/sky130_fd_sc_hs__nand2_1_29/B prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_41/Y
+ prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_53/a_132_392# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_45/a_206_368#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_15/a_437_503# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_37/a_651_503#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_39/a_544_485# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_53/a_735_102#
+ prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_45/a_52_123# prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_1/B
+ prbs_generator_syn_5/sky130_fd_sc_hs__nand2_2_3/B prbs_generator_syn_5/sky130_fd_sc_hs__clkbuf_16_1/A
+ prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_21/X prbs_generator_syn_5/sky130_fd_sc_hs__nand2_1_25/B
+ prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_39/a_376_368# prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_63/X
+ prbs_generator_syn_5/m3_13600_3481# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_69/a_1178_124#
+ prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_21/a_138_385# prbs_generator_syn_5/sky130_fd_sc_hs__nor2b_1_8/Y
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_19/a_1178_124# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_49/a_27_74#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_45/a_437_503# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_27/a_651_503#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_71/a_1141_508# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_65/a_651_503#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_29/a_544_485# prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_3/a_138_385#
+ prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_55/X prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_43/a_735_102#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_41/a_1034_424# prbs_generator_syn_5/sky130_fd_sc_hs__nand2_1_9/B
+ prbs_generator_syn_5/sky130_fd_sc_hs__nor2b_1_9/Y prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_59/a_1034_424#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_39/a_1141_508# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_33/a_1226_296#
+ prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_49/a_52_123# prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_47/Y
+ prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_43/Y prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_4/a_651_503#
+ prbs_generator_syn_5/sky130_fd_sc_hs__nand2_1_49/B prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_19/A
+ prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_11/a_138_385# prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_5/X
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_63/a_206_368# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_17/a_651_503#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_19/a_544_485# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_55/a_651_503#
+ prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_9/Y prbs_generator_syn_5/sky130_fd_sc_hs__nand2_1_17/B
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_57/a_544_485# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_67/a_696_458#
+ prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_35/X prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_19/a_27_74#
+ prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_45/a_222_392# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_32/a_1226_296#
+ prbs_generator_syn_5/sky130_fd_sc_hs__nand2_1_43/B prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_25/A
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_1/a_206_368# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_49/a_1226_296#
+ prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_1/a_112_119# prbs_generator_syn_5/sky130_fd_sc_hs__or2_1_1/X
+ prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_59/a_376_368# prbs_generator_syn_5/sky130_fd_sc_hs__nand2_1_19/B
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_5/a_696_458# prbs_generator_syn_5/sky130_fd_sc_hs__nor2b_1_1/Y
+ prbs_generator_syn_5/sky130_fd_sc_hs__nor2b_1_5/a_278_368# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_17/a_1178_124#
+ prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_39/X prbs_generator_syn_5/m3_13600_5433#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_63/a_437_503# prbs_generator_syn_5/sky130_fd_sc_hs__nand2_2_5/B
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_23/a_735_102# prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_53/A
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_61/a_735_102# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_57/a_1034_424#
+ prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_63/B prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_37/a_1141_508#
+ prbs_generator_syn_5/sky130_fd_sc_hs__nand2_1_47/B prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_29/X
+ prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_65/Y prbs_generator_syn_5/m3_13600_4701#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_1/a_437_503# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_67/a_1178_124#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_9/a_735_102# prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_13/a_132_392#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_15/a_1178_124# prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_15/A
+ prbs_generator_syn_5/sky130_fd_sc_hs__nand2_1_1/B prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_43/B
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_35/a_651_503# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_8/D
+ prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_29/A prbs_generator_syn_5/sky130_fd_sc_hs__nand2_1_7/B
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_13/a_735_102# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_47/a_696_458#
+ prbs_generator_syn_5/sky130_fd_sc_hs__nand2_1_31/B prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_51/a_735_102#
+ prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_59/X prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_35/a_1141_508#
+ prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_25/a_222_392# prbs_generator_syn_5/sky130_fd_sc_hs__sdlclkp_2_1/a_288_48#
+ prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_55/B prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_17/B
+ prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_43/A prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_7/A
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_65/a_1178_124# prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_59/Y
+ prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_41/X prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_21/a_230_79#
+ prbs_generator_syn_5/sky130_fd_sc_hs__nand2_1_57/a_117_74# prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_1/a_222_392#
+ prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_19/B prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_35/a_293_74#
+ prbs_generator_syn_5/sky130_fd_sc_hs__nand2_1_23/a_117_74# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_73/a_206_368#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_25/a_651_503# prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_1/a_138_385#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_37/a_696_458# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_67/a_544_485#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_43/a_27_74# prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_9/X
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_55/a_1034_424# prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_39/a_112_119#
+ prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_15/a_222_392# prbs_generator_syn_5/sky130_fd_sc_hs__conb_1_1/HI
+ prbs_generator_syn_5/sky130_fd_sc_hs__nand2_1_23/B prbs_generator_syn_5/sky130_fd_sc_hs__nand2_1_53/B
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_9/a_1178_124# prbs_generator_syn_5/sky130_fd_sc_hs__nor2b_1_4/A
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_47/a_1226_296# prbs_generator_syn_5/m3_13600_11045#
+ prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_17/X prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_29/a_376_368#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_5/a_544_485# prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_3/X
+ prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_31/a_132_392# prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_61/A
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_15/a_651_503# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_73/a_437_503#
+ prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_25/a_230_79# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_27/a_696_458#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_65/a_696_458# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_33/a_735_102#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_71/a_735_102# prbs_generator_syn_5/m3_13600_7263#
+ prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_43/a_222_392# prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_50/Y
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_8/a_1178_124# prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_53/B
+ prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_19/a_376_368# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_63/a_1178_124#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_4/a_696_458# prbs_generator_syn_5/sky130_fd_sc_hs__nor2b_1_4/a_278_368#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_13/a_1178_124# prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_61/a_132_392#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_53/a_206_368# prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_21/a_52_123#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_45/a_651_503# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_17/a_696_458#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_47/a_544_485# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_55/a_696_458#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_21/a_735_102# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_37/a_27_74#
+ prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_61/B prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_61/X
+ prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_59/a_112_119# prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_31/A
+ prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_33/a_222_392# prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_29/a_230_79#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_45/a_1226_296# prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_9/a_132_392#
+ prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_5/A prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_57/Y
+ prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_31/X prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_51/a_27_74#
+ prbs_generator_syn_5/sky130_fd_sc_hs__nor2b_1_8/a_27_112# prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_47/a_376_368#
+ prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_53/a_293_74# prbs_generator_syn_5/sky130_fd_sc_hs__nand2_1_43/a_117_74#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_8/a_735_102# prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_21/a_293_74#
+ prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_39/a_138_385# prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_63/Y
+ prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_51/a_132_392# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_43/a_206_368#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_53/a_437_503# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_37/a_544_485#
+ prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_57/X prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_53/a_1034_424#
+ prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_25/a_52_123# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_33/a_1141_508#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_63/Q prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_23/a_222_392#
+ prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_63/a_222_392# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_7/a_1178_124#
+ prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_53/X prbs_generator_syn_5/sky130_fd_sc_hs__nand2_2_5/Y
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_61/a_1178_124# prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_1/a_230_79#
+ prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_43/a_230_79# prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_11/a_230_79#
+ prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_41/a_132_392# prbs_generator_syn_5/sky130_fd_sc_hs__nand2_1_13/a_117_74#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_43/a_437_503# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_27/a_544_485#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_63/a_651_503# prbs_generator_syn_5/sky130_fd_sc_hs__nand2_1_7/a_117_74#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_35/a_696_458# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_65/a_544_485#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_51/a_1034_424# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_41/a_735_102#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_32/a_1141_508# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_49/a_1141_508#
+ prbs_generator_syn_5/sky130_fd_sc_hs__nand2_1_55/B prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_53/a_222_392#
+ prbs_generator_syn_5/sky130_fd_sc_hs__sdlclkp_2_1/a_114_112# prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_9/a_293_74#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_43/a_1226_296# prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_29/a_52_123#
+ prbs_generator_syn_5/sky130_fd_sc_hs__nand2_1_37/B prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_1/a_651_503#
+ prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_27/a_376_368# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_4/a_544_485#
+ prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_67/a_376_368# prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_27/X
+ prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_1/X prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_59/a_138_385#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_29/a_1178_124# prbs_generator_syn_5/m3_13600_2871#
+ prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_5/a_230_79# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_23/a_206_368#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_61/a_206_368# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_17/a_544_485#
+ prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_15/a_230_79# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_25/a_696_458#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_55/a_544_485# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_32/a_735_102#
+ prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_29/a_293_74# prbs_generator_syn_5/sky130_fd_sc_hs__nand2_1_17/a_117_74#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_69/a_1034_424# prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_29/a_112_119#
+ prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_37/X prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_31/B
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_19/a_1034_424# prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_33/A
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_9/a_206_368# prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_57/a_376_368#
+ prbs_generator_syn_5/sky130_fd_sc_hs__sdlclkp_2_1/a_706_317# prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_11/B
+ prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_1/a_52_123# prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_39/B
+ prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_21/a_132_392# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_13/a_206_368#
+ prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_43/a_52_123# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_51/a_206_368#
+ prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_47/X prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_23/a_437_503#
+ prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_11/a_52_123# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_61/a_437_503#
+ prbs_generator_syn_5/sky130_fd_sc_hs__nor2b_1_7/Y prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_51/A
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_15/a_696_458# prbs_generator_syn_5/sky130_fd_sc_hs__nor2b_1_5/Y
+ prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_9/a_230_79# prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_25/X
+ prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_19/a_112_119# prbs_generator_syn_5/sky130_fd_sc_hs__nand2_1_45/B
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_5/a_1178_124# prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_19/a_230_79#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_41/a_1226_296# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_59/a_1226_296#
+ prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_63/a_230_79# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_51/Q
+ prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_7/a_132_392# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_9/a_437_503#
+ prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_46/a_376_368# prbs_generator_syn_5/sky130_fd_sc_hs__nand2_1_33/a_117_74#
+ prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_11/a_293_74# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_27/a_1178_124#
+ prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_11/a_132_392# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_13/a_437_503#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_51/a_437_503# prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_5/a_52_123#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_35/a_544_485# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_73/a_651_503#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_45/a_696_458# prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_15/a_52_123#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_47/a_1141_508# prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_47/a_112_119#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_4/a_1178_124# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_17/a_1034_424#
+ prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_23/B prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_37/a_376_368#
+ prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_15/B prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_7/Y
+ prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_29/a_138_385# prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_33/a_230_79#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_25/a_1178_124# prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_47/a_293_74#
+ prbs_generator_syn_5/sky130_fd_sc_hs__nand2_1_37/a_117_74# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_33/a_206_368#
+ prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_15/a_293_74# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_71/a_206_368#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_25/a_544_485# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_67/a_1034_424#
+ prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_13/a_222_392# prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_9/a_52_123#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_15/a_1034_424# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_57/a_1226_296#
+ prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_19/a_52_123# prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_23/X
+ prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_63/a_52_123# prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_19/a_138_385#
+ prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_9/a_376_368# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_21/a_206_368#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_33/a_437_503# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_71/a_437_503#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_53/a_651_503# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_15/a_544_485#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_63/a_696_458# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_65/a_1034_424#
+ prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_19/a_293_74# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_45/a_1141_508#
+ prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_27/a_112_119# prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_67/a_112_119#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_1/a_1178_124# prbs_generator_syn_5/sky130_fd_sc_hs__conb_1_1/a_21_290#
+ prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_63/a_293_74# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_8/a_206_368#
+ prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_17/a_376_368# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_63/a_27_74#
+ prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_21/A prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_55/a_376_368#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_1/a_696_458# prbs_generator_syn_5/sky130_fd_sc_hs__nor2b_1_1/a_278_368#
+ prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_47/a_138_385# prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_33/a_52_123#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_9/a_1034_424# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_21/a_437_503#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_1/a_27_74# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_43/a_651_503#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_1/Q prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_45/a_544_485#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_69/a_735_102# prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_57/a_112_119#
+ prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_31/a_222_392# prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_13/A
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_55/a_1226_296# prbs_generator_syn_5/sky130_fd_sc_hs__nand2_2_5/a_27_74#
+ prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_53/a_230_79# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_8/a_437_503#
+ prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_67/a_293_74# prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_33/a_293_74#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_7/a_735_102# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_23/a_1178_124#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_41/a_206_368# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_8/a_1034_424#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_63/a_1034_424# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_59/a_735_102#
+ prbs_generator_syn_5/sky130_fd_sc_hs__nand2_1_5/B prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_43/a_1141_508#
+ prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_46/a_112_119# prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_61/a_222_392#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_13/a_1034_424# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_73/a_1178_124#
+ prbs_generator_syn_5/sky130_fd_sc_hs__nand2_1_27/B prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_13/B
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_57/a_27_74# prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_57/a_230_79#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_21/a_1178_124# prbs_generator_syn_5/sky130_fd_sc_hs__nor2b_1_1/a_27_112#
+ prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_27/a_138_385# prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_23/a_230_79#
+ prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_67/a_138_385# prbs_generator_syn_5/sky130_fd_sc_hs__nand2_1_41/B
+ prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_9/a_222_392# prbs_generator_syn_5/sky130_fd_sc_hs__nand2_1_27/a_117_74#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_32/a_206_368# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_23/a_651_503#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_41/a_437_503# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_73/a_27_74#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_61/a_651_503# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_63/a_544_485#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_49/a_735_102# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_73/a_696_458#
+ prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_37/a_112_119# prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_51/a_222_392#
+ prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_43/X prbs_generator_syn_5/sky130_fd_sc_hs__nand2_2_1/B
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_9/a_651_503# prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_53/a_52_123#
+ prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_49/X prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_25/a_376_368#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_1/a_544_485# prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_65/a_376_368#
+ prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_57/a_138_385# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_27/a_27_74#
+ prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_39/a_132_392# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_7/a_1034_424#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_13/a_651_503# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_32/a_437_503#
+ prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_27/a_230_79# prbs_generator_syn_5/m3_13600_12265#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_51/a_651_503# prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_59/B
+ prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_47/A prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_61/a_1034_424#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_41/a_1141_508# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_59/a_1141_508#
+ prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_41/a_222_392# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_53/a_1226_296#
+ prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_3/A prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_71/a_1178_124#
+ prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_9/a_112_119# prbs_generator_syn_5/sky130_fd_sc_hs__nand2_1_3/a_117_74#
+ prbs_generator_syn_5/m3_13600_8483# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_39/a_1178_124#
+ prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_57/a_52_123# prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_46/a_138_385#
+ prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_23/a_52_123# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_67/a_27_74#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_53/a_696_458# prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_17/a_112_119#
+ prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_11/A prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_55/a_112_119#
+ prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_1/A prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_51/a_1226_296#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_29/a_1034_424# prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_59/A
+ prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_23/A prbs_generator_syn_5/sky130_fd_sc_hs__nand2_1_39/B
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_5/a_27_74# prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_57/a_293_74#
+ prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_37/a_138_385# prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_59/a_132_392#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_33/a_651_503# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_71/a_651_503#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_43/a_696_458# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_73/a_544_485#
+ prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_27/a_52_123# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_57/a_1141_508#
+ prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_21/a_222_392# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_35/a_27_74#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_69/a_1226_296# prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_37/B
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_19/a_1226_296# prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_35/a_376_368#
+ prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_47/a_230_79# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_37/a_1178_124#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_5/a_1034_424# prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_49/a_132_392#
+ prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_7/a_222_392# prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_27/a_293_74#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_21/a_651_503# prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_9/a_138_385#
+ prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_11/a_222_392# prbs_generator_syn_5/m3_13600_14095#
+ prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_50/A prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_27/a_1034_424#
+ prbs_generator_syn_5/sky130_fd_sc_hs__nand2_1_13/B prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_8/a_651_503#
+ prbs_generator_syn_5/m3_13600_9703# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_35/a_1178_124#
+ prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_17/a_138_385# prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_55/a_138_385#
+ prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_7/a_230_79# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_4/a_1034_424#
+ prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_7/a_376_368# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_69/a_206_368#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_23/a_696_458# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_53/a_544_485#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_39/a_735_102# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_61/a_696_458#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_55/a_1141_508# prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_25/a_112_119#
+ prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_65/a_112_119# prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_43/a_293_74#
+ prbs_generator_syn_5/sky130_fd_sc_hs__nand2_1_57/B prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_25/a_1034_424#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_7/a_206_368# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_17/a_1226_296#
+ prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_15/a_376_368# prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_53/a_376_368#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_9/a_696_458# prbs_generator_syn_5/m3_13600_431#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_45/a_27_74# prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_47/a_52_123#
+ prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_29/a_132_392# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_59/a_206_368#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_69/a_437_503# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_41/a_651_503#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_43/a_544_485# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_13/a_696_458#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_29/a_735_102# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_51/a_696_458#
+ prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_61/Y prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_67/a_1226_296#
+ prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_5/a_132_392# prbs_generator_syn_5/sky130_fd_sc_hs__and2b_2_1/a_198_48#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_7/a_437_503# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_15/a_1226_296#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_69/a_27_74# prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_46/a_293_74#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_1/a_1034_424# prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_19/a_132_392#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_49/a_206_368# prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_7/a_52_123#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_59/a_437_503# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_32/a_651_503#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_7/a_27_74# prbs_generator_syn_5/sky130_fd_sc_hs__nand2_2_1/a_27_74#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_19/a_735_102# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_57/a_735_102#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_65/a_1226_296# prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_37/A
+ prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_33/a_376_368# prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_37/a_230_79#
+ prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_25/a_138_385# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_39/a_27_74#
+ prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_65/a_138_385# prbs_generator_syn_5/sky130_fd_sc_hs__nor2b_1_9/a_278_368#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_49/a_437_503# prbs_generator_syn_5/sky130_fd_sc_hs__and2b_2_1/a_505_74#
+ prbs_generator_syn_5/sky130_fd_sc_hs__nand2_1_51/a_117_74# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_23/a_544_485#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_33/a_696_458# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_61/a_544_485#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_9/a_1226_296# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_53/a_1141_508#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_71/a_696_458# prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_35/a_112_119#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_23/a_1034_424# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_9/a_544_485#
+ prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_63/a_376_368# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_33/a_1178_124#
+ prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_5/a_376_368# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_13/a_544_485#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_73/a_1034_424# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_21/a_696_458#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_51/a_544_485# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_8/a_1226_296#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_51/a_1141_508# prbs_generator_syn_5/sky130_fd_sc_hs__nand2_1_55/a_117_74#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_21/a_1034_424# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_63/a_1226_296#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_23/a_27_74# prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_7/a_112_119#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_13/a_1226_296# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_8/a_696_458#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_32/a_1178_124# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_49/a_1178_124#
+ prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_37/a_52_123# prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_27/a_132_392#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_71/Q prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_67/a_735_102#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_69/a_1141_508# prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_15/a_112_119#
+ prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_53/a_112_119# prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_39/a_222_392#
+ prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_55/a_230_79# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_19/a_1141_508#
+ prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_37/a_293_74# prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_43/a_376_368#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_5/a_735_102# prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_35/a_138_385#
+ prbs_generator_syn_5/sky130_fd_sc_hs__sdlclkp_2_1/a_114_424# prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_57/a_132_392#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_71/a_1034_424# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_7/a_1226_296#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_33/a_544_485# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_41/a_696_458#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_71/a_544_485# prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_21/B
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_61/a_1226_296# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_39/a_1034_424#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_17/a_27_74# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_9/a_27_74#
+ prbs_generator_syn_5/sky130_fd_sc_hs__nor2b_1_5/a_27_112# prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_47/a_132_392#
+ prbs_generator_syn_5/sky130_fd_sc_hs__nor2b_1_8/a_278_368# prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_9/B
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_39/a_206_368# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_33/a_27_74#
+ prbs_generator_syn_5/sky130_fd_sc_hs__nand2_1_41/a_117_74# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_69/a_651_503#
+ prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_51/a_293_74# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_21/a_544_485#
+ prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_7/a_138_385# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_32/a_696_458#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_47/a_735_102# prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_33/a_112_119#
+ prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_59/a_222_392# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_17/a_1141_508#
+ prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_55/a_52_123# prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_3/a_293_74#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_7/a_651_503# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_29/a_1226_296#
+ prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_23/a_376_368# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_8/a_544_485#
+ prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_47/B prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_47/a_1178_124#
+ prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_15/a_138_385# prbs_generator_syn_5/sky130_fd_sc_hs__sdlclkp_2_1/a_1195_374#
+ prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_53/a_138_385# prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_37/a_132_392#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_29/a_206_368# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_39/a_437_503#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_59/a_651_503# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_37/a_735_102#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_67/a_1141_508# prbs_generator_syn_5/sky130_fd_sc_hs__and2b_2_1/a_27_74#
+ prbs_generator_syn_5/sky130_fd_sc_hs__conb_1_1/a_165_290# prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_55/a_293_74#
+ prbs_generator_syn_5/sky130_fd_sc_hs__nand2_1_45/a_117_74# prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_63/a_112_119#
+ prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_49/a_222_392# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_37/a_1034_424#
+ prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_23/a_293_74# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_15/a_1141_508#
+ prbs_generator_syn_5/sky130_fd_sc_hs__nand2_1_5/a_117_74# prbs_generator_syn_5/m3_13600_13485#
+ prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_5/a_112_119# prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_13/a_376_368#
+ prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_51/a_376_368# prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_7/a_293_74#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_19/a_206_368# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_57/a_206_368#
+ prbs_generator_syn_5/sky130_fd_sc_hs__sdlclkp_2_1/a_318_74# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_29/a_437_503#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_49/a_651_503# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_25/a_27_74#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_5/a_1226_296# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_41/a_544_485#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_27/a_735_102# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_65/a_1141_508#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_65/a_735_102# prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_3/a_230_79#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_35/a_1034_424# prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_13/a_230_79#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_41/a_27_74# prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_3/a_132_392#
+ prbs_generator_syn_5/sky130_fd_sc_hs__nand2_1_49/a_117_74# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_27/a_1226_296#
+ prbs_generator_syn_5/sky130_fd_sc_hs__nand2_1_15/a_117_74# prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_41/a_376_368#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_45/a_1178_124# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_4/a_735_102#
+ prbs_generator_syn_5/sky130_fd_sc_hs__nand2_1_9/a_117_74# prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_33/a_138_385#
+ prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_17/a_132_392# prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_55/a_132_392#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_9/a_1141_508# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_19/a_437_503#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_57/a_437_503# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_4/a_1226_296#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_32/a_544_485# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_17/a_735_102#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_55/a_735_102# prbs_generator_syn_5/m3_13600_2261#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_65/a_27_74# prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_29/a_222_392#
+ prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_43/a_112_119# prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_19/X
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_25/a_1226_296# prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_31/a_376_368#
+ prbs_generator_syn_5/sky130_fd_sc_hs__or2_1_1/a_63_368# prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_17/a_230_79#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_4/a_27_74# prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_61/a_230_79#
+ prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_63/a_138_385# prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_5/a_222_392#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_8/a_1141_508# prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_41/a_293_74#
+ prbs_generator_syn_5/sky130_fd_sc_hs__nand2_1_31/a_117_74# prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_5/a_138_385#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_63/a_1141_508# prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_19/a_222_392#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_13/a_1141_508# prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_3/a_52_123#
+ prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_13/a_52_123# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_43/a_1178_124#
+ prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_61/a_376_368# prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_35/a_132_392#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_67/a_206_368# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_1/a_1226_296#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_69/a_696_458# prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_31/a_230_79#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_35/a_735_102# prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_23/a_112_119#
+ prbs_generator_syn_5/sky130_fd_sc_hs__nand2_1_35/a_117_74# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_59/a_27_74#
+ prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_13/a_293_74# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_5/a_206_368#
+ prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_50/a_376_368# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_7/a_696_458#
+ prbs_generator_syn_5/sky130_fd_sc_hs__nor2b_1_7/a_278_368# prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_17/a_52_123#
+ prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_43/a_138_385# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_7/a_1141_508#
+ prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_61/a_52_123# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_67/a_437_503#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_61/a_1141_508# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_25/a_735_102#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_59/a_696_458# prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_13/a_112_119#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_33/a_1034_424# prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_51/a_112_119#
+ prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_35/a_230_79# prbs_generator_syn_5/m3_13600_4091#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_23/a_1226_296# prbs_generator_syn_5/sky130_fd_sc_hs__nand2_1_39/a_117_74#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_29/a_27_74# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_5/a_437_503#
+ prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_17/a_293_74# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_41/a_1178_124#
+ prbs_generator_syn_5/sky130_fd_sc_hs__or2_1_1/a_152_368# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_59/a_1178_124#
+ prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_61/a_293_74# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_47/a_206_368#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_39/a_651_503# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_49/a_696_458#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_15/a_735_102# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_32/a_1034_424#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_73/a_1226_296# prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_27/a_222_392#
+ prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_41/a_112_119# prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_31/a_52_123#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_49/a_1034_424# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_29/a_1141_508#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_21/a_1226_296# prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_39/a_230_79#
+ prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_23/a_138_385# prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_51/a_230_79#
+ prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_45/a_132_392# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_37/a_206_368#
+ prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_65/a_293_74# prbs_generator_syn_5/sky130_fd_sc_hs__nand2_1_53/a_117_74#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_47/a_437_503# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_29/a_651_503#
+ prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_31/a_293_74# prbs_generator_syn_5/sky130_fd_sc_hs__nand2_1_21/a_117_74#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_69/a_544_485# prbs_generator_syn_5/sky130_fd_sc_hs__clkbuf_16_1/a_114_74#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_45/a_735_102# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_13/a_27_74#
+ prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_31/a_112_119# prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_57/a_222_392#
+ prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_35/a_52_123# prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_21/a_376_368#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_7/a_544_485# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_57/a_1178_124#
+ prbs_generator_syn_5/m3_13600_6043# prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_13/a_138_385#
+ prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_51/a_138_385# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_5/a_1141_508#
+ prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_3/a_376_368# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_27/a_206_368#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_65/a_206_368# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_37/a_437_503#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_19/a_651_503# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_57/a_651_503#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_59/a_544_485# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_71/a_1226_296#
+ prbs_generator_syn_5/sky130_fd_sc_hs__nand2_1_25/a_117_74# prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_61/a_112_119#
+ prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_47/a_222_392# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_27/a_1141_508#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_53/a_27_74# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_4/a_206_368#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_39/a_1226_296# prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_11/a_376_368#
+ prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_39/a_52_123# prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_41/a_138_385#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_4/a_1141_508# prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_25/a_132_392#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_17/a_206_368# prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_41/A
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_55/a_206_368# prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_51/a_52_123#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_27/a_437_503# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_65/a_437_503#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_49/a_544_485# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_63/a_735_102#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_47/a_1034_424# prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_50/a_112_119#
+ prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_37/a_222_392# prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_59/a_230_79#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_25/a_1141_508# prbs_generator_syn_5/sky130_fd_sc_hs__nor2b_1_4/a_27_112#
+ prbs_generator_syn_5/sky130_fd_sc_hs__sdlclkp_2_1/a_685_81# prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_1/a_132_392#
+ prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_39/a_293_74# prbs_generator_syn_5/sky130_fd_sc_hs__nand2_1_29/a_117_74#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_4/a_437_503# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_55/a_1178_124#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_21/a_27_74# prbs_generator_syn_5/m3_13600_12875#
+ prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_50/a_293_74# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_1/a_735_102#
+ prbs_generator_syn_5/sky130_fd_sc_hs__xnor2_1_31/a_138_385# prbs_generator_syn_5/sky130_fd_sc_hs__a22o_1_15/a_132_392#
+ prbs_generator_syn_5/sky130_fd_sc_hs__nand2_1_1/a_117_74# prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_17/a_437_503#
+ prbs_generator_syn_5/sky130_fd_sc_hs__dfxtp_4_55/a_437_503# prbs_generator_syn
Xsky130_fd_sc_hs__clkbuf_4_130 DVSS: DVDD: DVDD: DVSS: pi5_con[2] sky130_fd_sc_hs__clkbuf_4_131/X
+ sky130_fd_sc_hs__clkbuf_4_131/a_83_270# sky130_fd_sc_hs__clkbuf_4
Xsky130_fd_sc_hs__clkdlyinv5sd2_1_4 DVSS: DVDD: DVSS: DVDD: dout_n sky130_fd_sc_hs__and2_2_1/B
+ sky130_fd_sc_hs__clkdlyinv5sd2_1_5/a_28_74# sky130_fd_sc_hs__clkdlyinv5sd2_1_5/a_682_74#
+ sky130_fd_sc_hs__clkdlyinv5sd2_1_5/a_549_74# sky130_fd_sc_hs__clkdlyinv5sd2_1_5/a_288_74#
+ sky130_fd_sc_hs__clkdlyinv5sd2_1
Xsky130_fd_sc_hs__clkbuf_4_70 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__nand2_2_5/Y
+ sky130_fd_sc_hs__inv_4_11/A sky130_fd_sc_hs__clkbuf_4_71/a_83_270# sky130_fd_sc_hs__clkbuf_4
Xsky130_fd_sc_hs__clkbuf_4_81 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__nand2_8_1/Y
+ sky130_fd_sc_hs__clkbuf_4_81/X sky130_fd_sc_hs__clkbuf_4_81/a_83_270# sky130_fd_sc_hs__clkbuf_4
Xsky130_fd_sc_hs__clkbuf_4_92 DVSS: DVDD: DVDD: DVSS: div_ratio_half[3] sky130_fd_sc_hs__clkbuf_4_93/X
+ sky130_fd_sc_hs__clkbuf_4_93/a_83_270# sky130_fd_sc_hs__clkbuf_4
Xsky130_fd_sc_hs__o21ai_2_17 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__inv_4_17/Y sky130_fd_sc_hs__or2b_4_5/X
+ sky130_fd_sc_hs__nand2_2_7/A sky130_fd_sc_hs__o21ai_2_17/Y sky130_fd_sc_hs__o21ai_2_17/a_116_368#
+ sky130_fd_sc_hs__o21ai_2_17/a_27_74# sky130_fd_sc_hs__o21ai_2
Xsky130_fd_sc_hs__o21ai_2_28 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__inv_4_21/Y sky130_fd_sc_hs__or2b_4_1/A
+ sky130_fd_sc_hs__buf_8_3/X sky130_fd_sc_hs__buf_2_95/A sky130_fd_sc_hs__o21ai_2_29/a_116_368#
+ sky130_fd_sc_hs__o21ai_2_29/a_27_74# sky130_fd_sc_hs__o21ai_2
Xsky130_fd_sc_hs__o21ai_2_39 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__inv_4_23/Y sky130_fd_sc_hs__or2b_4_1/X
+ sky130_fd_sc_hs__nand2_2_15/B sky130_fd_sc_hs__o21ai_2_39/Y sky130_fd_sc_hs__o21ai_2_39/a_116_368#
+ sky130_fd_sc_hs__o21ai_2_39/a_27_74# sky130_fd_sc_hs__o21ai_2
Xqr_4t1_mux_top_0 qr_4t1_mux_top_1/clk_Q hr_16t4_mux_top_1/clk qr_4t1_mux_top_3/clk_I
+ qr_4t1_mux_top_1/clk_IB qr_4t1_mux_top_1/din[3] qr_4t1_mux_top_1/din[2] qr_4t1_mux_top_1/din[1]
+ qr_4t1_mux_top_1/din[0] qr_4t1_mux_top_1/rst qr_4t1_mux_top_1/din_3_dummy qr_4t1_mux_top_1/din_3_dummy
+ qr_4t1_mux_top_1/din_3_dummy qr_4t1_mux_top_1/din_3_dummy dout_p qr_4t1_mux_top_1/mux_out_dummy
+ DVSS: DVDD: qr_4t1_mux_top_1/sky130_fd_sc_hs__dfxtp_2_1/a_1172_124# qr_4t1_mux_top_1/sky130_fd_sc_hs__dfxtp_2_3/a_1217_314#
+ qr_4t1_mux_top_1/sky130_fd_sc_hs__dfxtp_4_1/a_1141_508# qr_4t1_mux_top_1/sky130_fd_sc_hs__dfxtp_2_3/a_695_459#
+ qr_4t1_mux_top_1/sky130_fd_sc_hs__dfxtp_4_3/a_651_503# qr_4t1_mux_top_1/sky130_fd_sc_hs__dfxtp_2_1/a_538_429#
+ qr_4t1_mux_top_1/sky130_fd_sc_hs__mux4_1_1/A0 qr_4t1_mux_top_1/sky130_fd_sc_hs__mux4_1_1/a_264_74#
+ qr_4t1_mux_top_1/sky130_fd_sc_hs__dfxtp_2_1/a_1217_314# qr_4t1_mux_top_1/sky130_fd_sc_hs__mux4_1_1/a_1338_125#
+ qr_4t1_mux_top_1/sky130_fd_sc_hs__mux4_4_1/a_758_306# qr_4t1_mux_top_1/sky130_fd_sc_hs__mux4_1_1/A2
+ qr_4t1_mux_top_1/sky130_fd_sc_hs__dfxtp_2_7/a_206_368# qr_4t1_mux_top_1/sky130_fd_sc_hs__dfxtp_2_5/a_431_508#
+ qr_4t1_mux_top_1/sky130_fd_sc_hs__mux4_1_1/A1 qr_4t1_mux_top_1/sky130_fd_sc_hs__dfxtp_2_7/D
+ qr_4t1_mux_top_1/sky130_fd_sc_hs__dfxtp_4_1/a_206_368# qr_4t1_mux_top_1/sky130_fd_sc_hs__dfxtp_2_7/a_708_101#
+ qr_4t1_mux_top_1/sky130_fd_sc_hs__dfxtp_4_3/a_696_458# qr_4t1_mux_top_1/sky130_fd_sc_hs__dfxtp_2_9/a_644_504#
+ qr_4t1_mux_top_1/sky130_fd_sc_hs__mux4_1_1/X qr_4t1_mux_top_1/sky130_fd_sc_hs__dfxtp_2_11/a_206_368#
+ qr_4t1_mux_top_1/sky130_fd_sc_hs__dfxtp_4_1/a_437_503# qr_4t1_mux_top_1/sky130_fd_sc_hs__clkbuf_1_1/a_27_74#
+ qr_4t1_mux_top_1/sky130_fd_sc_hs__dfxtp_2_3/a_431_508# qr_4t1_mux_top_1/sky130_fd_sc_hs__dfxtp_4_3/a_544_485#
+ qr_4t1_mux_top_1/sky130_fd_sc_hs__dfxtp_2_9/a_538_429# qr_4t1_mux_top_1/sky130_fd_sc_hs__dfxtp_2_11/a_708_101#
+ qr_4t1_mux_top_1/sky130_fd_sc_hs__dfxtp_2_11/a_1125_508# qr_4t1_mux_top_1/sky130_fd_sc_hs__mux4_1_1/a_27_74#
+ qr_4t1_mux_top_1/sky130_fd_sc_hs__mux4_1_1/a_342_74# qr_4t1_mux_top_1/sky130_fd_sc_hs__dfxtp_2_11/a_27_74#
+ qr_4t1_mux_top_1/sky130_fd_sc_hs__dfxtp_2_1/a_695_459# qr_4t1_mux_top_1/sky130_fd_sc_hs__dfxtp_4_1/a_651_503#
+ qr_4t1_mux_top_1/sky130_fd_sc_hs__dfxtp_4_1/D qr_4t1_mux_top_1/sky130_fd_sc_hs__dfxtp_2_7/a_644_504#
+ qr_4t1_mux_top_1/sky130_fd_sc_hs__dfxtp_4_3/a_1178_124# qr_4t1_mux_top_1/sky130_fd_sc_hs__clkbuf_2_1/a_43_192#
+ qr_4t1_mux_top_1/sky130_fd_sc_hs__dfxtp_2_5/a_206_368# qr_4t1_mux_top_1/sky130_fd_sc_hs__clkbuf_1_5/X
+ qr_4t1_mux_top_1/sky130_fd_sc_hs__dfxtp_2_9/a_1125_508# qr_4t1_mux_top_1/sky130_fd_sc_hs__clkbuf_2_3/X
+ qr_4t1_mux_top_1/sky130_fd_sc_hs__dfxtp_2_7/a_538_429# qr_4t1_mux_top_1/sky130_fd_sc_hs__dfxtp_2_9/Q
+ qr_4t1_mux_top_1/sky130_fd_sc_hs__dfxtp_4_1/a_1178_124# qr_4t1_mux_top_1/sky130_fd_sc_hs__dfxtp_2_11/a_644_504#
+ qr_4t1_mux_top_1/sky130_fd_sc_hs__dfxtp_4_1/a_696_458# qr_4t1_mux_top_1/sky130_fd_sc_hs__dfxtp_2_5/a_27_74#
+ qr_4t1_mux_top_1/sky130_fd_sc_hs__dfxtp_2_5/a_708_101# qr_4t1_mux_top_1/sky130_fd_sc_hs__dfxtp_4_1/a_27_74#
+ qr_4t1_mux_top_1/sky130_fd_sc_hs__mux4_4_1/a_1285_377# qr_4t1_mux_top_1/sky130_fd_sc_hs__dfxtp_2_7/a_1125_508#
+ qr_4t1_mux_top_1/sky130_fd_sc_hs__mux4_1_1/a_537_341# qr_4t1_mux_top_1/sky130_fd_sc_hs__mux4_1_1/a_255_341#
+ qr_4t1_mux_top_1/sky130_fd_sc_hs__mux4_4_1/A0 qr_4t1_mux_top_1/sky130_fd_sc_hs__clkbuf_1_3/X
+ qr_4t1_mux_top_1/sky130_fd_sc_hs__mux4_1_1/A3 qr_4t1_mux_top_1/sky130_fd_sc_hs__dfxtp_2_11/a_538_429#
+ qr_4t1_mux_top_1/sky130_fd_sc_hs__dfxtp_2_3/a_206_368# qr_4t1_mux_top_1/sky130_fd_sc_hs__dfxtp_2_1/a_431_508#
+ qr_4t1_mux_top_1/sky130_fd_sc_hs__clkbuf_1_1/X qr_4t1_mux_top_1/sky130_fd_sc_hs__dfxtp_2_9/a_695_459#
+ qr_4t1_mux_top_1/sky130_fd_sc_hs__dfxtp_4_1/a_544_485# qr_4t1_mux_top_1/sky130_fd_sc_hs__dfxtp_2_5/a_1125_508#
+ qr_4t1_mux_top_1/sky130_fd_sc_hs__mux4_4_1/A2 qr_4t1_mux_top_1/sky130_fd_sc_hs__dfxtp_2_7/a_27_74#
+ qr_4t1_mux_top_1/sky130_fd_sc_hs__dfxtp_2_3/a_708_101# qr_4t1_mux_top_1/sky130_fd_sc_hs__dfxtp_2_3/a_1125_508#
+ qr_4t1_mux_top_1/sky130_fd_sc_hs__dfxtp_4_3/a_27_74# qr_4t1_mux_top_1/sky130_fd_sc_hs__dfxtp_2_11/a_1019_424#
+ qr_4t1_mux_top_1/sky130_fd_sc_hs__mux4_1_1/a_450_74# qr_4t1_mux_top_1/sky130_fd_sc_hs__dfxtp_4_3/a_1034_424#
+ qr_4t1_mux_top_1/sky130_fd_sc_hs__clkbuf_1_3/a_27_74# qr_4t1_mux_top_1/sky130_fd_sc_hs__dfxtp_2_1/a_1125_508#
+ qr_4t1_mux_top_1/sky130_fd_sc_hs__mux4_4_1/a_114_126# qr_4t1_mux_top_1/sky130_fd_sc_hs__dfxtp_2_1/a_27_74#
+ qr_4t1_mux_top_1/sky130_fd_sc_hs__dfxtp_2_5/a_644_504# qr_4t1_mux_top_1/sky130_fd_sc_hs__dfxtp_4_1/a_1034_424#
+ qr_4t1_mux_top_1/sky130_fd_sc_hs__dfxtp_2_11/a_1172_124# qr_4t1_mux_top_1/sky130_fd_sc_hs__mux4_4_1/a_1450_121#
+ qr_4t1_mux_top_1/sky130_fd_sc_hs__dfxtp_2_9/a_431_508# qr_4t1_mux_top_1/sky130_fd_sc_hs__dfxtp_2_7/a_695_459#
+ qr_4t1_mux_top_1/sky130_fd_sc_hs__mux4_4_1/a_1191_121# qr_4t1_mux_top_1/sky130_fd_sc_hs__mux4_1_1/a_768_74#
+ qr_4t1_mux_top_1/sky130_fd_sc_hs__dfxtp_2_5/a_538_429# qr_4t1_mux_top_1/sky130_fd_sc_hs__dfxtp_2_9/a_1019_424#
+ qr_4t1_mux_top_1/sky130_fd_sc_hs__mux4_1_1/a_1396_99# qr_4t1_mux_top_1/sky130_fd_sc_hs__dfxtp_2_3/a_644_504#
+ qr_4t1_mux_top_1/sky130_fd_sc_hs__mux4_1_1/a_1065_387# qr_4t1_mux_top_1/sky130_fd_sc_hs__dfxtp_4_3/a_735_102#
+ qr_4t1_mux_top_1/sky130_fd_sc_hs__dfxtp_2_3/a_27_74# qr_4t1_mux_top_1/sky130_fd_sc_hs__dfxtp_2_11/a_695_459#
+ qr_4t1_mux_top_1/sky130_fd_sc_hs__dfxtp_2_11/a_1217_314# qr_4t1_mux_top_1/sky130_fd_sc_hs__dfxtp_2_7/a_1019_424#
+ qr_4t1_mux_top_1/sky130_fd_sc_hs__dfxtp_2_1/a_206_368# qr_4t1_mux_top_1/sky130_fd_sc_hs__mux4_4_1/a_1278_121#
+ qr_4t1_mux_top_1/sky130_fd_sc_hs__dfxtp_2_3/a_538_429# qr_4t1_mux_top_1/sky130_fd_sc_hs__dfxtp_4_3/a_1226_296#
+ qr_4t1_mux_top_1/sky130_fd_sc_hs__dfxtp_2_1/a_708_101# qr_4t1_mux_top_1/sky130_fd_sc_hs__dfxtp_2_9/a_1172_124#
+ qr_4t1_mux_top_1/sky130_fd_sc_hs__mux4_4_1/a_509_392# qr_4t1_mux_top_1/sky130_fd_sc_hs__dfxtp_2_5/a_1019_424#
+ qr_4t1_mux_top_1/sky130_fd_sc_hs__dfxtp_2_3/a_1019_424# qr_4t1_mux_top_1/sky130_fd_sc_hs__dfxtp_2_7/a_431_508#
+ qr_4t1_mux_top_1/sky130_fd_sc_hs__dfxtp_2_7/a_1172_124# qr_4t1_mux_top_1/sky130_fd_sc_hs__dfxtp_4_1/a_1226_296#
+ qr_4t1_mux_top_1/sky130_fd_sc_hs__mux4_4_1/a_1465_377# qr_4t1_mux_top_1/sky130_fd_sc_hs__mux4_1_1/a_846_74#
+ qr_4t1_mux_top_1/sky130_fd_sc_hs__mux4_4_1/a_2199_74# qr_4t1_mux_top_1/sky130_fd_sc_hs__dfxtp_2_9/a_1217_314#
+ qr_4t1_mux_top_1/sky130_fd_sc_hs__dfxtp_4_3/a_206_368# qr_4t1_mux_top_1/sky130_fd_sc_hs__clkbuf_2_3/a_43_192#
+ qr_4t1_mux_top_1/sky130_fd_sc_hs__mux4_4_1/a_296_392# qr_4t1_mux_top_1/sky130_fd_sc_hs__dfxtp_2_1/a_1019_424#
+ qr_4t1_mux_top_1/sky130_fd_sc_hs__dfxtp_4_3/a_437_503# qr_4t1_mux_top_1/sky130_fd_sc_hs__dfxtp_2_11/a_431_508#
+ qr_4t1_mux_top_1/sky130_fd_sc_hs__dfxtp_2_5/a_1172_124# qr_4t1_mux_top_1/sky130_fd_sc_hs__dfxtp_2_9/a_27_74#
+ qr_4t1_mux_top_1/sky130_fd_sc_hs__dfxtp_2_7/a_1217_314# qr_4t1_mux_top_1/sky130_fd_sc_hs__dfxtp_2_9/a_206_368#
+ qr_4t1_mux_top_1/sky130_fd_sc_hs__dfxtp_2_3/a_1172_124# qr_4t1_mux_top_1/sky130_fd_sc_hs__dfxtp_2_5/a_695_459#
+ qr_4t1_mux_top_1/sky130_fd_sc_hs__mux4_4_1/a_2489_347# qr_4t1_mux_top_1/sky130_fd_sc_hs__mux4_1_1/a_763_341#
+ qr_4t1_mux_top_1/sky130_fd_sc_hs__dfxtp_4_3/a_1141_508# qr_4t1_mux_top_1/sky130_fd_sc_hs__mux4_4_1/a_299_126#
+ qr_4t1_mux_top_1/sky130_fd_sc_hs__dfxtp_2_9/a_708_101# qr_4t1_mux_top_1/sky130_fd_sc_hs__mux4_4_1/a_116_392#
+ qr_4t1_mux_top_1/sky130_fd_sc_hs__dfxtp_2_1/a_644_504# qr_4t1_mux_top_1/sky130_fd_sc_hs__mux4_1_1/a_979_74#
+ qr_4t1_mux_top_1/sky130_fd_sc_hs__dfxtp_2_5/a_1217_314# qr_4t1_mux_top_1/sky130_fd_sc_hs__dfxtp_4_1/a_735_102#
+ qr_4t1_mux_top_1/sky130_fd_sc_hs__clkbuf_1_5/a_27_74# qr_4t1_mux_top
Xsky130_fd_sc_hs__buf_1_0 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__buf_1_1/A sky130_fd_sc_hs__buf_1_1/X
+ sky130_fd_sc_hs__buf_1_1/a_27_164# sky130_fd_sc_hs__buf_1
Xsky130_fd_sc_hs__buf_2_109 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__buf_2_109/A sky130_fd_sc_hs__buf_2_109/X
+ sky130_fd_sc_hs__buf_2_109/a_21_260# sky130_fd_sc_hs__buf_2
Xsky130_fd_sc_hs__inv_4_16 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__inv_4_17/Y sky130_fd_sc_hs__inv_4_17/A
+ sky130_fd_sc_hs__inv_4
Xsky130_fd_sc_hs__inv_4_27 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__inv_4_27/Y osc_core_1/p1
+ sky130_fd_sc_hs__inv_4
Xsky130_fd_sc_hs__inv_4_38 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__inv_4_39/Y sky130_fd_sc_hs__inv_4_39/A
+ sky130_fd_sc_hs__inv_4
Xsky130_fd_sc_hs__inv_4_49 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__inv_4_49/Y osc_core_1/p3
+ sky130_fd_sc_hs__inv_4
Xsky130_fd_sc_hs__conb_1_160 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__conb_1_161/LO
+ sky130_fd_sc_hs__conb_1_161/HI sky130_fd_sc_hs__conb_1_161/a_165_290# sky130_fd_sc_hs__conb_1_161/a_21_290#
+ sky130_fd_sc_hs__conb_1
Xsky130_fd_sc_hs__conb_1_171 DVSS: DVDD: DVDD: DVSS: qr_4t1_mux_top_3/din_3_dummy
+ sky130_fd_sc_hs__conb_1_171/HI sky130_fd_sc_hs__conb_1_171/a_165_290# sky130_fd_sc_hs__conb_1_171/a_21_290#
+ sky130_fd_sc_hs__conb_1
Xsky130_fd_sc_hs__conb_1_182 DVSS: DVDD: DVDD: DVSS: prbs_generator_syn_23/eqn[8]
+ prbs_generator_syn_23/eqn[1] sky130_fd_sc_hs__conb_1_183/a_165_290# sky130_fd_sc_hs__conb_1_183/a_21_290#
+ sky130_fd_sc_hs__conb_1
Xsky130_fd_sc_hs__conb_1_193 DVSS: DVDD: DVDD: DVSS: prbs_generator_syn_19/eqn[13]
+ sky130_fd_sc_hs__conb_1_193/HI sky130_fd_sc_hs__conb_1_193/a_165_290# sky130_fd_sc_hs__conb_1_193/a_21_290#
+ sky130_fd_sc_hs__conb_1
Xsky130_fd_sc_hs__nand2_1_1 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__or2b_2_1/A sky130_fd_sc_hs__nor4_2_1/D
+ sky130_fd_sc_hs__nor2_4_1/Y sky130_fd_sc_hs__nand2_1_1/a_117_74# sky130_fd_sc_hs__nand2_1
Xsky130_fd_sc_hs__clkbuf_16_10 DVSS: DVDD: DVDD: DVSS: osc_core_1/pi1_l[3] sky130_fd_sc_hs__clkbuf_4_13/X
+ sky130_fd_sc_hs__clkbuf_16_11/a_114_74# sky130_fd_sc_hs__clkbuf_16
Xsky130_fd_sc_hs__clkbuf_16_21 DVSS: DVDD: DVDD: DVSS: osc_core_1/pi1_l[2] sky130_fd_sc_hs__clkbuf_4_21/X
+ sky130_fd_sc_hs__clkbuf_16_21/a_114_74# sky130_fd_sc_hs__clkbuf_16
Xsky130_fd_sc_hs__clkbuf_16_32 DVSS: DVDD: DVDD: DVSS: osc_core_1/pi3_l[0] sky130_fd_sc_hs__clkbuf_16_1/X
+ sky130_fd_sc_hs__clkbuf_16_33/a_114_74# sky130_fd_sc_hs__clkbuf_16
Xsky130_fd_sc_hs__clkbuf_16_43 DVSS: DVDD: DVDD: DVSS: test_mux_misc sky130_fd_sc_hs__inv_4_39/Y
+ sky130_fd_sc_hs__clkbuf_16_43/a_114_74# sky130_fd_sc_hs__clkbuf_16
Xsky130_fd_sc_hs__clkbuf_16_54 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__einvp_2_99/A
+ sky130_fd_sc_hs__einvp_2_65/A sky130_fd_sc_hs__clkbuf_16_55/a_114_74# sky130_fd_sc_hs__clkbuf_16
Xsky130_fd_sc_hs__clkbuf_16_65 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__nand2_2_3/B
+ sky130_fd_sc_hs__or2b_2_5/X sky130_fd_sc_hs__clkbuf_16_65/a_114_74# sky130_fd_sc_hs__clkbuf_16
Xsky130_fd_sc_hs__clkbuf_16_76 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__nor4_2_1/A
+ sky130_fd_sc_hs__clkbuf_8_79/X sky130_fd_sc_hs__clkbuf_16_77/a_114_74# sky130_fd_sc_hs__clkbuf_16
Xsky130_fd_sc_hs__clkbuf_16_87 DVSS: DVDD: DVDD: DVSS: hr_16t4_mux_top_1/clk sky130_fd_sc_hs__buf_1_1/X
+ sky130_fd_sc_hs__clkbuf_16_87/a_114_74# sky130_fd_sc_hs__clkbuf_16
Xsky130_fd_sc_hs__clkbuf_16_98 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__clkbuf_16_99/X
+ sky130_fd_sc_hs__clkbuf_4_123/X sky130_fd_sc_hs__clkbuf_16_99/a_114_74# sky130_fd_sc_hs__clkbuf_16
Xsky130_fd_sc_hs__clkbuf_16_120 DVSS: DVDD: DVDD: DVSS: prbs_generator_syn_31/clk
+ prbs_generator_syn_19/clk sky130_fd_sc_hs__clkbuf_16_121/a_114_74# sky130_fd_sc_hs__clkbuf_16
Xsky130_fd_sc_hs__clkbuf_16_131 DVSS: DVDD: DVDD: DVSS: osc_core_1/pi4_l[3] pi4_con[3]
+ sky130_fd_sc_hs__clkbuf_16_131/a_114_74# sky130_fd_sc_hs__clkbuf_16
Xsky130_fd_sc_hs__nand2_2_17 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__nand2_2_17/Y
+ sky130_fd_sc_hs__or2b_2_3/A sky130_fd_sc_hs__nand2_2_27/B sky130_fd_sc_hs__nand2_2_17/a_27_74#
+ sky130_fd_sc_hs__nand2_2
Xsky130_fd_sc_hs__nand2_2_28 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__nand2_2_29/Y
+ sky130_fd_sc_hs__nor2_4_1/B sky130_fd_sc_hs__nor2_4_1/A sky130_fd_sc_hs__nand2_2_29/a_27_74#
+ sky130_fd_sc_hs__nand2_2
Xprbs_generator_syn_6 prbs_generator_syn_9/clk prbs_generator_syn_9/rst prbs_generator_syn_7/cke
+ sky130_fd_sc_hs__conb_1_75/LO sky130_fd_sc_hs__conb_1_75/LO sky130_fd_sc_hs__conb_1_75/HI
+ sky130_fd_sc_hs__conb_1_75/HI sky130_fd_sc_hs__conb_1_75/HI sky130_fd_sc_hs__conb_1_75/LO
+ sky130_fd_sc_hs__conb_1_75/LO sky130_fd_sc_hs__conb_1_75/LO sky130_fd_sc_hs__conb_1_75/LO
+ sky130_fd_sc_hs__conb_1_75/LO sky130_fd_sc_hs__conb_1_75/LO sky130_fd_sc_hs__conb_1_73/LO
+ sky130_fd_sc_hs__conb_1_73/LO sky130_fd_sc_hs__conb_1_73/HI sky130_fd_sc_hs__conb_1_73/LO
+ sky130_fd_sc_hs__conb_1_73/LO sky130_fd_sc_hs__conb_1_73/LO sky130_fd_sc_hs__conb_1_73/LO
+ sky130_fd_sc_hs__conb_1_63/HI prbs_generator_syn_7/eqn[0] sky130_fd_sc_hs__conb_1_65/HI
+ sky130_fd_sc_hs__conb_1_65/LO sky130_fd_sc_hs__conb_1_65/HI sky130_fd_sc_hs__conb_1_65/HI
+ sky130_fd_sc_hs__conb_1_77/LO sky130_fd_sc_hs__conb_1_77/LO sky130_fd_sc_hs__conb_1_77/LO
+ sky130_fd_sc_hs__conb_1_79/LO sky130_fd_sc_hs__conb_1_79/LO sky130_fd_sc_hs__conb_1_79/LO
+ sky130_fd_sc_hs__conb_1_79/LO sky130_fd_sc_hs__conb_1_79/LO prbs_generator_syn_7/eqn[31]
+ prbs_generator_syn_7/eqn[31] prbs_generator_syn_7/eqn[31] prbs_generator_syn_7/eqn[28]
+ prbs_generator_syn_7/eqn[28] prbs_generator_syn_7/eqn[28] prbs_generator_syn_7/eqn[28]
+ prbs_generator_syn_7/eqn[28] prbs_generator_syn_7/eqn[28] prbs_generator_syn_7/eqn[28]
+ prbs_generator_syn_7/eqn[21] prbs_generator_syn_7/eqn[20] prbs_generator_syn_7/eqn[21]
+ prbs_generator_syn_7/eqn[21] prbs_generator_syn_7/eqn[21] prbs_generator_syn_7/eqn[21]
+ prbs_generator_syn_7/eqn[21] prbs_generator_syn_7/eqn[21] prbs_generator_syn_7/eqn[21]
+ prbs_generator_syn_7/eqn[9] prbs_generator_syn_7/eqn[9] prbs_generator_syn_7/eqn[9]
+ prbs_generator_syn_7/eqn[9] prbs_generator_syn_7/eqn[8] prbs_generator_syn_7/eqn[8]
+ prbs_generator_syn_7/eqn[8] prbs_generator_syn_7/eqn[8] prbs_generator_syn_7/eqn[8]
+ prbs_generator_syn_7/eqn[8] prbs_generator_syn_7/eqn[8] prbs_generator_syn_7/eqn[1]
+ prbs_generator_syn_7/eqn[0] prbs_generator_syn_9/inj_err sky130_fd_sc_hs__conb_1_73/LO
+ sky130_fd_sc_hs__conb_1_73/LO prbs_generator_syn_7/out DVSS: DVDD: prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_1/a_293_74#
+ prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_15/X prbs_generator_syn_7/sky130_fd_sc_hs__nand2_1_35/B
+ prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_51/Y prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_9/A
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_9/CLK prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_47/a_27_74#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_37/a_1226_296# prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_3/B
+ prbs_generator_syn_7/sky130_fd_sc_hs__nor2b_1_7/a_27_112# prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_29/B
+ prbs_generator_syn_7/sky130_fd_sc_hs__sdlclkp_2_1/a_580_74# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_1/a_1141_508#
+ prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_5/Y prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_41/a_230_79#
+ prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_61/a_138_385# prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_43/a_132_392#
+ prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_3/a_222_392# prbs_generator_syn_7/sky130_fd_sc_hs__nor2b_1_9/a_27_112#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_61/a_27_74# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_35/a_206_368#
+ prbs_generator_syn_7/sky130_fd_sc_hs__nand2_2_3/Y prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_25/B
+ prbs_generator_syn_7/sky130_fd_sc_hs__nand2_1_11/a_117_74# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_67/a_651_503#
+ prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_45/X prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_39/a_696_458#
+ prbs_generator_syn_7/sky130_fd_sc_hs__sdlclkp_2_1/a_1198_74# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_45/a_1034_424#
+ prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_17/a_222_392# prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_55/a_222_392#
+ prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_53/Y prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_35/A
+ prbs_generator_syn_7/m3_13600_1651# prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_59/a_52_123#
+ prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_5/a_293_74# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_35/a_1226_296#
+ prbs_generator_syn_7/sky130_fd_sc_hs__nand2_1_51/B prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_5/a_651_503#
+ prbs_generator_syn_7/sky130_fd_sc_hs__nand2_1_21/B prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_8/a_27_74#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_15/a_27_74# prbs_generator_syn_7/sky130_fd_sc_hs__and2b_2_1/X
+ prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_13/X prbs_generator_syn_7/sky130_fd_sc_hs__nand2_2_3/a_27_74#
+ prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_50/a_138_385# prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_33/a_132_392#
+ prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_1/a_376_368# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_25/a_206_368#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_35/a_437_503# prbs_generator_syn_7/sky130_fd_sc_hs__sdlclkp_2_1/a_708_451#
+ prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_45/a_230_79# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_29/a_696_458#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_32/a_27_74# prbs_generator_syn_7/sky130_fd_sc_hs__nor2b_1_4/Y
+ prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_59/a_293_74# prbs_generator_syn_7/sky130_fd_sc_hs__nand2_1_47/a_117_74#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_73/a_735_102# prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_21/a_112_119#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_23/a_1141_508# prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_25/a_293_74#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_7/Q prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_3/a_112_119#
+ prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_35/B prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_51/X
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_53/a_1178_124# prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_23/a_132_392#
+ prbs_generator_syn_7/sky130_fd_sc_hs__nand2_1_3/B prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_15/a_206_368#
+ prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_63/a_132_392# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_55/a_27_74#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_25/a_437_503# prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_41/a_52_123#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_47/a_651_503# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_73/a_1141_508#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_19/a_696_458# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_57/a_696_458#
+ prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_7/X prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_43/a_1034_424#
+ prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_55/A prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_11/a_112_119#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_21/a_1141_508# prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_35/a_222_392#
+ prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_49/a_230_79# prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_67/Y
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_71/a_27_74# prbs_generator_syn_7/sky130_fd_sc_hs__nand2_1_33/B
+ prbs_generator_syn_7/sky130_fd_sc_hs__conb_1_1/LO prbs_generator_syn_7/sky130_fd_sc_hs__nand2_1_19/a_117_74#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_51/a_1178_124# prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_33/X
+ prbs_generator_syn_7/sky130_fd_sc_hs__nand2_1_29/B prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_41/Y
+ prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_53/a_132_392# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_45/a_206_368#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_15/a_437_503# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_37/a_651_503#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_39/a_544_485# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_53/a_735_102#
+ prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_45/a_52_123# prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_1/B
+ prbs_generator_syn_7/sky130_fd_sc_hs__nand2_2_3/B prbs_generator_syn_7/sky130_fd_sc_hs__clkbuf_16_1/A
+ prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_21/X prbs_generator_syn_7/sky130_fd_sc_hs__nand2_1_25/B
+ prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_39/a_376_368# prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_63/X
+ prbs_generator_syn_7/m3_13600_3481# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_69/a_1178_124#
+ prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_21/a_138_385# prbs_generator_syn_7/sky130_fd_sc_hs__nor2b_1_8/Y
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_19/a_1178_124# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_49/a_27_74#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_45/a_437_503# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_27/a_651_503#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_71/a_1141_508# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_65/a_651_503#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_29/a_544_485# prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_3/a_138_385#
+ prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_55/X prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_43/a_735_102#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_41/a_1034_424# prbs_generator_syn_7/sky130_fd_sc_hs__nand2_1_9/B
+ prbs_generator_syn_7/sky130_fd_sc_hs__nor2b_1_9/Y prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_59/a_1034_424#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_39/a_1141_508# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_33/a_1226_296#
+ prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_49/a_52_123# prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_47/Y
+ prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_43/Y prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_4/a_651_503#
+ prbs_generator_syn_7/sky130_fd_sc_hs__nand2_1_49/B prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_19/A
+ prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_11/a_138_385# prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_5/X
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_63/a_206_368# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_17/a_651_503#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_19/a_544_485# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_55/a_651_503#
+ prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_9/Y prbs_generator_syn_7/sky130_fd_sc_hs__nand2_1_17/B
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_57/a_544_485# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_67/a_696_458#
+ prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_35/X prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_19/a_27_74#
+ prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_45/a_222_392# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_32/a_1226_296#
+ prbs_generator_syn_7/sky130_fd_sc_hs__nand2_1_43/B prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_25/A
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_1/a_206_368# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_49/a_1226_296#
+ prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_1/a_112_119# prbs_generator_syn_7/sky130_fd_sc_hs__or2_1_1/X
+ prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_59/a_376_368# prbs_generator_syn_7/sky130_fd_sc_hs__nand2_1_19/B
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_5/a_696_458# prbs_generator_syn_7/sky130_fd_sc_hs__nor2b_1_1/Y
+ prbs_generator_syn_7/sky130_fd_sc_hs__nor2b_1_5/a_278_368# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_17/a_1178_124#
+ prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_39/X prbs_generator_syn_7/m3_13600_5433#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_63/a_437_503# prbs_generator_syn_7/sky130_fd_sc_hs__nand2_2_5/B
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_23/a_735_102# prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_53/A
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_61/a_735_102# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_57/a_1034_424#
+ prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_63/B prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_37/a_1141_508#
+ prbs_generator_syn_7/sky130_fd_sc_hs__nand2_1_47/B prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_29/X
+ prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_65/Y prbs_generator_syn_7/m3_13600_4701#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_1/a_437_503# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_67/a_1178_124#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_9/a_735_102# prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_13/a_132_392#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_15/a_1178_124# prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_15/A
+ prbs_generator_syn_7/sky130_fd_sc_hs__nand2_1_1/B prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_43/B
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_35/a_651_503# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_8/D
+ prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_29/A prbs_generator_syn_7/sky130_fd_sc_hs__nand2_1_7/B
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_13/a_735_102# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_47/a_696_458#
+ prbs_generator_syn_7/sky130_fd_sc_hs__nand2_1_31/B prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_51/a_735_102#
+ prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_59/X prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_35/a_1141_508#
+ prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_25/a_222_392# prbs_generator_syn_7/sky130_fd_sc_hs__sdlclkp_2_1/a_288_48#
+ prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_55/B prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_17/B
+ prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_43/A prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_7/A
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_65/a_1178_124# prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_59/Y
+ prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_41/X prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_21/a_230_79#
+ prbs_generator_syn_7/sky130_fd_sc_hs__nand2_1_57/a_117_74# prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_1/a_222_392#
+ prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_19/B prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_35/a_293_74#
+ prbs_generator_syn_7/sky130_fd_sc_hs__nand2_1_23/a_117_74# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_73/a_206_368#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_25/a_651_503# prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_1/a_138_385#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_37/a_696_458# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_67/a_544_485#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_43/a_27_74# prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_9/X
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_55/a_1034_424# prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_39/a_112_119#
+ prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_15/a_222_392# prbs_generator_syn_7/sky130_fd_sc_hs__conb_1_1/HI
+ prbs_generator_syn_7/sky130_fd_sc_hs__nand2_1_23/B prbs_generator_syn_7/sky130_fd_sc_hs__nand2_1_53/B
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_9/a_1178_124# prbs_generator_syn_7/sky130_fd_sc_hs__nor2b_1_4/A
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_47/a_1226_296# prbs_generator_syn_7/m3_13600_11045#
+ prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_17/X prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_29/a_376_368#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_5/a_544_485# prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_3/X
+ prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_31/a_132_392# prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_61/A
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_15/a_651_503# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_73/a_437_503#
+ prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_25/a_230_79# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_27/a_696_458#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_65/a_696_458# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_33/a_735_102#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_71/a_735_102# prbs_generator_syn_7/m3_13600_7263#
+ prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_43/a_222_392# prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_50/Y
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_8/a_1178_124# prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_53/B
+ prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_19/a_376_368# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_63/a_1178_124#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_4/a_696_458# prbs_generator_syn_7/sky130_fd_sc_hs__nor2b_1_4/a_278_368#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_13/a_1178_124# prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_61/a_132_392#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_53/a_206_368# prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_21/a_52_123#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_45/a_651_503# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_17/a_696_458#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_47/a_544_485# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_55/a_696_458#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_21/a_735_102# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_37/a_27_74#
+ prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_61/B prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_61/X
+ prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_59/a_112_119# prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_31/A
+ prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_33/a_222_392# prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_29/a_230_79#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_45/a_1226_296# prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_9/a_132_392#
+ prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_5/A prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_57/Y
+ prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_31/X prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_51/a_27_74#
+ prbs_generator_syn_7/sky130_fd_sc_hs__nor2b_1_8/a_27_112# prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_47/a_376_368#
+ prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_53/a_293_74# prbs_generator_syn_7/sky130_fd_sc_hs__nand2_1_43/a_117_74#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_8/a_735_102# prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_21/a_293_74#
+ prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_39/a_138_385# prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_63/Y
+ prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_51/a_132_392# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_43/a_206_368#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_53/a_437_503# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_37/a_544_485#
+ prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_57/X prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_53/a_1034_424#
+ prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_25/a_52_123# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_33/a_1141_508#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_63/Q prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_23/a_222_392#
+ prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_63/a_222_392# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_7/a_1178_124#
+ prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_53/X prbs_generator_syn_7/sky130_fd_sc_hs__nand2_2_5/Y
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_61/a_1178_124# prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_1/a_230_79#
+ prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_43/a_230_79# prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_11/a_230_79#
+ prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_41/a_132_392# prbs_generator_syn_7/sky130_fd_sc_hs__nand2_1_13/a_117_74#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_43/a_437_503# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_27/a_544_485#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_63/a_651_503# prbs_generator_syn_7/sky130_fd_sc_hs__nand2_1_7/a_117_74#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_35/a_696_458# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_65/a_544_485#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_51/a_1034_424# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_41/a_735_102#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_32/a_1141_508# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_49/a_1141_508#
+ prbs_generator_syn_7/sky130_fd_sc_hs__nand2_1_55/B prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_53/a_222_392#
+ prbs_generator_syn_7/sky130_fd_sc_hs__sdlclkp_2_1/a_114_112# prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_9/a_293_74#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_43/a_1226_296# prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_29/a_52_123#
+ prbs_generator_syn_7/sky130_fd_sc_hs__nand2_1_37/B prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_1/a_651_503#
+ prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_27/a_376_368# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_4/a_544_485#
+ prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_67/a_376_368# prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_27/X
+ prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_1/X prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_59/a_138_385#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_29/a_1178_124# prbs_generator_syn_7/m3_13600_2871#
+ prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_5/a_230_79# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_23/a_206_368#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_61/a_206_368# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_17/a_544_485#
+ prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_15/a_230_79# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_25/a_696_458#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_55/a_544_485# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_32/a_735_102#
+ prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_29/a_293_74# prbs_generator_syn_7/sky130_fd_sc_hs__nand2_1_17/a_117_74#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_69/a_1034_424# prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_29/a_112_119#
+ prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_37/X prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_31/B
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_19/a_1034_424# prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_33/A
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_9/a_206_368# prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_57/a_376_368#
+ prbs_generator_syn_7/sky130_fd_sc_hs__sdlclkp_2_1/a_706_317# prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_11/B
+ prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_1/a_52_123# prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_39/B
+ prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_21/a_132_392# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_13/a_206_368#
+ prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_43/a_52_123# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_51/a_206_368#
+ prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_47/X prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_23/a_437_503#
+ prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_11/a_52_123# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_61/a_437_503#
+ prbs_generator_syn_7/sky130_fd_sc_hs__nor2b_1_7/Y prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_51/A
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_15/a_696_458# prbs_generator_syn_7/sky130_fd_sc_hs__nor2b_1_5/Y
+ prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_9/a_230_79# prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_25/X
+ prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_19/a_112_119# prbs_generator_syn_7/sky130_fd_sc_hs__nand2_1_45/B
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_5/a_1178_124# prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_19/a_230_79#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_41/a_1226_296# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_59/a_1226_296#
+ prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_63/a_230_79# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_51/Q
+ prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_7/a_132_392# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_9/a_437_503#
+ prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_46/a_376_368# prbs_generator_syn_7/sky130_fd_sc_hs__nand2_1_33/a_117_74#
+ prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_11/a_293_74# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_27/a_1178_124#
+ prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_11/a_132_392# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_13/a_437_503#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_51/a_437_503# prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_5/a_52_123#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_35/a_544_485# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_73/a_651_503#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_45/a_696_458# prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_15/a_52_123#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_47/a_1141_508# prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_47/a_112_119#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_4/a_1178_124# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_17/a_1034_424#
+ prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_23/B prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_37/a_376_368#
+ prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_15/B prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_7/Y
+ prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_29/a_138_385# prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_33/a_230_79#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_25/a_1178_124# prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_47/a_293_74#
+ prbs_generator_syn_7/sky130_fd_sc_hs__nand2_1_37/a_117_74# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_33/a_206_368#
+ prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_15/a_293_74# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_71/a_206_368#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_25/a_544_485# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_67/a_1034_424#
+ prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_13/a_222_392# prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_9/a_52_123#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_15/a_1034_424# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_57/a_1226_296#
+ prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_19/a_52_123# prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_23/X
+ prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_63/a_52_123# prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_19/a_138_385#
+ prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_9/a_376_368# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_21/a_206_368#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_33/a_437_503# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_71/a_437_503#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_53/a_651_503# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_15/a_544_485#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_63/a_696_458# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_65/a_1034_424#
+ prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_19/a_293_74# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_45/a_1141_508#
+ prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_27/a_112_119# prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_67/a_112_119#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_1/a_1178_124# prbs_generator_syn_7/sky130_fd_sc_hs__conb_1_1/a_21_290#
+ prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_63/a_293_74# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_8/a_206_368#
+ prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_17/a_376_368# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_63/a_27_74#
+ prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_21/A prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_55/a_376_368#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_1/a_696_458# prbs_generator_syn_7/sky130_fd_sc_hs__nor2b_1_1/a_278_368#
+ prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_47/a_138_385# prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_33/a_52_123#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_9/a_1034_424# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_21/a_437_503#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_1/a_27_74# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_43/a_651_503#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_1/Q prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_45/a_544_485#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_69/a_735_102# prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_57/a_112_119#
+ prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_31/a_222_392# prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_13/A
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_55/a_1226_296# prbs_generator_syn_7/sky130_fd_sc_hs__nand2_2_5/a_27_74#
+ prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_53/a_230_79# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_8/a_437_503#
+ prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_67/a_293_74# prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_33/a_293_74#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_7/a_735_102# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_23/a_1178_124#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_41/a_206_368# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_8/a_1034_424#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_63/a_1034_424# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_59/a_735_102#
+ prbs_generator_syn_7/sky130_fd_sc_hs__nand2_1_5/B prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_43/a_1141_508#
+ prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_46/a_112_119# prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_61/a_222_392#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_13/a_1034_424# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_73/a_1178_124#
+ prbs_generator_syn_7/sky130_fd_sc_hs__nand2_1_27/B prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_13/B
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_57/a_27_74# prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_57/a_230_79#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_21/a_1178_124# prbs_generator_syn_7/sky130_fd_sc_hs__nor2b_1_1/a_27_112#
+ prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_27/a_138_385# prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_23/a_230_79#
+ prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_67/a_138_385# prbs_generator_syn_7/sky130_fd_sc_hs__nand2_1_41/B
+ prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_9/a_222_392# prbs_generator_syn_7/sky130_fd_sc_hs__nand2_1_27/a_117_74#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_32/a_206_368# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_23/a_651_503#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_41/a_437_503# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_73/a_27_74#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_61/a_651_503# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_63/a_544_485#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_49/a_735_102# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_73/a_696_458#
+ prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_37/a_112_119# prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_51/a_222_392#
+ prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_43/X prbs_generator_syn_7/sky130_fd_sc_hs__nand2_2_1/B
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_9/a_651_503# prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_53/a_52_123#
+ prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_49/X prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_25/a_376_368#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_1/a_544_485# prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_65/a_376_368#
+ prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_57/a_138_385# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_27/a_27_74#
+ prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_39/a_132_392# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_7/a_1034_424#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_13/a_651_503# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_32/a_437_503#
+ prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_27/a_230_79# prbs_generator_syn_7/m3_13600_12265#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_51/a_651_503# prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_59/B
+ prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_47/A prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_61/a_1034_424#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_41/a_1141_508# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_59/a_1141_508#
+ prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_41/a_222_392# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_53/a_1226_296#
+ prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_3/A prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_71/a_1178_124#
+ prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_9/a_112_119# prbs_generator_syn_7/sky130_fd_sc_hs__nand2_1_3/a_117_74#
+ prbs_generator_syn_7/m3_13600_8483# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_39/a_1178_124#
+ prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_57/a_52_123# prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_46/a_138_385#
+ prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_23/a_52_123# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_67/a_27_74#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_53/a_696_458# prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_17/a_112_119#
+ prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_11/A prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_55/a_112_119#
+ prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_1/A prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_51/a_1226_296#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_29/a_1034_424# prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_59/A
+ prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_23/A prbs_generator_syn_7/sky130_fd_sc_hs__nand2_1_39/B
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_5/a_27_74# prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_57/a_293_74#
+ prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_37/a_138_385# prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_59/a_132_392#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_33/a_651_503# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_71/a_651_503#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_43/a_696_458# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_73/a_544_485#
+ prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_27/a_52_123# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_57/a_1141_508#
+ prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_21/a_222_392# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_35/a_27_74#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_69/a_1226_296# prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_37/B
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_19/a_1226_296# prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_35/a_376_368#
+ prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_47/a_230_79# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_37/a_1178_124#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_5/a_1034_424# prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_49/a_132_392#
+ prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_7/a_222_392# prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_27/a_293_74#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_21/a_651_503# prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_9/a_138_385#
+ prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_11/a_222_392# prbs_generator_syn_7/m3_13600_14095#
+ prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_50/A prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_27/a_1034_424#
+ prbs_generator_syn_7/sky130_fd_sc_hs__nand2_1_13/B prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_8/a_651_503#
+ prbs_generator_syn_7/m3_13600_9703# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_35/a_1178_124#
+ prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_17/a_138_385# prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_55/a_138_385#
+ prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_7/a_230_79# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_4/a_1034_424#
+ prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_7/a_376_368# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_69/a_206_368#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_23/a_696_458# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_53/a_544_485#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_39/a_735_102# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_61/a_696_458#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_55/a_1141_508# prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_25/a_112_119#
+ prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_65/a_112_119# prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_43/a_293_74#
+ prbs_generator_syn_7/sky130_fd_sc_hs__nand2_1_57/B prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_25/a_1034_424#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_7/a_206_368# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_17/a_1226_296#
+ prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_15/a_376_368# prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_53/a_376_368#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_9/a_696_458# prbs_generator_syn_7/m3_13600_431#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_45/a_27_74# prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_47/a_52_123#
+ prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_29/a_132_392# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_59/a_206_368#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_69/a_437_503# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_41/a_651_503#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_43/a_544_485# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_13/a_696_458#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_29/a_735_102# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_51/a_696_458#
+ prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_61/Y prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_67/a_1226_296#
+ prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_5/a_132_392# prbs_generator_syn_7/sky130_fd_sc_hs__and2b_2_1/a_198_48#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_7/a_437_503# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_15/a_1226_296#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_69/a_27_74# prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_46/a_293_74#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_1/a_1034_424# prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_19/a_132_392#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_49/a_206_368# prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_7/a_52_123#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_59/a_437_503# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_32/a_651_503#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_7/a_27_74# prbs_generator_syn_7/sky130_fd_sc_hs__nand2_2_1/a_27_74#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_19/a_735_102# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_57/a_735_102#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_65/a_1226_296# prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_37/A
+ prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_33/a_376_368# prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_37/a_230_79#
+ prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_25/a_138_385# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_39/a_27_74#
+ prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_65/a_138_385# prbs_generator_syn_7/sky130_fd_sc_hs__nor2b_1_9/a_278_368#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_49/a_437_503# prbs_generator_syn_7/sky130_fd_sc_hs__and2b_2_1/a_505_74#
+ prbs_generator_syn_7/sky130_fd_sc_hs__nand2_1_51/a_117_74# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_23/a_544_485#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_33/a_696_458# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_61/a_544_485#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_9/a_1226_296# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_53/a_1141_508#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_71/a_696_458# prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_35/a_112_119#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_23/a_1034_424# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_9/a_544_485#
+ prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_63/a_376_368# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_33/a_1178_124#
+ prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_5/a_376_368# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_13/a_544_485#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_73/a_1034_424# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_21/a_696_458#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_51/a_544_485# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_8/a_1226_296#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_51/a_1141_508# prbs_generator_syn_7/sky130_fd_sc_hs__nand2_1_55/a_117_74#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_21/a_1034_424# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_63/a_1226_296#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_23/a_27_74# prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_7/a_112_119#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_13/a_1226_296# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_8/a_696_458#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_32/a_1178_124# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_49/a_1178_124#
+ prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_37/a_52_123# prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_27/a_132_392#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_71/Q prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_67/a_735_102#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_69/a_1141_508# prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_15/a_112_119#
+ prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_53/a_112_119# prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_39/a_222_392#
+ prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_55/a_230_79# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_19/a_1141_508#
+ prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_37/a_293_74# prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_43/a_376_368#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_5/a_735_102# prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_35/a_138_385#
+ prbs_generator_syn_7/sky130_fd_sc_hs__sdlclkp_2_1/a_114_424# prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_57/a_132_392#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_71/a_1034_424# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_7/a_1226_296#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_33/a_544_485# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_41/a_696_458#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_71/a_544_485# prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_21/B
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_61/a_1226_296# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_39/a_1034_424#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_17/a_27_74# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_9/a_27_74#
+ prbs_generator_syn_7/sky130_fd_sc_hs__nor2b_1_5/a_27_112# prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_47/a_132_392#
+ prbs_generator_syn_7/sky130_fd_sc_hs__nor2b_1_8/a_278_368# prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_9/B
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_39/a_206_368# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_33/a_27_74#
+ prbs_generator_syn_7/sky130_fd_sc_hs__nand2_1_41/a_117_74# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_69/a_651_503#
+ prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_51/a_293_74# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_21/a_544_485#
+ prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_7/a_138_385# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_32/a_696_458#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_47/a_735_102# prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_33/a_112_119#
+ prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_59/a_222_392# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_17/a_1141_508#
+ prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_55/a_52_123# prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_3/a_293_74#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_7/a_651_503# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_29/a_1226_296#
+ prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_23/a_376_368# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_8/a_544_485#
+ prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_47/B prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_47/a_1178_124#
+ prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_15/a_138_385# prbs_generator_syn_7/sky130_fd_sc_hs__sdlclkp_2_1/a_1195_374#
+ prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_53/a_138_385# prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_37/a_132_392#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_29/a_206_368# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_39/a_437_503#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_59/a_651_503# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_37/a_735_102#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_67/a_1141_508# prbs_generator_syn_7/sky130_fd_sc_hs__and2b_2_1/a_27_74#
+ prbs_generator_syn_7/sky130_fd_sc_hs__conb_1_1/a_165_290# prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_55/a_293_74#
+ prbs_generator_syn_7/sky130_fd_sc_hs__nand2_1_45/a_117_74# prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_63/a_112_119#
+ prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_49/a_222_392# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_37/a_1034_424#
+ prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_23/a_293_74# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_15/a_1141_508#
+ prbs_generator_syn_7/sky130_fd_sc_hs__nand2_1_5/a_117_74# prbs_generator_syn_7/m3_13600_13485#
+ prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_5/a_112_119# prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_13/a_376_368#
+ prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_51/a_376_368# prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_7/a_293_74#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_19/a_206_368# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_57/a_206_368#
+ prbs_generator_syn_7/sky130_fd_sc_hs__sdlclkp_2_1/a_318_74# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_29/a_437_503#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_49/a_651_503# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_25/a_27_74#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_5/a_1226_296# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_41/a_544_485#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_27/a_735_102# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_65/a_1141_508#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_65/a_735_102# prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_3/a_230_79#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_35/a_1034_424# prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_13/a_230_79#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_41/a_27_74# prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_3/a_132_392#
+ prbs_generator_syn_7/sky130_fd_sc_hs__nand2_1_49/a_117_74# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_27/a_1226_296#
+ prbs_generator_syn_7/sky130_fd_sc_hs__nand2_1_15/a_117_74# prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_41/a_376_368#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_45/a_1178_124# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_4/a_735_102#
+ prbs_generator_syn_7/sky130_fd_sc_hs__nand2_1_9/a_117_74# prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_33/a_138_385#
+ prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_17/a_132_392# prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_55/a_132_392#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_9/a_1141_508# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_19/a_437_503#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_57/a_437_503# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_4/a_1226_296#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_32/a_544_485# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_17/a_735_102#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_55/a_735_102# prbs_generator_syn_7/m3_13600_2261#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_65/a_27_74# prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_29/a_222_392#
+ prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_43/a_112_119# prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_19/X
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_25/a_1226_296# prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_31/a_376_368#
+ prbs_generator_syn_7/sky130_fd_sc_hs__or2_1_1/a_63_368# prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_17/a_230_79#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_4/a_27_74# prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_61/a_230_79#
+ prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_63/a_138_385# prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_5/a_222_392#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_8/a_1141_508# prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_41/a_293_74#
+ prbs_generator_syn_7/sky130_fd_sc_hs__nand2_1_31/a_117_74# prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_5/a_138_385#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_63/a_1141_508# prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_19/a_222_392#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_13/a_1141_508# prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_3/a_52_123#
+ prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_13/a_52_123# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_43/a_1178_124#
+ prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_61/a_376_368# prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_35/a_132_392#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_67/a_206_368# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_1/a_1226_296#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_69/a_696_458# prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_31/a_230_79#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_35/a_735_102# prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_23/a_112_119#
+ prbs_generator_syn_7/sky130_fd_sc_hs__nand2_1_35/a_117_74# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_59/a_27_74#
+ prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_13/a_293_74# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_5/a_206_368#
+ prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_50/a_376_368# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_7/a_696_458#
+ prbs_generator_syn_7/sky130_fd_sc_hs__nor2b_1_7/a_278_368# prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_17/a_52_123#
+ prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_43/a_138_385# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_7/a_1141_508#
+ prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_61/a_52_123# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_67/a_437_503#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_61/a_1141_508# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_25/a_735_102#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_59/a_696_458# prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_13/a_112_119#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_33/a_1034_424# prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_51/a_112_119#
+ prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_35/a_230_79# prbs_generator_syn_7/m3_13600_4091#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_23/a_1226_296# prbs_generator_syn_7/sky130_fd_sc_hs__nand2_1_39/a_117_74#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_29/a_27_74# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_5/a_437_503#
+ prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_17/a_293_74# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_41/a_1178_124#
+ prbs_generator_syn_7/sky130_fd_sc_hs__or2_1_1/a_152_368# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_59/a_1178_124#
+ prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_61/a_293_74# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_47/a_206_368#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_39/a_651_503# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_49/a_696_458#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_15/a_735_102# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_32/a_1034_424#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_73/a_1226_296# prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_27/a_222_392#
+ prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_41/a_112_119# prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_31/a_52_123#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_49/a_1034_424# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_29/a_1141_508#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_21/a_1226_296# prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_39/a_230_79#
+ prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_23/a_138_385# prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_51/a_230_79#
+ prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_45/a_132_392# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_37/a_206_368#
+ prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_65/a_293_74# prbs_generator_syn_7/sky130_fd_sc_hs__nand2_1_53/a_117_74#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_47/a_437_503# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_29/a_651_503#
+ prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_31/a_293_74# prbs_generator_syn_7/sky130_fd_sc_hs__nand2_1_21/a_117_74#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_69/a_544_485# prbs_generator_syn_7/sky130_fd_sc_hs__clkbuf_16_1/a_114_74#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_45/a_735_102# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_13/a_27_74#
+ prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_31/a_112_119# prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_57/a_222_392#
+ prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_35/a_52_123# prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_21/a_376_368#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_7/a_544_485# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_57/a_1178_124#
+ prbs_generator_syn_7/m3_13600_6043# prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_13/a_138_385#
+ prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_51/a_138_385# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_5/a_1141_508#
+ prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_3/a_376_368# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_27/a_206_368#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_65/a_206_368# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_37/a_437_503#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_19/a_651_503# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_57/a_651_503#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_59/a_544_485# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_71/a_1226_296#
+ prbs_generator_syn_7/sky130_fd_sc_hs__nand2_1_25/a_117_74# prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_61/a_112_119#
+ prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_47/a_222_392# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_27/a_1141_508#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_53/a_27_74# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_4/a_206_368#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_39/a_1226_296# prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_11/a_376_368#
+ prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_39/a_52_123# prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_41/a_138_385#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_4/a_1141_508# prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_25/a_132_392#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_17/a_206_368# prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_41/A
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_55/a_206_368# prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_51/a_52_123#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_27/a_437_503# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_65/a_437_503#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_49/a_544_485# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_63/a_735_102#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_47/a_1034_424# prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_50/a_112_119#
+ prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_37/a_222_392# prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_59/a_230_79#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_25/a_1141_508# prbs_generator_syn_7/sky130_fd_sc_hs__nor2b_1_4/a_27_112#
+ prbs_generator_syn_7/sky130_fd_sc_hs__sdlclkp_2_1/a_685_81# prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_1/a_132_392#
+ prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_39/a_293_74# prbs_generator_syn_7/sky130_fd_sc_hs__nand2_1_29/a_117_74#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_4/a_437_503# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_55/a_1178_124#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_21/a_27_74# prbs_generator_syn_7/m3_13600_12875#
+ prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_50/a_293_74# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_1/a_735_102#
+ prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_31/a_138_385# prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_15/a_132_392#
+ prbs_generator_syn_7/sky130_fd_sc_hs__nand2_1_1/a_117_74# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_17/a_437_503#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_55/a_437_503# prbs_generator_syn
Xsky130_fd_sc_hs__clkbuf_4_120 DVSS: DVDD: DVDD: DVSS: CTL_BUF_P[0] sky130_fd_sc_hs__clkbuf_8_79/A
+ sky130_fd_sc_hs__clkbuf_4_121/a_83_270# sky130_fd_sc_hs__clkbuf_4
Xsky130_fd_sc_hs__clkbuf_4_131 DVSS: DVDD: DVDD: DVSS: pi5_con[2] sky130_fd_sc_hs__clkbuf_4_131/X
+ sky130_fd_sc_hs__clkbuf_4_131/a_83_270# sky130_fd_sc_hs__clkbuf_4
Xsky130_fd_sc_hs__o21ai_2_0 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__inv_4_11/Y sky130_fd_sc_hs__o21ai_2_3/A2
+ sky130_fd_sc_hs__nand2_2_3/B sky130_fd_sc_hs__buf_2_39/A sky130_fd_sc_hs__o21ai_2_1/a_116_368#
+ sky130_fd_sc_hs__o21ai_2_1/a_27_74# sky130_fd_sc_hs__o21ai_2
Xsky130_fd_sc_hs__clkdlyinv5sd2_1_5 DVSS: DVDD: DVSS: DVDD: dout_n sky130_fd_sc_hs__and2_2_1/B
+ sky130_fd_sc_hs__clkdlyinv5sd2_1_5/a_28_74# sky130_fd_sc_hs__clkdlyinv5sd2_1_5/a_682_74#
+ sky130_fd_sc_hs__clkdlyinv5sd2_1_5/a_549_74# sky130_fd_sc_hs__clkdlyinv5sd2_1_5/a_288_74#
+ sky130_fd_sc_hs__clkdlyinv5sd2_1
Xsky130_fd_sc_hs__clkbuf_4_60 DVSS: DVDD: DVDD: DVSS: fine_control_avg_window_select[3]
+ sky130_fd_sc_hs__clkbuf_4_61/X sky130_fd_sc_hs__clkbuf_4_61/a_83_270# sky130_fd_sc_hs__clkbuf_4
Xsky130_fd_sc_hs__clkbuf_4_71 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__nand2_2_5/Y
+ sky130_fd_sc_hs__inv_4_11/A sky130_fd_sc_hs__clkbuf_4_71/a_83_270# sky130_fd_sc_hs__clkbuf_4
Xsky130_fd_sc_hs__clkbuf_4_82 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__nand2_2_15/Y
+ sky130_fd_sc_hs__dlrtp_1_24/D sky130_fd_sc_hs__clkbuf_4_83/a_83_270# sky130_fd_sc_hs__clkbuf_4
Xsky130_fd_sc_hs__clkbuf_4_93 DVSS: DVDD: DVDD: DVSS: div_ratio_half[3] sky130_fd_sc_hs__clkbuf_4_93/X
+ sky130_fd_sc_hs__clkbuf_4_93/a_83_270# sky130_fd_sc_hs__clkbuf_4
Xsky130_fd_sc_hs__o21ai_2_18 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__inv_4_17/Y sky130_fd_sc_hs__o21ai_2_23/A2
+ sky130_fd_sc_hs__nand2_2_7/A sky130_fd_sc_hs__o21ai_2_19/Y sky130_fd_sc_hs__o21ai_2_19/a_116_368#
+ sky130_fd_sc_hs__o21ai_2_19/a_27_74# sky130_fd_sc_hs__o21ai_2
Xsky130_fd_sc_hs__o21ai_2_29 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__inv_4_21/Y sky130_fd_sc_hs__or2b_4_1/A
+ sky130_fd_sc_hs__buf_8_3/X sky130_fd_sc_hs__buf_2_95/A sky130_fd_sc_hs__o21ai_2_29/a_116_368#
+ sky130_fd_sc_hs__o21ai_2_29/a_27_74# sky130_fd_sc_hs__o21ai_2
Xqr_4t1_mux_top_1 qr_4t1_mux_top_1/clk_Q hr_16t4_mux_top_1/clk qr_4t1_mux_top_3/clk_I
+ qr_4t1_mux_top_1/clk_IB qr_4t1_mux_top_1/din[3] qr_4t1_mux_top_1/din[2] qr_4t1_mux_top_1/din[1]
+ qr_4t1_mux_top_1/din[0] qr_4t1_mux_top_1/rst qr_4t1_mux_top_1/din_3_dummy qr_4t1_mux_top_1/din_3_dummy
+ qr_4t1_mux_top_1/din_3_dummy qr_4t1_mux_top_1/din_3_dummy dout_p qr_4t1_mux_top_1/mux_out_dummy
+ DVSS: DVDD: qr_4t1_mux_top_1/sky130_fd_sc_hs__dfxtp_2_1/a_1172_124# qr_4t1_mux_top_1/sky130_fd_sc_hs__dfxtp_2_3/a_1217_314#
+ qr_4t1_mux_top_1/sky130_fd_sc_hs__dfxtp_4_1/a_1141_508# qr_4t1_mux_top_1/sky130_fd_sc_hs__dfxtp_2_3/a_695_459#
+ qr_4t1_mux_top_1/sky130_fd_sc_hs__dfxtp_4_3/a_651_503# qr_4t1_mux_top_1/sky130_fd_sc_hs__dfxtp_2_1/a_538_429#
+ qr_4t1_mux_top_1/sky130_fd_sc_hs__mux4_1_1/A0 qr_4t1_mux_top_1/sky130_fd_sc_hs__mux4_1_1/a_264_74#
+ qr_4t1_mux_top_1/sky130_fd_sc_hs__dfxtp_2_1/a_1217_314# qr_4t1_mux_top_1/sky130_fd_sc_hs__mux4_1_1/a_1338_125#
+ qr_4t1_mux_top_1/sky130_fd_sc_hs__mux4_4_1/a_758_306# qr_4t1_mux_top_1/sky130_fd_sc_hs__mux4_1_1/A2
+ qr_4t1_mux_top_1/sky130_fd_sc_hs__dfxtp_2_7/a_206_368# qr_4t1_mux_top_1/sky130_fd_sc_hs__dfxtp_2_5/a_431_508#
+ qr_4t1_mux_top_1/sky130_fd_sc_hs__mux4_1_1/A1 qr_4t1_mux_top_1/sky130_fd_sc_hs__dfxtp_2_7/D
+ qr_4t1_mux_top_1/sky130_fd_sc_hs__dfxtp_4_1/a_206_368# qr_4t1_mux_top_1/sky130_fd_sc_hs__dfxtp_2_7/a_708_101#
+ qr_4t1_mux_top_1/sky130_fd_sc_hs__dfxtp_4_3/a_696_458# qr_4t1_mux_top_1/sky130_fd_sc_hs__dfxtp_2_9/a_644_504#
+ qr_4t1_mux_top_1/sky130_fd_sc_hs__mux4_1_1/X qr_4t1_mux_top_1/sky130_fd_sc_hs__dfxtp_2_11/a_206_368#
+ qr_4t1_mux_top_1/sky130_fd_sc_hs__dfxtp_4_1/a_437_503# qr_4t1_mux_top_1/sky130_fd_sc_hs__clkbuf_1_1/a_27_74#
+ qr_4t1_mux_top_1/sky130_fd_sc_hs__dfxtp_2_3/a_431_508# qr_4t1_mux_top_1/sky130_fd_sc_hs__dfxtp_4_3/a_544_485#
+ qr_4t1_mux_top_1/sky130_fd_sc_hs__dfxtp_2_9/a_538_429# qr_4t1_mux_top_1/sky130_fd_sc_hs__dfxtp_2_11/a_708_101#
+ qr_4t1_mux_top_1/sky130_fd_sc_hs__dfxtp_2_11/a_1125_508# qr_4t1_mux_top_1/sky130_fd_sc_hs__mux4_1_1/a_27_74#
+ qr_4t1_mux_top_1/sky130_fd_sc_hs__mux4_1_1/a_342_74# qr_4t1_mux_top_1/sky130_fd_sc_hs__dfxtp_2_11/a_27_74#
+ qr_4t1_mux_top_1/sky130_fd_sc_hs__dfxtp_2_1/a_695_459# qr_4t1_mux_top_1/sky130_fd_sc_hs__dfxtp_4_1/a_651_503#
+ qr_4t1_mux_top_1/sky130_fd_sc_hs__dfxtp_4_1/D qr_4t1_mux_top_1/sky130_fd_sc_hs__dfxtp_2_7/a_644_504#
+ qr_4t1_mux_top_1/sky130_fd_sc_hs__dfxtp_4_3/a_1178_124# qr_4t1_mux_top_1/sky130_fd_sc_hs__clkbuf_2_1/a_43_192#
+ qr_4t1_mux_top_1/sky130_fd_sc_hs__dfxtp_2_5/a_206_368# qr_4t1_mux_top_1/sky130_fd_sc_hs__clkbuf_1_5/X
+ qr_4t1_mux_top_1/sky130_fd_sc_hs__dfxtp_2_9/a_1125_508# qr_4t1_mux_top_1/sky130_fd_sc_hs__clkbuf_2_3/X
+ qr_4t1_mux_top_1/sky130_fd_sc_hs__dfxtp_2_7/a_538_429# qr_4t1_mux_top_1/sky130_fd_sc_hs__dfxtp_2_9/Q
+ qr_4t1_mux_top_1/sky130_fd_sc_hs__dfxtp_4_1/a_1178_124# qr_4t1_mux_top_1/sky130_fd_sc_hs__dfxtp_2_11/a_644_504#
+ qr_4t1_mux_top_1/sky130_fd_sc_hs__dfxtp_4_1/a_696_458# qr_4t1_mux_top_1/sky130_fd_sc_hs__dfxtp_2_5/a_27_74#
+ qr_4t1_mux_top_1/sky130_fd_sc_hs__dfxtp_2_5/a_708_101# qr_4t1_mux_top_1/sky130_fd_sc_hs__dfxtp_4_1/a_27_74#
+ qr_4t1_mux_top_1/sky130_fd_sc_hs__mux4_4_1/a_1285_377# qr_4t1_mux_top_1/sky130_fd_sc_hs__dfxtp_2_7/a_1125_508#
+ qr_4t1_mux_top_1/sky130_fd_sc_hs__mux4_1_1/a_537_341# qr_4t1_mux_top_1/sky130_fd_sc_hs__mux4_1_1/a_255_341#
+ qr_4t1_mux_top_1/sky130_fd_sc_hs__mux4_4_1/A0 qr_4t1_mux_top_1/sky130_fd_sc_hs__clkbuf_1_3/X
+ qr_4t1_mux_top_1/sky130_fd_sc_hs__mux4_1_1/A3 qr_4t1_mux_top_1/sky130_fd_sc_hs__dfxtp_2_11/a_538_429#
+ qr_4t1_mux_top_1/sky130_fd_sc_hs__dfxtp_2_3/a_206_368# qr_4t1_mux_top_1/sky130_fd_sc_hs__dfxtp_2_1/a_431_508#
+ qr_4t1_mux_top_1/sky130_fd_sc_hs__clkbuf_1_1/X qr_4t1_mux_top_1/sky130_fd_sc_hs__dfxtp_2_9/a_695_459#
+ qr_4t1_mux_top_1/sky130_fd_sc_hs__dfxtp_4_1/a_544_485# qr_4t1_mux_top_1/sky130_fd_sc_hs__dfxtp_2_5/a_1125_508#
+ qr_4t1_mux_top_1/sky130_fd_sc_hs__mux4_4_1/A2 qr_4t1_mux_top_1/sky130_fd_sc_hs__dfxtp_2_7/a_27_74#
+ qr_4t1_mux_top_1/sky130_fd_sc_hs__dfxtp_2_3/a_708_101# qr_4t1_mux_top_1/sky130_fd_sc_hs__dfxtp_2_3/a_1125_508#
+ qr_4t1_mux_top_1/sky130_fd_sc_hs__dfxtp_4_3/a_27_74# qr_4t1_mux_top_1/sky130_fd_sc_hs__dfxtp_2_11/a_1019_424#
+ qr_4t1_mux_top_1/sky130_fd_sc_hs__mux4_1_1/a_450_74# qr_4t1_mux_top_1/sky130_fd_sc_hs__dfxtp_4_3/a_1034_424#
+ qr_4t1_mux_top_1/sky130_fd_sc_hs__clkbuf_1_3/a_27_74# qr_4t1_mux_top_1/sky130_fd_sc_hs__dfxtp_2_1/a_1125_508#
+ qr_4t1_mux_top_1/sky130_fd_sc_hs__mux4_4_1/a_114_126# qr_4t1_mux_top_1/sky130_fd_sc_hs__dfxtp_2_1/a_27_74#
+ qr_4t1_mux_top_1/sky130_fd_sc_hs__dfxtp_2_5/a_644_504# qr_4t1_mux_top_1/sky130_fd_sc_hs__dfxtp_4_1/a_1034_424#
+ qr_4t1_mux_top_1/sky130_fd_sc_hs__dfxtp_2_11/a_1172_124# qr_4t1_mux_top_1/sky130_fd_sc_hs__mux4_4_1/a_1450_121#
+ qr_4t1_mux_top_1/sky130_fd_sc_hs__dfxtp_2_9/a_431_508# qr_4t1_mux_top_1/sky130_fd_sc_hs__dfxtp_2_7/a_695_459#
+ qr_4t1_mux_top_1/sky130_fd_sc_hs__mux4_4_1/a_1191_121# qr_4t1_mux_top_1/sky130_fd_sc_hs__mux4_1_1/a_768_74#
+ qr_4t1_mux_top_1/sky130_fd_sc_hs__dfxtp_2_5/a_538_429# qr_4t1_mux_top_1/sky130_fd_sc_hs__dfxtp_2_9/a_1019_424#
+ qr_4t1_mux_top_1/sky130_fd_sc_hs__mux4_1_1/a_1396_99# qr_4t1_mux_top_1/sky130_fd_sc_hs__dfxtp_2_3/a_644_504#
+ qr_4t1_mux_top_1/sky130_fd_sc_hs__mux4_1_1/a_1065_387# qr_4t1_mux_top_1/sky130_fd_sc_hs__dfxtp_4_3/a_735_102#
+ qr_4t1_mux_top_1/sky130_fd_sc_hs__dfxtp_2_3/a_27_74# qr_4t1_mux_top_1/sky130_fd_sc_hs__dfxtp_2_11/a_695_459#
+ qr_4t1_mux_top_1/sky130_fd_sc_hs__dfxtp_2_11/a_1217_314# qr_4t1_mux_top_1/sky130_fd_sc_hs__dfxtp_2_7/a_1019_424#
+ qr_4t1_mux_top_1/sky130_fd_sc_hs__dfxtp_2_1/a_206_368# qr_4t1_mux_top_1/sky130_fd_sc_hs__mux4_4_1/a_1278_121#
+ qr_4t1_mux_top_1/sky130_fd_sc_hs__dfxtp_2_3/a_538_429# qr_4t1_mux_top_1/sky130_fd_sc_hs__dfxtp_4_3/a_1226_296#
+ qr_4t1_mux_top_1/sky130_fd_sc_hs__dfxtp_2_1/a_708_101# qr_4t1_mux_top_1/sky130_fd_sc_hs__dfxtp_2_9/a_1172_124#
+ qr_4t1_mux_top_1/sky130_fd_sc_hs__mux4_4_1/a_509_392# qr_4t1_mux_top_1/sky130_fd_sc_hs__dfxtp_2_5/a_1019_424#
+ qr_4t1_mux_top_1/sky130_fd_sc_hs__dfxtp_2_3/a_1019_424# qr_4t1_mux_top_1/sky130_fd_sc_hs__dfxtp_2_7/a_431_508#
+ qr_4t1_mux_top_1/sky130_fd_sc_hs__dfxtp_2_7/a_1172_124# qr_4t1_mux_top_1/sky130_fd_sc_hs__dfxtp_4_1/a_1226_296#
+ qr_4t1_mux_top_1/sky130_fd_sc_hs__mux4_4_1/a_1465_377# qr_4t1_mux_top_1/sky130_fd_sc_hs__mux4_1_1/a_846_74#
+ qr_4t1_mux_top_1/sky130_fd_sc_hs__mux4_4_1/a_2199_74# qr_4t1_mux_top_1/sky130_fd_sc_hs__dfxtp_2_9/a_1217_314#
+ qr_4t1_mux_top_1/sky130_fd_sc_hs__dfxtp_4_3/a_206_368# qr_4t1_mux_top_1/sky130_fd_sc_hs__clkbuf_2_3/a_43_192#
+ qr_4t1_mux_top_1/sky130_fd_sc_hs__mux4_4_1/a_296_392# qr_4t1_mux_top_1/sky130_fd_sc_hs__dfxtp_2_1/a_1019_424#
+ qr_4t1_mux_top_1/sky130_fd_sc_hs__dfxtp_4_3/a_437_503# qr_4t1_mux_top_1/sky130_fd_sc_hs__dfxtp_2_11/a_431_508#
+ qr_4t1_mux_top_1/sky130_fd_sc_hs__dfxtp_2_5/a_1172_124# qr_4t1_mux_top_1/sky130_fd_sc_hs__dfxtp_2_9/a_27_74#
+ qr_4t1_mux_top_1/sky130_fd_sc_hs__dfxtp_2_7/a_1217_314# qr_4t1_mux_top_1/sky130_fd_sc_hs__dfxtp_2_9/a_206_368#
+ qr_4t1_mux_top_1/sky130_fd_sc_hs__dfxtp_2_3/a_1172_124# qr_4t1_mux_top_1/sky130_fd_sc_hs__dfxtp_2_5/a_695_459#
+ qr_4t1_mux_top_1/sky130_fd_sc_hs__mux4_4_1/a_2489_347# qr_4t1_mux_top_1/sky130_fd_sc_hs__mux4_1_1/a_763_341#
+ qr_4t1_mux_top_1/sky130_fd_sc_hs__dfxtp_4_3/a_1141_508# qr_4t1_mux_top_1/sky130_fd_sc_hs__mux4_4_1/a_299_126#
+ qr_4t1_mux_top_1/sky130_fd_sc_hs__dfxtp_2_9/a_708_101# qr_4t1_mux_top_1/sky130_fd_sc_hs__mux4_4_1/a_116_392#
+ qr_4t1_mux_top_1/sky130_fd_sc_hs__dfxtp_2_1/a_644_504# qr_4t1_mux_top_1/sky130_fd_sc_hs__mux4_1_1/a_979_74#
+ qr_4t1_mux_top_1/sky130_fd_sc_hs__dfxtp_2_5/a_1217_314# qr_4t1_mux_top_1/sky130_fd_sc_hs__dfxtp_4_1/a_735_102#
+ qr_4t1_mux_top_1/sky130_fd_sc_hs__clkbuf_1_5/a_27_74# qr_4t1_mux_top
Xsky130_fd_sc_hs__buf_1_1 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__buf_1_1/A sky130_fd_sc_hs__buf_1_1/X
+ sky130_fd_sc_hs__buf_1_1/a_27_164# sky130_fd_sc_hs__buf_1
Xsky130_fd_sc_hs__inv_4_17 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__inv_4_17/Y sky130_fd_sc_hs__inv_4_17/A
+ sky130_fd_sc_hs__inv_4
Xsky130_fd_sc_hs__inv_4_28 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__inv_4_29/Y sky130_fd_sc_hs__inv_4_29/A
+ sky130_fd_sc_hs__inv_4
Xsky130_fd_sc_hs__inv_4_39 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__inv_4_39/Y sky130_fd_sc_hs__inv_4_39/A
+ sky130_fd_sc_hs__inv_4
Xsky130_fd_sc_hs__conb_1_150 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__conb_1_151/LO
+ sky130_fd_sc_hs__conb_1_151/HI sky130_fd_sc_hs__conb_1_151/a_165_290# sky130_fd_sc_hs__conb_1_151/a_21_290#
+ sky130_fd_sc_hs__conb_1
Xsky130_fd_sc_hs__conb_1_161 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__conb_1_161/LO
+ sky130_fd_sc_hs__conb_1_161/HI sky130_fd_sc_hs__conb_1_161/a_165_290# sky130_fd_sc_hs__conb_1_161/a_21_290#
+ sky130_fd_sc_hs__conb_1
Xsky130_fd_sc_hs__conb_1_172 DVSS: DVDD: DVDD: DVSS: prbs_generator_syn_21/eqn[8]
+ prbs_generator_syn_21/eqn[1] sky130_fd_sc_hs__conb_1_173/a_165_290# sky130_fd_sc_hs__conb_1_173/a_21_290#
+ sky130_fd_sc_hs__conb_1
Xsky130_fd_sc_hs__conb_1_183 DVSS: DVDD: DVDD: DVSS: prbs_generator_syn_23/eqn[8]
+ prbs_generator_syn_23/eqn[1] sky130_fd_sc_hs__conb_1_183/a_165_290# sky130_fd_sc_hs__conb_1_183/a_21_290#
+ sky130_fd_sc_hs__conb_1
Xsky130_fd_sc_hs__conb_1_194 DVSS: DVDD: DVDD: DVSS: prbs_generator_syn_19/eqn[9]
+ sky130_fd_sc_hs__conb_1_195/HI sky130_fd_sc_hs__conb_1_195/a_165_290# sky130_fd_sc_hs__conb_1_195/a_21_290#
+ sky130_fd_sc_hs__conb_1
Xsky130_fd_sc_hs__nand2_1_2 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__or2b_4_3/A sky130_fd_sc_hs__or4_2_1/D
+ sky130_fd_sc_hs__nor2_4_3/Y sky130_fd_sc_hs__nand2_1_3/a_117_74# sky130_fd_sc_hs__nand2_1
Xsky130_fd_sc_hs__einvp_2_150 DVSS: DVDD: DVDD: DVSS: dout_p sky130_fd_sc_hs__einvp_2_99/A
+ sky130_fd_sc_hs__buf_2_155/X sky130_fd_sc_hs__einvp_2_151/a_263_323# sky130_fd_sc_hs__einvp_2_151/a_36_74#
+ sky130_fd_sc_hs__einvp_2_151/a_27_368# sky130_fd_sc_hs__einvp_2
Xsky130_fd_sc_hs__clkbuf_16_11 DVSS: DVDD: DVDD: DVSS: osc_core_1/pi1_l[3] sky130_fd_sc_hs__clkbuf_4_13/X
+ sky130_fd_sc_hs__clkbuf_16_11/a_114_74# sky130_fd_sc_hs__clkbuf_16
Xsky130_fd_sc_hs__clkbuf_16_22 DVSS: DVDD: DVDD: DVSS: osc_core_1/pi1_l[0] sky130_fd_sc_hs__clkbuf_8_5/X
+ sky130_fd_sc_hs__clkbuf_16_23/a_114_74# sky130_fd_sc_hs__clkbuf_16
Xsky130_fd_sc_hs__clkbuf_16_33 DVSS: DVDD: DVDD: DVSS: osc_core_1/pi3_l[0] sky130_fd_sc_hs__clkbuf_16_1/X
+ sky130_fd_sc_hs__clkbuf_16_33/a_114_74# sky130_fd_sc_hs__clkbuf_16
Xsky130_fd_sc_hs__clkbuf_16_44 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__dlrtp_1_9/GATE
+ sky130_fd_sc_hs__clkbuf_2_3/A sky130_fd_sc_hs__clkbuf_16_45/a_114_74# sky130_fd_sc_hs__clkbuf_16
Xsky130_fd_sc_hs__clkbuf_16_55 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__einvp_2_99/A
+ sky130_fd_sc_hs__einvp_2_65/A sky130_fd_sc_hs__clkbuf_16_55/a_114_74# sky130_fd_sc_hs__clkbuf_16
Xsky130_fd_sc_hs__clkbuf_16_66 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__nand2_2_9/B
+ sky130_fd_sc_hs__or2b_2_5/A sky130_fd_sc_hs__clkbuf_16_67/a_114_74# sky130_fd_sc_hs__clkbuf_16
Xsky130_fd_sc_hs__clkbuf_16_77 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__nor4_2_1/A
+ sky130_fd_sc_hs__clkbuf_8_79/X sky130_fd_sc_hs__clkbuf_16_77/a_114_74# sky130_fd_sc_hs__clkbuf_16
Xsky130_fd_sc_hs__clkbuf_16_88 DVSS: DVDD: DVDD: DVSS: qr_4t1_mux_top_1/clk_IB qr_4t1_mux_top_3/clk_IB
+ sky130_fd_sc_hs__clkbuf_16_89/a_114_74# sky130_fd_sc_hs__clkbuf_16
Xsky130_fd_sc_hs__clkbuf_16_99 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__clkbuf_16_99/X
+ sky130_fd_sc_hs__clkbuf_4_123/X sky130_fd_sc_hs__clkbuf_16_99/a_114_74# sky130_fd_sc_hs__clkbuf_16
Xsky130_fd_sc_hs__clkbuf_16_110 DVSS: DVDD: DVDD: DVSS: prbs_generator_syn_31/rst
+ prbs_generator_syn_27/rst sky130_fd_sc_hs__clkbuf_16_111/a_114_74# sky130_fd_sc_hs__clkbuf_16
Xsky130_fd_sc_hs__clkbuf_16_121 DVSS: DVDD: DVDD: DVSS: prbs_generator_syn_31/clk
+ prbs_generator_syn_19/clk sky130_fd_sc_hs__clkbuf_16_121/a_114_74# sky130_fd_sc_hs__clkbuf_16
Xsky130_fd_sc_hs__clkbuf_16_132 DVSS: DVDD: DVDD: DVSS: osc_core_1/pi5_l[0] pi5_con[0]
+ sky130_fd_sc_hs__clkbuf_16_133/a_114_74# sky130_fd_sc_hs__clkbuf_16
Xsky130_fd_sc_hs__nand2_2_18 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__buf_8_3/A sky130_fd_sc_hs__nor2_4_1/B
+ sky130_fd_sc_hs__or2b_2_1/A sky130_fd_sc_hs__nand2_2_19/a_27_74# sky130_fd_sc_hs__nand2_2
Xsky130_fd_sc_hs__nand2_2_29 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__nand2_2_29/Y
+ sky130_fd_sc_hs__nor2_4_1/B sky130_fd_sc_hs__nor2_4_1/A sky130_fd_sc_hs__nand2_2_29/a_27_74#
+ sky130_fd_sc_hs__nand2_2
Xprbs_generator_syn_7 prbs_generator_syn_9/clk prbs_generator_syn_9/rst prbs_generator_syn_7/cke
+ sky130_fd_sc_hs__conb_1_75/LO sky130_fd_sc_hs__conb_1_75/LO sky130_fd_sc_hs__conb_1_75/HI
+ sky130_fd_sc_hs__conb_1_75/HI sky130_fd_sc_hs__conb_1_75/HI sky130_fd_sc_hs__conb_1_75/LO
+ sky130_fd_sc_hs__conb_1_75/LO sky130_fd_sc_hs__conb_1_75/LO sky130_fd_sc_hs__conb_1_75/LO
+ sky130_fd_sc_hs__conb_1_75/LO sky130_fd_sc_hs__conb_1_75/LO sky130_fd_sc_hs__conb_1_73/LO
+ sky130_fd_sc_hs__conb_1_73/LO sky130_fd_sc_hs__conb_1_73/HI sky130_fd_sc_hs__conb_1_73/LO
+ sky130_fd_sc_hs__conb_1_73/LO sky130_fd_sc_hs__conb_1_73/LO sky130_fd_sc_hs__conb_1_73/LO
+ sky130_fd_sc_hs__conb_1_63/HI prbs_generator_syn_7/eqn[0] sky130_fd_sc_hs__conb_1_65/HI
+ sky130_fd_sc_hs__conb_1_65/LO sky130_fd_sc_hs__conb_1_65/HI sky130_fd_sc_hs__conb_1_65/HI
+ sky130_fd_sc_hs__conb_1_77/LO sky130_fd_sc_hs__conb_1_77/LO sky130_fd_sc_hs__conb_1_77/LO
+ sky130_fd_sc_hs__conb_1_79/LO sky130_fd_sc_hs__conb_1_79/LO sky130_fd_sc_hs__conb_1_79/LO
+ sky130_fd_sc_hs__conb_1_79/LO sky130_fd_sc_hs__conb_1_79/LO prbs_generator_syn_7/eqn[31]
+ prbs_generator_syn_7/eqn[31] prbs_generator_syn_7/eqn[31] prbs_generator_syn_7/eqn[28]
+ prbs_generator_syn_7/eqn[28] prbs_generator_syn_7/eqn[28] prbs_generator_syn_7/eqn[28]
+ prbs_generator_syn_7/eqn[28] prbs_generator_syn_7/eqn[28] prbs_generator_syn_7/eqn[28]
+ prbs_generator_syn_7/eqn[21] prbs_generator_syn_7/eqn[20] prbs_generator_syn_7/eqn[21]
+ prbs_generator_syn_7/eqn[21] prbs_generator_syn_7/eqn[21] prbs_generator_syn_7/eqn[21]
+ prbs_generator_syn_7/eqn[21] prbs_generator_syn_7/eqn[21] prbs_generator_syn_7/eqn[21]
+ prbs_generator_syn_7/eqn[9] prbs_generator_syn_7/eqn[9] prbs_generator_syn_7/eqn[9]
+ prbs_generator_syn_7/eqn[9] prbs_generator_syn_7/eqn[8] prbs_generator_syn_7/eqn[8]
+ prbs_generator_syn_7/eqn[8] prbs_generator_syn_7/eqn[8] prbs_generator_syn_7/eqn[8]
+ prbs_generator_syn_7/eqn[8] prbs_generator_syn_7/eqn[8] prbs_generator_syn_7/eqn[1]
+ prbs_generator_syn_7/eqn[0] prbs_generator_syn_9/inj_err sky130_fd_sc_hs__conb_1_73/LO
+ sky130_fd_sc_hs__conb_1_73/LO prbs_generator_syn_7/out DVSS: DVDD: prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_1/a_293_74#
+ prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_15/X prbs_generator_syn_7/sky130_fd_sc_hs__nand2_1_35/B
+ prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_51/Y prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_9/A
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_9/CLK prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_47/a_27_74#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_37/a_1226_296# prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_3/B
+ prbs_generator_syn_7/sky130_fd_sc_hs__nor2b_1_7/a_27_112# prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_29/B
+ prbs_generator_syn_7/sky130_fd_sc_hs__sdlclkp_2_1/a_580_74# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_1/a_1141_508#
+ prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_5/Y prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_41/a_230_79#
+ prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_61/a_138_385# prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_43/a_132_392#
+ prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_3/a_222_392# prbs_generator_syn_7/sky130_fd_sc_hs__nor2b_1_9/a_27_112#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_61/a_27_74# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_35/a_206_368#
+ prbs_generator_syn_7/sky130_fd_sc_hs__nand2_2_3/Y prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_25/B
+ prbs_generator_syn_7/sky130_fd_sc_hs__nand2_1_11/a_117_74# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_67/a_651_503#
+ prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_45/X prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_39/a_696_458#
+ prbs_generator_syn_7/sky130_fd_sc_hs__sdlclkp_2_1/a_1198_74# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_45/a_1034_424#
+ prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_17/a_222_392# prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_55/a_222_392#
+ prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_53/Y prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_35/A
+ prbs_generator_syn_7/m3_13600_1651# prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_59/a_52_123#
+ prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_5/a_293_74# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_35/a_1226_296#
+ prbs_generator_syn_7/sky130_fd_sc_hs__nand2_1_51/B prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_5/a_651_503#
+ prbs_generator_syn_7/sky130_fd_sc_hs__nand2_1_21/B prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_8/a_27_74#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_15/a_27_74# prbs_generator_syn_7/sky130_fd_sc_hs__and2b_2_1/X
+ prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_13/X prbs_generator_syn_7/sky130_fd_sc_hs__nand2_2_3/a_27_74#
+ prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_50/a_138_385# prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_33/a_132_392#
+ prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_1/a_376_368# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_25/a_206_368#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_35/a_437_503# prbs_generator_syn_7/sky130_fd_sc_hs__sdlclkp_2_1/a_708_451#
+ prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_45/a_230_79# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_29/a_696_458#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_32/a_27_74# prbs_generator_syn_7/sky130_fd_sc_hs__nor2b_1_4/Y
+ prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_59/a_293_74# prbs_generator_syn_7/sky130_fd_sc_hs__nand2_1_47/a_117_74#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_73/a_735_102# prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_21/a_112_119#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_23/a_1141_508# prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_25/a_293_74#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_7/Q prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_3/a_112_119#
+ prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_35/B prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_51/X
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_53/a_1178_124# prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_23/a_132_392#
+ prbs_generator_syn_7/sky130_fd_sc_hs__nand2_1_3/B prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_15/a_206_368#
+ prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_63/a_132_392# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_55/a_27_74#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_25/a_437_503# prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_41/a_52_123#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_47/a_651_503# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_73/a_1141_508#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_19/a_696_458# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_57/a_696_458#
+ prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_7/X prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_43/a_1034_424#
+ prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_55/A prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_11/a_112_119#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_21/a_1141_508# prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_35/a_222_392#
+ prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_49/a_230_79# prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_67/Y
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_71/a_27_74# prbs_generator_syn_7/sky130_fd_sc_hs__nand2_1_33/B
+ prbs_generator_syn_7/sky130_fd_sc_hs__conb_1_1/LO prbs_generator_syn_7/sky130_fd_sc_hs__nand2_1_19/a_117_74#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_51/a_1178_124# prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_33/X
+ prbs_generator_syn_7/sky130_fd_sc_hs__nand2_1_29/B prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_41/Y
+ prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_53/a_132_392# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_45/a_206_368#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_15/a_437_503# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_37/a_651_503#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_39/a_544_485# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_53/a_735_102#
+ prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_45/a_52_123# prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_1/B
+ prbs_generator_syn_7/sky130_fd_sc_hs__nand2_2_3/B prbs_generator_syn_7/sky130_fd_sc_hs__clkbuf_16_1/A
+ prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_21/X prbs_generator_syn_7/sky130_fd_sc_hs__nand2_1_25/B
+ prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_39/a_376_368# prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_63/X
+ prbs_generator_syn_7/m3_13600_3481# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_69/a_1178_124#
+ prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_21/a_138_385# prbs_generator_syn_7/sky130_fd_sc_hs__nor2b_1_8/Y
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_19/a_1178_124# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_49/a_27_74#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_45/a_437_503# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_27/a_651_503#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_71/a_1141_508# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_65/a_651_503#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_29/a_544_485# prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_3/a_138_385#
+ prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_55/X prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_43/a_735_102#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_41/a_1034_424# prbs_generator_syn_7/sky130_fd_sc_hs__nand2_1_9/B
+ prbs_generator_syn_7/sky130_fd_sc_hs__nor2b_1_9/Y prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_59/a_1034_424#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_39/a_1141_508# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_33/a_1226_296#
+ prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_49/a_52_123# prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_47/Y
+ prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_43/Y prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_4/a_651_503#
+ prbs_generator_syn_7/sky130_fd_sc_hs__nand2_1_49/B prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_19/A
+ prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_11/a_138_385# prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_5/X
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_63/a_206_368# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_17/a_651_503#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_19/a_544_485# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_55/a_651_503#
+ prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_9/Y prbs_generator_syn_7/sky130_fd_sc_hs__nand2_1_17/B
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_57/a_544_485# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_67/a_696_458#
+ prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_35/X prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_19/a_27_74#
+ prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_45/a_222_392# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_32/a_1226_296#
+ prbs_generator_syn_7/sky130_fd_sc_hs__nand2_1_43/B prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_25/A
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_1/a_206_368# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_49/a_1226_296#
+ prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_1/a_112_119# prbs_generator_syn_7/sky130_fd_sc_hs__or2_1_1/X
+ prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_59/a_376_368# prbs_generator_syn_7/sky130_fd_sc_hs__nand2_1_19/B
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_5/a_696_458# prbs_generator_syn_7/sky130_fd_sc_hs__nor2b_1_1/Y
+ prbs_generator_syn_7/sky130_fd_sc_hs__nor2b_1_5/a_278_368# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_17/a_1178_124#
+ prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_39/X prbs_generator_syn_7/m3_13600_5433#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_63/a_437_503# prbs_generator_syn_7/sky130_fd_sc_hs__nand2_2_5/B
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_23/a_735_102# prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_53/A
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_61/a_735_102# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_57/a_1034_424#
+ prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_63/B prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_37/a_1141_508#
+ prbs_generator_syn_7/sky130_fd_sc_hs__nand2_1_47/B prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_29/X
+ prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_65/Y prbs_generator_syn_7/m3_13600_4701#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_1/a_437_503# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_67/a_1178_124#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_9/a_735_102# prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_13/a_132_392#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_15/a_1178_124# prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_15/A
+ prbs_generator_syn_7/sky130_fd_sc_hs__nand2_1_1/B prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_43/B
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_35/a_651_503# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_8/D
+ prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_29/A prbs_generator_syn_7/sky130_fd_sc_hs__nand2_1_7/B
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_13/a_735_102# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_47/a_696_458#
+ prbs_generator_syn_7/sky130_fd_sc_hs__nand2_1_31/B prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_51/a_735_102#
+ prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_59/X prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_35/a_1141_508#
+ prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_25/a_222_392# prbs_generator_syn_7/sky130_fd_sc_hs__sdlclkp_2_1/a_288_48#
+ prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_55/B prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_17/B
+ prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_43/A prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_7/A
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_65/a_1178_124# prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_59/Y
+ prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_41/X prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_21/a_230_79#
+ prbs_generator_syn_7/sky130_fd_sc_hs__nand2_1_57/a_117_74# prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_1/a_222_392#
+ prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_19/B prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_35/a_293_74#
+ prbs_generator_syn_7/sky130_fd_sc_hs__nand2_1_23/a_117_74# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_73/a_206_368#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_25/a_651_503# prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_1/a_138_385#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_37/a_696_458# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_67/a_544_485#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_43/a_27_74# prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_9/X
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_55/a_1034_424# prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_39/a_112_119#
+ prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_15/a_222_392# prbs_generator_syn_7/sky130_fd_sc_hs__conb_1_1/HI
+ prbs_generator_syn_7/sky130_fd_sc_hs__nand2_1_23/B prbs_generator_syn_7/sky130_fd_sc_hs__nand2_1_53/B
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_9/a_1178_124# prbs_generator_syn_7/sky130_fd_sc_hs__nor2b_1_4/A
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_47/a_1226_296# prbs_generator_syn_7/m3_13600_11045#
+ prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_17/X prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_29/a_376_368#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_5/a_544_485# prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_3/X
+ prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_31/a_132_392# prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_61/A
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_15/a_651_503# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_73/a_437_503#
+ prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_25/a_230_79# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_27/a_696_458#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_65/a_696_458# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_33/a_735_102#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_71/a_735_102# prbs_generator_syn_7/m3_13600_7263#
+ prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_43/a_222_392# prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_50/Y
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_8/a_1178_124# prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_53/B
+ prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_19/a_376_368# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_63/a_1178_124#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_4/a_696_458# prbs_generator_syn_7/sky130_fd_sc_hs__nor2b_1_4/a_278_368#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_13/a_1178_124# prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_61/a_132_392#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_53/a_206_368# prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_21/a_52_123#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_45/a_651_503# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_17/a_696_458#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_47/a_544_485# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_55/a_696_458#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_21/a_735_102# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_37/a_27_74#
+ prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_61/B prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_61/X
+ prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_59/a_112_119# prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_31/A
+ prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_33/a_222_392# prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_29/a_230_79#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_45/a_1226_296# prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_9/a_132_392#
+ prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_5/A prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_57/Y
+ prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_31/X prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_51/a_27_74#
+ prbs_generator_syn_7/sky130_fd_sc_hs__nor2b_1_8/a_27_112# prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_47/a_376_368#
+ prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_53/a_293_74# prbs_generator_syn_7/sky130_fd_sc_hs__nand2_1_43/a_117_74#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_8/a_735_102# prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_21/a_293_74#
+ prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_39/a_138_385# prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_63/Y
+ prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_51/a_132_392# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_43/a_206_368#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_53/a_437_503# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_37/a_544_485#
+ prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_57/X prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_53/a_1034_424#
+ prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_25/a_52_123# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_33/a_1141_508#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_63/Q prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_23/a_222_392#
+ prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_63/a_222_392# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_7/a_1178_124#
+ prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_53/X prbs_generator_syn_7/sky130_fd_sc_hs__nand2_2_5/Y
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_61/a_1178_124# prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_1/a_230_79#
+ prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_43/a_230_79# prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_11/a_230_79#
+ prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_41/a_132_392# prbs_generator_syn_7/sky130_fd_sc_hs__nand2_1_13/a_117_74#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_43/a_437_503# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_27/a_544_485#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_63/a_651_503# prbs_generator_syn_7/sky130_fd_sc_hs__nand2_1_7/a_117_74#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_35/a_696_458# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_65/a_544_485#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_51/a_1034_424# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_41/a_735_102#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_32/a_1141_508# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_49/a_1141_508#
+ prbs_generator_syn_7/sky130_fd_sc_hs__nand2_1_55/B prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_53/a_222_392#
+ prbs_generator_syn_7/sky130_fd_sc_hs__sdlclkp_2_1/a_114_112# prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_9/a_293_74#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_43/a_1226_296# prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_29/a_52_123#
+ prbs_generator_syn_7/sky130_fd_sc_hs__nand2_1_37/B prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_1/a_651_503#
+ prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_27/a_376_368# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_4/a_544_485#
+ prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_67/a_376_368# prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_27/X
+ prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_1/X prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_59/a_138_385#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_29/a_1178_124# prbs_generator_syn_7/m3_13600_2871#
+ prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_5/a_230_79# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_23/a_206_368#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_61/a_206_368# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_17/a_544_485#
+ prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_15/a_230_79# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_25/a_696_458#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_55/a_544_485# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_32/a_735_102#
+ prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_29/a_293_74# prbs_generator_syn_7/sky130_fd_sc_hs__nand2_1_17/a_117_74#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_69/a_1034_424# prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_29/a_112_119#
+ prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_37/X prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_31/B
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_19/a_1034_424# prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_33/A
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_9/a_206_368# prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_57/a_376_368#
+ prbs_generator_syn_7/sky130_fd_sc_hs__sdlclkp_2_1/a_706_317# prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_11/B
+ prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_1/a_52_123# prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_39/B
+ prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_21/a_132_392# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_13/a_206_368#
+ prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_43/a_52_123# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_51/a_206_368#
+ prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_47/X prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_23/a_437_503#
+ prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_11/a_52_123# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_61/a_437_503#
+ prbs_generator_syn_7/sky130_fd_sc_hs__nor2b_1_7/Y prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_51/A
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_15/a_696_458# prbs_generator_syn_7/sky130_fd_sc_hs__nor2b_1_5/Y
+ prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_9/a_230_79# prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_25/X
+ prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_19/a_112_119# prbs_generator_syn_7/sky130_fd_sc_hs__nand2_1_45/B
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_5/a_1178_124# prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_19/a_230_79#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_41/a_1226_296# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_59/a_1226_296#
+ prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_63/a_230_79# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_51/Q
+ prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_7/a_132_392# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_9/a_437_503#
+ prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_46/a_376_368# prbs_generator_syn_7/sky130_fd_sc_hs__nand2_1_33/a_117_74#
+ prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_11/a_293_74# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_27/a_1178_124#
+ prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_11/a_132_392# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_13/a_437_503#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_51/a_437_503# prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_5/a_52_123#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_35/a_544_485# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_73/a_651_503#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_45/a_696_458# prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_15/a_52_123#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_47/a_1141_508# prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_47/a_112_119#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_4/a_1178_124# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_17/a_1034_424#
+ prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_23/B prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_37/a_376_368#
+ prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_15/B prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_7/Y
+ prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_29/a_138_385# prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_33/a_230_79#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_25/a_1178_124# prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_47/a_293_74#
+ prbs_generator_syn_7/sky130_fd_sc_hs__nand2_1_37/a_117_74# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_33/a_206_368#
+ prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_15/a_293_74# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_71/a_206_368#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_25/a_544_485# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_67/a_1034_424#
+ prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_13/a_222_392# prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_9/a_52_123#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_15/a_1034_424# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_57/a_1226_296#
+ prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_19/a_52_123# prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_23/X
+ prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_63/a_52_123# prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_19/a_138_385#
+ prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_9/a_376_368# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_21/a_206_368#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_33/a_437_503# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_71/a_437_503#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_53/a_651_503# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_15/a_544_485#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_63/a_696_458# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_65/a_1034_424#
+ prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_19/a_293_74# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_45/a_1141_508#
+ prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_27/a_112_119# prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_67/a_112_119#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_1/a_1178_124# prbs_generator_syn_7/sky130_fd_sc_hs__conb_1_1/a_21_290#
+ prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_63/a_293_74# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_8/a_206_368#
+ prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_17/a_376_368# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_63/a_27_74#
+ prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_21/A prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_55/a_376_368#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_1/a_696_458# prbs_generator_syn_7/sky130_fd_sc_hs__nor2b_1_1/a_278_368#
+ prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_47/a_138_385# prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_33/a_52_123#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_9/a_1034_424# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_21/a_437_503#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_1/a_27_74# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_43/a_651_503#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_1/Q prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_45/a_544_485#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_69/a_735_102# prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_57/a_112_119#
+ prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_31/a_222_392# prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_13/A
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_55/a_1226_296# prbs_generator_syn_7/sky130_fd_sc_hs__nand2_2_5/a_27_74#
+ prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_53/a_230_79# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_8/a_437_503#
+ prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_67/a_293_74# prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_33/a_293_74#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_7/a_735_102# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_23/a_1178_124#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_41/a_206_368# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_8/a_1034_424#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_63/a_1034_424# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_59/a_735_102#
+ prbs_generator_syn_7/sky130_fd_sc_hs__nand2_1_5/B prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_43/a_1141_508#
+ prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_46/a_112_119# prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_61/a_222_392#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_13/a_1034_424# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_73/a_1178_124#
+ prbs_generator_syn_7/sky130_fd_sc_hs__nand2_1_27/B prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_13/B
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_57/a_27_74# prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_57/a_230_79#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_21/a_1178_124# prbs_generator_syn_7/sky130_fd_sc_hs__nor2b_1_1/a_27_112#
+ prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_27/a_138_385# prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_23/a_230_79#
+ prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_67/a_138_385# prbs_generator_syn_7/sky130_fd_sc_hs__nand2_1_41/B
+ prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_9/a_222_392# prbs_generator_syn_7/sky130_fd_sc_hs__nand2_1_27/a_117_74#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_32/a_206_368# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_23/a_651_503#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_41/a_437_503# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_73/a_27_74#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_61/a_651_503# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_63/a_544_485#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_49/a_735_102# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_73/a_696_458#
+ prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_37/a_112_119# prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_51/a_222_392#
+ prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_43/X prbs_generator_syn_7/sky130_fd_sc_hs__nand2_2_1/B
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_9/a_651_503# prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_53/a_52_123#
+ prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_49/X prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_25/a_376_368#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_1/a_544_485# prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_65/a_376_368#
+ prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_57/a_138_385# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_27/a_27_74#
+ prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_39/a_132_392# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_7/a_1034_424#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_13/a_651_503# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_32/a_437_503#
+ prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_27/a_230_79# prbs_generator_syn_7/m3_13600_12265#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_51/a_651_503# prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_59/B
+ prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_47/A prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_61/a_1034_424#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_41/a_1141_508# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_59/a_1141_508#
+ prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_41/a_222_392# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_53/a_1226_296#
+ prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_3/A prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_71/a_1178_124#
+ prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_9/a_112_119# prbs_generator_syn_7/sky130_fd_sc_hs__nand2_1_3/a_117_74#
+ prbs_generator_syn_7/m3_13600_8483# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_39/a_1178_124#
+ prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_57/a_52_123# prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_46/a_138_385#
+ prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_23/a_52_123# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_67/a_27_74#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_53/a_696_458# prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_17/a_112_119#
+ prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_11/A prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_55/a_112_119#
+ prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_1/A prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_51/a_1226_296#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_29/a_1034_424# prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_59/A
+ prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_23/A prbs_generator_syn_7/sky130_fd_sc_hs__nand2_1_39/B
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_5/a_27_74# prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_57/a_293_74#
+ prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_37/a_138_385# prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_59/a_132_392#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_33/a_651_503# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_71/a_651_503#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_43/a_696_458# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_73/a_544_485#
+ prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_27/a_52_123# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_57/a_1141_508#
+ prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_21/a_222_392# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_35/a_27_74#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_69/a_1226_296# prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_37/B
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_19/a_1226_296# prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_35/a_376_368#
+ prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_47/a_230_79# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_37/a_1178_124#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_5/a_1034_424# prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_49/a_132_392#
+ prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_7/a_222_392# prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_27/a_293_74#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_21/a_651_503# prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_9/a_138_385#
+ prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_11/a_222_392# prbs_generator_syn_7/m3_13600_14095#
+ prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_50/A prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_27/a_1034_424#
+ prbs_generator_syn_7/sky130_fd_sc_hs__nand2_1_13/B prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_8/a_651_503#
+ prbs_generator_syn_7/m3_13600_9703# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_35/a_1178_124#
+ prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_17/a_138_385# prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_55/a_138_385#
+ prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_7/a_230_79# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_4/a_1034_424#
+ prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_7/a_376_368# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_69/a_206_368#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_23/a_696_458# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_53/a_544_485#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_39/a_735_102# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_61/a_696_458#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_55/a_1141_508# prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_25/a_112_119#
+ prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_65/a_112_119# prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_43/a_293_74#
+ prbs_generator_syn_7/sky130_fd_sc_hs__nand2_1_57/B prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_25/a_1034_424#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_7/a_206_368# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_17/a_1226_296#
+ prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_15/a_376_368# prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_53/a_376_368#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_9/a_696_458# prbs_generator_syn_7/m3_13600_431#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_45/a_27_74# prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_47/a_52_123#
+ prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_29/a_132_392# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_59/a_206_368#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_69/a_437_503# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_41/a_651_503#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_43/a_544_485# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_13/a_696_458#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_29/a_735_102# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_51/a_696_458#
+ prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_61/Y prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_67/a_1226_296#
+ prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_5/a_132_392# prbs_generator_syn_7/sky130_fd_sc_hs__and2b_2_1/a_198_48#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_7/a_437_503# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_15/a_1226_296#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_69/a_27_74# prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_46/a_293_74#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_1/a_1034_424# prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_19/a_132_392#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_49/a_206_368# prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_7/a_52_123#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_59/a_437_503# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_32/a_651_503#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_7/a_27_74# prbs_generator_syn_7/sky130_fd_sc_hs__nand2_2_1/a_27_74#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_19/a_735_102# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_57/a_735_102#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_65/a_1226_296# prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_37/A
+ prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_33/a_376_368# prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_37/a_230_79#
+ prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_25/a_138_385# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_39/a_27_74#
+ prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_65/a_138_385# prbs_generator_syn_7/sky130_fd_sc_hs__nor2b_1_9/a_278_368#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_49/a_437_503# prbs_generator_syn_7/sky130_fd_sc_hs__and2b_2_1/a_505_74#
+ prbs_generator_syn_7/sky130_fd_sc_hs__nand2_1_51/a_117_74# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_23/a_544_485#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_33/a_696_458# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_61/a_544_485#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_9/a_1226_296# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_53/a_1141_508#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_71/a_696_458# prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_35/a_112_119#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_23/a_1034_424# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_9/a_544_485#
+ prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_63/a_376_368# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_33/a_1178_124#
+ prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_5/a_376_368# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_13/a_544_485#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_73/a_1034_424# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_21/a_696_458#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_51/a_544_485# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_8/a_1226_296#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_51/a_1141_508# prbs_generator_syn_7/sky130_fd_sc_hs__nand2_1_55/a_117_74#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_21/a_1034_424# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_63/a_1226_296#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_23/a_27_74# prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_7/a_112_119#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_13/a_1226_296# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_8/a_696_458#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_32/a_1178_124# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_49/a_1178_124#
+ prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_37/a_52_123# prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_27/a_132_392#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_71/Q prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_67/a_735_102#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_69/a_1141_508# prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_15/a_112_119#
+ prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_53/a_112_119# prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_39/a_222_392#
+ prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_55/a_230_79# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_19/a_1141_508#
+ prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_37/a_293_74# prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_43/a_376_368#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_5/a_735_102# prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_35/a_138_385#
+ prbs_generator_syn_7/sky130_fd_sc_hs__sdlclkp_2_1/a_114_424# prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_57/a_132_392#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_71/a_1034_424# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_7/a_1226_296#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_33/a_544_485# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_41/a_696_458#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_71/a_544_485# prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_21/B
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_61/a_1226_296# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_39/a_1034_424#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_17/a_27_74# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_9/a_27_74#
+ prbs_generator_syn_7/sky130_fd_sc_hs__nor2b_1_5/a_27_112# prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_47/a_132_392#
+ prbs_generator_syn_7/sky130_fd_sc_hs__nor2b_1_8/a_278_368# prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_9/B
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_39/a_206_368# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_33/a_27_74#
+ prbs_generator_syn_7/sky130_fd_sc_hs__nand2_1_41/a_117_74# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_69/a_651_503#
+ prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_51/a_293_74# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_21/a_544_485#
+ prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_7/a_138_385# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_32/a_696_458#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_47/a_735_102# prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_33/a_112_119#
+ prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_59/a_222_392# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_17/a_1141_508#
+ prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_55/a_52_123# prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_3/a_293_74#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_7/a_651_503# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_29/a_1226_296#
+ prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_23/a_376_368# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_8/a_544_485#
+ prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_47/B prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_47/a_1178_124#
+ prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_15/a_138_385# prbs_generator_syn_7/sky130_fd_sc_hs__sdlclkp_2_1/a_1195_374#
+ prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_53/a_138_385# prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_37/a_132_392#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_29/a_206_368# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_39/a_437_503#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_59/a_651_503# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_37/a_735_102#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_67/a_1141_508# prbs_generator_syn_7/sky130_fd_sc_hs__and2b_2_1/a_27_74#
+ prbs_generator_syn_7/sky130_fd_sc_hs__conb_1_1/a_165_290# prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_55/a_293_74#
+ prbs_generator_syn_7/sky130_fd_sc_hs__nand2_1_45/a_117_74# prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_63/a_112_119#
+ prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_49/a_222_392# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_37/a_1034_424#
+ prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_23/a_293_74# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_15/a_1141_508#
+ prbs_generator_syn_7/sky130_fd_sc_hs__nand2_1_5/a_117_74# prbs_generator_syn_7/m3_13600_13485#
+ prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_5/a_112_119# prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_13/a_376_368#
+ prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_51/a_376_368# prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_7/a_293_74#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_19/a_206_368# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_57/a_206_368#
+ prbs_generator_syn_7/sky130_fd_sc_hs__sdlclkp_2_1/a_318_74# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_29/a_437_503#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_49/a_651_503# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_25/a_27_74#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_5/a_1226_296# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_41/a_544_485#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_27/a_735_102# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_65/a_1141_508#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_65/a_735_102# prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_3/a_230_79#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_35/a_1034_424# prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_13/a_230_79#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_41/a_27_74# prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_3/a_132_392#
+ prbs_generator_syn_7/sky130_fd_sc_hs__nand2_1_49/a_117_74# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_27/a_1226_296#
+ prbs_generator_syn_7/sky130_fd_sc_hs__nand2_1_15/a_117_74# prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_41/a_376_368#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_45/a_1178_124# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_4/a_735_102#
+ prbs_generator_syn_7/sky130_fd_sc_hs__nand2_1_9/a_117_74# prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_33/a_138_385#
+ prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_17/a_132_392# prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_55/a_132_392#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_9/a_1141_508# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_19/a_437_503#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_57/a_437_503# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_4/a_1226_296#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_32/a_544_485# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_17/a_735_102#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_55/a_735_102# prbs_generator_syn_7/m3_13600_2261#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_65/a_27_74# prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_29/a_222_392#
+ prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_43/a_112_119# prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_19/X
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_25/a_1226_296# prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_31/a_376_368#
+ prbs_generator_syn_7/sky130_fd_sc_hs__or2_1_1/a_63_368# prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_17/a_230_79#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_4/a_27_74# prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_61/a_230_79#
+ prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_63/a_138_385# prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_5/a_222_392#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_8/a_1141_508# prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_41/a_293_74#
+ prbs_generator_syn_7/sky130_fd_sc_hs__nand2_1_31/a_117_74# prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_5/a_138_385#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_63/a_1141_508# prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_19/a_222_392#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_13/a_1141_508# prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_3/a_52_123#
+ prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_13/a_52_123# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_43/a_1178_124#
+ prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_61/a_376_368# prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_35/a_132_392#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_67/a_206_368# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_1/a_1226_296#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_69/a_696_458# prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_31/a_230_79#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_35/a_735_102# prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_23/a_112_119#
+ prbs_generator_syn_7/sky130_fd_sc_hs__nand2_1_35/a_117_74# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_59/a_27_74#
+ prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_13/a_293_74# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_5/a_206_368#
+ prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_50/a_376_368# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_7/a_696_458#
+ prbs_generator_syn_7/sky130_fd_sc_hs__nor2b_1_7/a_278_368# prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_17/a_52_123#
+ prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_43/a_138_385# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_7/a_1141_508#
+ prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_61/a_52_123# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_67/a_437_503#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_61/a_1141_508# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_25/a_735_102#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_59/a_696_458# prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_13/a_112_119#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_33/a_1034_424# prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_51/a_112_119#
+ prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_35/a_230_79# prbs_generator_syn_7/m3_13600_4091#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_23/a_1226_296# prbs_generator_syn_7/sky130_fd_sc_hs__nand2_1_39/a_117_74#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_29/a_27_74# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_5/a_437_503#
+ prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_17/a_293_74# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_41/a_1178_124#
+ prbs_generator_syn_7/sky130_fd_sc_hs__or2_1_1/a_152_368# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_59/a_1178_124#
+ prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_61/a_293_74# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_47/a_206_368#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_39/a_651_503# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_49/a_696_458#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_15/a_735_102# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_32/a_1034_424#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_73/a_1226_296# prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_27/a_222_392#
+ prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_41/a_112_119# prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_31/a_52_123#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_49/a_1034_424# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_29/a_1141_508#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_21/a_1226_296# prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_39/a_230_79#
+ prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_23/a_138_385# prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_51/a_230_79#
+ prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_45/a_132_392# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_37/a_206_368#
+ prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_65/a_293_74# prbs_generator_syn_7/sky130_fd_sc_hs__nand2_1_53/a_117_74#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_47/a_437_503# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_29/a_651_503#
+ prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_31/a_293_74# prbs_generator_syn_7/sky130_fd_sc_hs__nand2_1_21/a_117_74#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_69/a_544_485# prbs_generator_syn_7/sky130_fd_sc_hs__clkbuf_16_1/a_114_74#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_45/a_735_102# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_13/a_27_74#
+ prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_31/a_112_119# prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_57/a_222_392#
+ prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_35/a_52_123# prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_21/a_376_368#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_7/a_544_485# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_57/a_1178_124#
+ prbs_generator_syn_7/m3_13600_6043# prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_13/a_138_385#
+ prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_51/a_138_385# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_5/a_1141_508#
+ prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_3/a_376_368# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_27/a_206_368#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_65/a_206_368# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_37/a_437_503#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_19/a_651_503# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_57/a_651_503#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_59/a_544_485# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_71/a_1226_296#
+ prbs_generator_syn_7/sky130_fd_sc_hs__nand2_1_25/a_117_74# prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_61/a_112_119#
+ prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_47/a_222_392# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_27/a_1141_508#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_53/a_27_74# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_4/a_206_368#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_39/a_1226_296# prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_11/a_376_368#
+ prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_39/a_52_123# prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_41/a_138_385#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_4/a_1141_508# prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_25/a_132_392#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_17/a_206_368# prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_41/A
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_55/a_206_368# prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_51/a_52_123#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_27/a_437_503# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_65/a_437_503#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_49/a_544_485# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_63/a_735_102#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_47/a_1034_424# prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_50/a_112_119#
+ prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_37/a_222_392# prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_59/a_230_79#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_25/a_1141_508# prbs_generator_syn_7/sky130_fd_sc_hs__nor2b_1_4/a_27_112#
+ prbs_generator_syn_7/sky130_fd_sc_hs__sdlclkp_2_1/a_685_81# prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_1/a_132_392#
+ prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_39/a_293_74# prbs_generator_syn_7/sky130_fd_sc_hs__nand2_1_29/a_117_74#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_4/a_437_503# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_55/a_1178_124#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_21/a_27_74# prbs_generator_syn_7/m3_13600_12875#
+ prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_50/a_293_74# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_1/a_735_102#
+ prbs_generator_syn_7/sky130_fd_sc_hs__xnor2_1_31/a_138_385# prbs_generator_syn_7/sky130_fd_sc_hs__a22o_1_15/a_132_392#
+ prbs_generator_syn_7/sky130_fd_sc_hs__nand2_1_1/a_117_74# prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_17/a_437_503#
+ prbs_generator_syn_7/sky130_fd_sc_hs__dfxtp_4_55/a_437_503# prbs_generator_syn
Xsky130_fd_sc_hs__clkbuf_4_110 DVSS: DVDD: DVDD: DVSS: inj_en osc_core_1/inj_en sky130_fd_sc_hs__clkbuf_4_111/a_83_270#
+ sky130_fd_sc_hs__clkbuf_4
Xsky130_fd_sc_hs__clkbuf_4_121 DVSS: DVDD: DVDD: DVSS: CTL_BUF_P[0] sky130_fd_sc_hs__clkbuf_8_79/A
+ sky130_fd_sc_hs__clkbuf_4_121/a_83_270# sky130_fd_sc_hs__clkbuf_4
Xsky130_fd_sc_hs__clkbuf_4_132 DVSS: DVDD: DVDD: DVSS: inj_error sky130_fd_sc_hs__clkbuf_8_91/A
+ sky130_fd_sc_hs__clkbuf_4_133/a_83_270# sky130_fd_sc_hs__clkbuf_4
Xsky130_fd_sc_hs__o21ai_2_1 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__inv_4_11/Y sky130_fd_sc_hs__o21ai_2_3/A2
+ sky130_fd_sc_hs__nand2_2_3/B sky130_fd_sc_hs__buf_2_39/A sky130_fd_sc_hs__o21ai_2_1/a_116_368#
+ sky130_fd_sc_hs__o21ai_2_1/a_27_74# sky130_fd_sc_hs__o21ai_2
Xsky130_fd_sc_hs__clkdlyinv5sd2_1_6 DVSS: DVDD: DVSS: DVDD: dout_n sky130_fd_sc_hs__and2_2_1/A
+ sky130_fd_sc_hs__clkdlyinv5sd2_1_7/a_28_74# sky130_fd_sc_hs__clkdlyinv5sd2_1_7/a_682_74#
+ sky130_fd_sc_hs__clkdlyinv5sd2_1_7/a_549_74# sky130_fd_sc_hs__clkdlyinv5sd2_1_7/a_288_74#
+ sky130_fd_sc_hs__clkdlyinv5sd2_1
Xsky130_fd_sc_hs__clkbuf_4_50 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__clkbuf_4_51/A
+ sky130_fd_sc_hs__clkbuf_8_29/A sky130_fd_sc_hs__clkbuf_4_51/a_83_270# sky130_fd_sc_hs__clkbuf_4
Xsky130_fd_sc_hs__clkbuf_4_61 DVSS: DVDD: DVDD: DVSS: fine_control_avg_window_select[3]
+ sky130_fd_sc_hs__clkbuf_4_61/X sky130_fd_sc_hs__clkbuf_4_61/a_83_270# sky130_fd_sc_hs__clkbuf_4
Xsky130_fd_sc_hs__clkbuf_4_72 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__or2b_4_5/X
+ sky130_fd_sc_hs__o21ai_2_3/A2 sky130_fd_sc_hs__clkbuf_4_73/a_83_270# sky130_fd_sc_hs__clkbuf_4
Xsky130_fd_sc_hs__clkbuf_4_83 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__nand2_2_15/Y
+ sky130_fd_sc_hs__dlrtp_1_24/D sky130_fd_sc_hs__clkbuf_4_83/a_83_270# sky130_fd_sc_hs__clkbuf_4
Xsky130_fd_sc_hs__clkbuf_4_94 DVSS: DVDD: DVDD: DVSS: div_ratio_half[2] sky130_fd_sc_hs__clkbuf_4_95/X
+ sky130_fd_sc_hs__clkbuf_4_95/a_83_270# sky130_fd_sc_hs__clkbuf_4
Xsky130_fd_sc_hs__o21ai_2_19 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__inv_4_17/Y sky130_fd_sc_hs__o21ai_2_23/A2
+ sky130_fd_sc_hs__nand2_2_7/A sky130_fd_sc_hs__o21ai_2_19/Y sky130_fd_sc_hs__o21ai_2_19/a_116_368#
+ sky130_fd_sc_hs__o21ai_2_19/a_27_74# sky130_fd_sc_hs__o21ai_2
Xqr_4t1_mux_top_2 qr_4t1_mux_top_3/clk_Q hr_16t4_mux_top_3/clk qr_4t1_mux_top_3/clk_I
+ qr_4t1_mux_top_3/clk_IB qr_4t1_mux_top_3/din[3] qr_4t1_mux_top_3/din[2] qr_4t1_mux_top_3/din[1]
+ qr_4t1_mux_top_3/din[0] qr_4t1_mux_top_3/rst qr_4t1_mux_top_3/din_3_dummy qr_4t1_mux_top_3/din_3_dummy
+ qr_4t1_mux_top_3/din_3_dummy qr_4t1_mux_top_3/din_3_dummy dout_n qr_4t1_mux_top_3/mux_out_dummy
+ DVSS: DVDD: qr_4t1_mux_top_3/sky130_fd_sc_hs__dfxtp_2_1/a_1172_124# qr_4t1_mux_top_3/sky130_fd_sc_hs__dfxtp_2_3/a_1217_314#
+ qr_4t1_mux_top_3/sky130_fd_sc_hs__dfxtp_4_1/a_1141_508# qr_4t1_mux_top_3/sky130_fd_sc_hs__dfxtp_2_3/a_695_459#
+ qr_4t1_mux_top_3/sky130_fd_sc_hs__dfxtp_4_3/a_651_503# qr_4t1_mux_top_3/sky130_fd_sc_hs__dfxtp_2_1/a_538_429#
+ qr_4t1_mux_top_3/sky130_fd_sc_hs__mux4_1_1/A0 qr_4t1_mux_top_3/sky130_fd_sc_hs__mux4_1_1/a_264_74#
+ qr_4t1_mux_top_3/sky130_fd_sc_hs__dfxtp_2_1/a_1217_314# qr_4t1_mux_top_3/sky130_fd_sc_hs__mux4_1_1/a_1338_125#
+ qr_4t1_mux_top_3/sky130_fd_sc_hs__mux4_4_1/a_758_306# qr_4t1_mux_top_3/sky130_fd_sc_hs__mux4_1_1/A2
+ qr_4t1_mux_top_3/sky130_fd_sc_hs__dfxtp_2_7/a_206_368# qr_4t1_mux_top_3/sky130_fd_sc_hs__dfxtp_2_5/a_431_508#
+ qr_4t1_mux_top_3/sky130_fd_sc_hs__mux4_1_1/A1 qr_4t1_mux_top_3/sky130_fd_sc_hs__dfxtp_2_7/D
+ qr_4t1_mux_top_3/sky130_fd_sc_hs__dfxtp_4_1/a_206_368# qr_4t1_mux_top_3/sky130_fd_sc_hs__dfxtp_2_7/a_708_101#
+ qr_4t1_mux_top_3/sky130_fd_sc_hs__dfxtp_4_3/a_696_458# qr_4t1_mux_top_3/sky130_fd_sc_hs__dfxtp_2_9/a_644_504#
+ qr_4t1_mux_top_3/sky130_fd_sc_hs__mux4_1_1/X qr_4t1_mux_top_3/sky130_fd_sc_hs__dfxtp_2_11/a_206_368#
+ qr_4t1_mux_top_3/sky130_fd_sc_hs__dfxtp_4_1/a_437_503# qr_4t1_mux_top_3/sky130_fd_sc_hs__clkbuf_1_1/a_27_74#
+ qr_4t1_mux_top_3/sky130_fd_sc_hs__dfxtp_2_3/a_431_508# qr_4t1_mux_top_3/sky130_fd_sc_hs__dfxtp_4_3/a_544_485#
+ qr_4t1_mux_top_3/sky130_fd_sc_hs__dfxtp_2_9/a_538_429# qr_4t1_mux_top_3/sky130_fd_sc_hs__dfxtp_2_11/a_708_101#
+ qr_4t1_mux_top_3/sky130_fd_sc_hs__dfxtp_2_11/a_1125_508# qr_4t1_mux_top_3/sky130_fd_sc_hs__mux4_1_1/a_27_74#
+ qr_4t1_mux_top_3/sky130_fd_sc_hs__mux4_1_1/a_342_74# qr_4t1_mux_top_3/sky130_fd_sc_hs__dfxtp_2_11/a_27_74#
+ qr_4t1_mux_top_3/sky130_fd_sc_hs__dfxtp_2_1/a_695_459# qr_4t1_mux_top_3/sky130_fd_sc_hs__dfxtp_4_1/a_651_503#
+ qr_4t1_mux_top_3/sky130_fd_sc_hs__dfxtp_4_1/D qr_4t1_mux_top_3/sky130_fd_sc_hs__dfxtp_2_7/a_644_504#
+ qr_4t1_mux_top_3/sky130_fd_sc_hs__dfxtp_4_3/a_1178_124# qr_4t1_mux_top_3/sky130_fd_sc_hs__clkbuf_2_1/a_43_192#
+ qr_4t1_mux_top_3/sky130_fd_sc_hs__dfxtp_2_5/a_206_368# qr_4t1_mux_top_3/sky130_fd_sc_hs__clkbuf_1_5/X
+ qr_4t1_mux_top_3/sky130_fd_sc_hs__dfxtp_2_9/a_1125_508# qr_4t1_mux_top_3/sky130_fd_sc_hs__clkbuf_2_3/X
+ qr_4t1_mux_top_3/sky130_fd_sc_hs__dfxtp_2_7/a_538_429# qr_4t1_mux_top_3/sky130_fd_sc_hs__dfxtp_2_9/Q
+ qr_4t1_mux_top_3/sky130_fd_sc_hs__dfxtp_4_1/a_1178_124# qr_4t1_mux_top_3/sky130_fd_sc_hs__dfxtp_2_11/a_644_504#
+ qr_4t1_mux_top_3/sky130_fd_sc_hs__dfxtp_4_1/a_696_458# qr_4t1_mux_top_3/sky130_fd_sc_hs__dfxtp_2_5/a_27_74#
+ qr_4t1_mux_top_3/sky130_fd_sc_hs__dfxtp_2_5/a_708_101# qr_4t1_mux_top_3/sky130_fd_sc_hs__dfxtp_4_1/a_27_74#
+ qr_4t1_mux_top_3/sky130_fd_sc_hs__mux4_4_1/a_1285_377# qr_4t1_mux_top_3/sky130_fd_sc_hs__dfxtp_2_7/a_1125_508#
+ qr_4t1_mux_top_3/sky130_fd_sc_hs__mux4_1_1/a_537_341# qr_4t1_mux_top_3/sky130_fd_sc_hs__mux4_1_1/a_255_341#
+ qr_4t1_mux_top_3/sky130_fd_sc_hs__mux4_4_1/A0 qr_4t1_mux_top_3/sky130_fd_sc_hs__clkbuf_1_3/X
+ qr_4t1_mux_top_3/sky130_fd_sc_hs__mux4_1_1/A3 qr_4t1_mux_top_3/sky130_fd_sc_hs__dfxtp_2_11/a_538_429#
+ qr_4t1_mux_top_3/sky130_fd_sc_hs__dfxtp_2_3/a_206_368# qr_4t1_mux_top_3/sky130_fd_sc_hs__dfxtp_2_1/a_431_508#
+ qr_4t1_mux_top_3/sky130_fd_sc_hs__clkbuf_1_1/X qr_4t1_mux_top_3/sky130_fd_sc_hs__dfxtp_2_9/a_695_459#
+ qr_4t1_mux_top_3/sky130_fd_sc_hs__dfxtp_4_1/a_544_485# qr_4t1_mux_top_3/sky130_fd_sc_hs__dfxtp_2_5/a_1125_508#
+ qr_4t1_mux_top_3/sky130_fd_sc_hs__mux4_4_1/A2 qr_4t1_mux_top_3/sky130_fd_sc_hs__dfxtp_2_7/a_27_74#
+ qr_4t1_mux_top_3/sky130_fd_sc_hs__dfxtp_2_3/a_708_101# qr_4t1_mux_top_3/sky130_fd_sc_hs__dfxtp_2_3/a_1125_508#
+ qr_4t1_mux_top_3/sky130_fd_sc_hs__dfxtp_4_3/a_27_74# qr_4t1_mux_top_3/sky130_fd_sc_hs__dfxtp_2_11/a_1019_424#
+ qr_4t1_mux_top_3/sky130_fd_sc_hs__mux4_1_1/a_450_74# qr_4t1_mux_top_3/sky130_fd_sc_hs__dfxtp_4_3/a_1034_424#
+ qr_4t1_mux_top_3/sky130_fd_sc_hs__clkbuf_1_3/a_27_74# qr_4t1_mux_top_3/sky130_fd_sc_hs__dfxtp_2_1/a_1125_508#
+ qr_4t1_mux_top_3/sky130_fd_sc_hs__mux4_4_1/a_114_126# qr_4t1_mux_top_3/sky130_fd_sc_hs__dfxtp_2_1/a_27_74#
+ qr_4t1_mux_top_3/sky130_fd_sc_hs__dfxtp_2_5/a_644_504# qr_4t1_mux_top_3/sky130_fd_sc_hs__dfxtp_4_1/a_1034_424#
+ qr_4t1_mux_top_3/sky130_fd_sc_hs__dfxtp_2_11/a_1172_124# qr_4t1_mux_top_3/sky130_fd_sc_hs__mux4_4_1/a_1450_121#
+ qr_4t1_mux_top_3/sky130_fd_sc_hs__dfxtp_2_9/a_431_508# qr_4t1_mux_top_3/sky130_fd_sc_hs__dfxtp_2_7/a_695_459#
+ qr_4t1_mux_top_3/sky130_fd_sc_hs__mux4_4_1/a_1191_121# qr_4t1_mux_top_3/sky130_fd_sc_hs__mux4_1_1/a_768_74#
+ qr_4t1_mux_top_3/sky130_fd_sc_hs__dfxtp_2_5/a_538_429# qr_4t1_mux_top_3/sky130_fd_sc_hs__dfxtp_2_9/a_1019_424#
+ qr_4t1_mux_top_3/sky130_fd_sc_hs__mux4_1_1/a_1396_99# qr_4t1_mux_top_3/sky130_fd_sc_hs__dfxtp_2_3/a_644_504#
+ qr_4t1_mux_top_3/sky130_fd_sc_hs__mux4_1_1/a_1065_387# qr_4t1_mux_top_3/sky130_fd_sc_hs__dfxtp_4_3/a_735_102#
+ qr_4t1_mux_top_3/sky130_fd_sc_hs__dfxtp_2_3/a_27_74# qr_4t1_mux_top_3/sky130_fd_sc_hs__dfxtp_2_11/a_695_459#
+ qr_4t1_mux_top_3/sky130_fd_sc_hs__dfxtp_2_11/a_1217_314# qr_4t1_mux_top_3/sky130_fd_sc_hs__dfxtp_2_7/a_1019_424#
+ qr_4t1_mux_top_3/sky130_fd_sc_hs__dfxtp_2_1/a_206_368# qr_4t1_mux_top_3/sky130_fd_sc_hs__mux4_4_1/a_1278_121#
+ qr_4t1_mux_top_3/sky130_fd_sc_hs__dfxtp_2_3/a_538_429# qr_4t1_mux_top_3/sky130_fd_sc_hs__dfxtp_4_3/a_1226_296#
+ qr_4t1_mux_top_3/sky130_fd_sc_hs__dfxtp_2_1/a_708_101# qr_4t1_mux_top_3/sky130_fd_sc_hs__dfxtp_2_9/a_1172_124#
+ qr_4t1_mux_top_3/sky130_fd_sc_hs__mux4_4_1/a_509_392# qr_4t1_mux_top_3/sky130_fd_sc_hs__dfxtp_2_5/a_1019_424#
+ qr_4t1_mux_top_3/sky130_fd_sc_hs__dfxtp_2_3/a_1019_424# qr_4t1_mux_top_3/sky130_fd_sc_hs__dfxtp_2_7/a_431_508#
+ qr_4t1_mux_top_3/sky130_fd_sc_hs__dfxtp_2_7/a_1172_124# qr_4t1_mux_top_3/sky130_fd_sc_hs__dfxtp_4_1/a_1226_296#
+ qr_4t1_mux_top_3/sky130_fd_sc_hs__mux4_4_1/a_1465_377# qr_4t1_mux_top_3/sky130_fd_sc_hs__mux4_1_1/a_846_74#
+ qr_4t1_mux_top_3/sky130_fd_sc_hs__mux4_4_1/a_2199_74# qr_4t1_mux_top_3/sky130_fd_sc_hs__dfxtp_2_9/a_1217_314#
+ qr_4t1_mux_top_3/sky130_fd_sc_hs__dfxtp_4_3/a_206_368# qr_4t1_mux_top_3/sky130_fd_sc_hs__clkbuf_2_3/a_43_192#
+ qr_4t1_mux_top_3/sky130_fd_sc_hs__mux4_4_1/a_296_392# qr_4t1_mux_top_3/sky130_fd_sc_hs__dfxtp_2_1/a_1019_424#
+ qr_4t1_mux_top_3/sky130_fd_sc_hs__dfxtp_4_3/a_437_503# qr_4t1_mux_top_3/sky130_fd_sc_hs__dfxtp_2_11/a_431_508#
+ qr_4t1_mux_top_3/sky130_fd_sc_hs__dfxtp_2_5/a_1172_124# qr_4t1_mux_top_3/sky130_fd_sc_hs__dfxtp_2_9/a_27_74#
+ qr_4t1_mux_top_3/sky130_fd_sc_hs__dfxtp_2_7/a_1217_314# qr_4t1_mux_top_3/sky130_fd_sc_hs__dfxtp_2_9/a_206_368#
+ qr_4t1_mux_top_3/sky130_fd_sc_hs__dfxtp_2_3/a_1172_124# qr_4t1_mux_top_3/sky130_fd_sc_hs__dfxtp_2_5/a_695_459#
+ qr_4t1_mux_top_3/sky130_fd_sc_hs__mux4_4_1/a_2489_347# qr_4t1_mux_top_3/sky130_fd_sc_hs__mux4_1_1/a_763_341#
+ qr_4t1_mux_top_3/sky130_fd_sc_hs__dfxtp_4_3/a_1141_508# qr_4t1_mux_top_3/sky130_fd_sc_hs__mux4_4_1/a_299_126#
+ qr_4t1_mux_top_3/sky130_fd_sc_hs__dfxtp_2_9/a_708_101# qr_4t1_mux_top_3/sky130_fd_sc_hs__mux4_4_1/a_116_392#
+ qr_4t1_mux_top_3/sky130_fd_sc_hs__dfxtp_2_1/a_644_504# qr_4t1_mux_top_3/sky130_fd_sc_hs__mux4_1_1/a_979_74#
+ qr_4t1_mux_top_3/sky130_fd_sc_hs__dfxtp_2_5/a_1217_314# qr_4t1_mux_top_3/sky130_fd_sc_hs__dfxtp_4_1/a_735_102#
+ qr_4t1_mux_top_3/sky130_fd_sc_hs__clkbuf_1_5/a_27_74# qr_4t1_mux_top
Xsky130_fd_sc_hs__inv_4_18 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__inv_4_19/Y sky130_fd_sc_hs__inv_4_19/A
+ sky130_fd_sc_hs__inv_4
Xsky130_fd_sc_hs__inv_4_29 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__inv_4_29/Y sky130_fd_sc_hs__inv_4_29/A
+ sky130_fd_sc_hs__inv_4
Xsky130_fd_sc_hs__conb_1_140 DVSS: DVDD: DVDD: DVSS: prbs_generator_syn_15/eqn[30]
+ sky130_fd_sc_hs__conb_1_141/HI sky130_fd_sc_hs__conb_1_141/a_165_290# sky130_fd_sc_hs__conb_1_141/a_21_290#
+ sky130_fd_sc_hs__conb_1
Xsky130_fd_sc_hs__conb_1_151 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__conb_1_151/LO
+ sky130_fd_sc_hs__conb_1_151/HI sky130_fd_sc_hs__conb_1_151/a_165_290# sky130_fd_sc_hs__conb_1_151/a_21_290#
+ sky130_fd_sc_hs__conb_1
Xsky130_fd_sc_hs__conb_1_162 DVSS: DVDD: DVDD: DVSS: prbs_generator_syn_17/eqn[2]
+ prbs_generator_syn_17/eqn[1] sky130_fd_sc_hs__conb_1_163/a_165_290# sky130_fd_sc_hs__conb_1_163/a_21_290#
+ sky130_fd_sc_hs__conb_1
Xsky130_fd_sc_hs__conb_1_173 DVSS: DVDD: DVDD: DVSS: prbs_generator_syn_21/eqn[8]
+ prbs_generator_syn_21/eqn[1] sky130_fd_sc_hs__conb_1_173/a_165_290# sky130_fd_sc_hs__conb_1_173/a_21_290#
+ sky130_fd_sc_hs__conb_1
Xsky130_fd_sc_hs__conb_1_184 DVSS: DVDD: DVDD: DVSS: prbs_generator_syn_29/eqn[9]
+ sky130_fd_sc_hs__conb_1_185/HI sky130_fd_sc_hs__conb_1_185/a_165_290# sky130_fd_sc_hs__conb_1_185/a_21_290#
+ sky130_fd_sc_hs__conb_1
Xsky130_fd_sc_hs__conb_1_195 DVSS: DVDD: DVDD: DVSS: prbs_generator_syn_19/eqn[9]
+ sky130_fd_sc_hs__conb_1_195/HI sky130_fd_sc_hs__conb_1_195/a_165_290# sky130_fd_sc_hs__conb_1_195/a_21_290#
+ sky130_fd_sc_hs__conb_1
Xosc_core_0 osc_core_1/glob_en osc_core_1/delay_con_lsb[4] osc_core_1/delay_con_lsb[3]
+ osc_core_1/delay_con_lsb[2] osc_core_1/delay_con_lsb[1] osc_core_1/delay_con_lsb[0]
+ osc_core_1/delay_con_msb[7] osc_core_1/delay_con_msb[6] osc_core_1/delay_con_msb[5]
+ osc_core_1/delay_con_msb[4] osc_core_1/delay_con_msb[3] osc_core_1/delay_con_msb[2]
+ osc_core_1/delay_con_msb[1] osc_core_1/delay_con_msb[0] osc_core_1/con_perb_5[3]
+ osc_core_1/con_perb_5[2] osc_core_1/con_perb_5[1] osc_core_1/con_perb_5[0] osc_core_1/con_perb_5[3]
+ osc_core_1/con_perb_5[2] osc_core_1/con_perb_5[1] osc_core_1/con_perb_5[0] osc_core_1/con_perb_5[3]
+ osc_core_1/con_perb_5[2] osc_core_1/con_perb_5[1] osc_core_1/con_perb_5[0] osc_core_1/con_perb_5[3]
+ osc_core_1/con_perb_5[2] osc_core_1/con_perb_5[1] osc_core_1/con_perb_5[0] osc_core_1/con_perb_5[3]
+ osc_core_1/con_perb_5[2] osc_core_1/con_perb_5[1] osc_core_1/con_perb_5[0] osc_core_1/ref_clk
+ osc_core_1/pi1_l[3] osc_core_1/pi1_l[2] osc_core_1/pi1_l[1] osc_core_1/pi1_l[0]
+ osc_core_1/pi1_r[3] osc_core_1/pi1_r[2] osc_core_1/pi1_r[1] osc_core_1/pi1_r[0]
+ osc_core_1/pi2_l[3] osc_core_1/pi2_l[2] osc_core_1/pi2_l[1] osc_core_1/pi2_l[0]
+ osc_core_1/pi2_r[3] osc_core_1/pi2_r[2] osc_core_1/pi2_r[1] osc_core_1/pi2_r[0]
+ osc_core_1/pi3_l[3] osc_core_1/pi3_l[2] osc_core_1/pi3_l[1] osc_core_1/pi3_l[0]
+ osc_core_1/pi3_r[3] osc_core_1/pi3_r[2] osc_core_1/pi3_r[1] osc_core_1/pi3_r[0]
+ osc_core_1/pi4_l[3] osc_core_1/pi4_l[2] osc_core_1/pi4_l[1] osc_core_1/pi4_l[0]
+ osc_core_1/pi4_r[3] osc_core_1/pi4_r[2] osc_core_1/pi4_r[1] osc_core_1/pi4_r[0]
+ osc_core_1/pi5_l[3] osc_core_1/pi5_l[2] osc_core_1/pi5_l[1] osc_core_1/pi5_l[0]
+ osc_core_1/pi5_r[3] osc_core_1/pi5_r[2] osc_core_1/pi5_r[1] osc_core_1/pi5_r[0]
+ osc_core_1/osc_000 osc_core_1/osc_036 osc_core_1/osc_072 osc_core_1/osc_108 osc_core_1/osc_144
+ osc_core_1/inj_en osc_core_1/inj_out osc_core_1/osc_hold osc_core_1/p1 osc_core_1/p2
+ osc_core_1/p3 osc_core_1/p4 osc_core_1/p5 DVSS: AVDD osc_core_1/sky130_fd_sc_hs__einvp_2_5/a_36_74#
+ osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_75/X osc_core_1/sky130_fd_sc_hs__nand2_2_93/Y
+ osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_1/X osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_11/a_28_74#
+ osc_core_1/sky130_fd_sc_hs__inv_4_5/Y osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_27/a_289_74#
+ osc_core_1/sky130_fd_sc_hs__nand2_8_9/B osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_7/a_405_138#
+ osc_core_1/sky130_fd_sc_hs__nand2_4_40/a_27_74# osc_core_1/sky130_fd_sc_hs__dfrtp_4_3/a_890_138#
+ osc_core_1/sky130_fd_sc_hs__nand2_1_9/B osc_core_1/sky130_fd_sc_hs__nand2_4_137/a_27_74#
+ osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_56/A osc_core_1/sky130_fd_sc_hs__inv_4_17/Y
+ osc_core_1/sky130_fd_sc_hs__nand2_2_55/Y osc_core_1/sky130_fd_sc_hs__nand2_8_31/a_27_74#
+ osc_core_1/sky130_fd_sc_hs__nand2_4_53/a_27_74# osc_core_1/sky130_fd_sc_hs__nand2_4_123/Y
+ osc_core_1/sky130_fd_sc_hs__einvp_1_1/a_44_549# osc_core_1/sky130_fd_sc_hs__nand2_1_5/a_117_74#
+ osc_core_1/sky130_fd_sc_hs__inv_4_3/Y osc_core_1/sky130_fd_sc_hs__nand2_2_69/a_27_74#
+ osc_core_1/sky130_fd_sc_hs__einvp_2_11/a_263_323# osc_core_1/sky130_fd_sc_hs__einvp_8_3/a_27_368#
+ osc_core_1/sky130_fd_sc_hs__nand2_2_84/B osc_core_1/sky130_fd_sc_hs__a21oi_1_9/a_29_368#
+ osc_core_1/sky130_fd_sc_hs__nand2_4_51/Y osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_68/X
+ osc_core_1/sky130_fd_sc_hs__einvp_4_9/a_473_323# osc_core_1/sky130_fd_sc_hs__nand2_2_109/a_27_74#
+ osc_core_1/sky130_fd_sc_hs__inv_16_3/Y osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_31/X
+ osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_5/A osc_core_1/sky130_fd_sc_hs__nand2_2_45/B
+ osc_core_1/sky130_fd_sc_hs__nand2_2_3/a_27_74# osc_core_1/sky130_fd_sc_hs__einvp_8_14/a_802_323#
+ osc_core_1/sky130_fd_sc_hs__einvp_2_19/a_36_74# osc_core_1/sky130_fd_sc_hs__nand2_4_15/Y
+ osc_core_1/sky130_fd_sc_hs__nand2_4_153/Y osc_core_1/sky130_fd_sc_hs__nand2_4_107/a_27_74#
+ osc_core_1/sky130_fd_sc_hs__and4_2_3/X osc_core_1/sky130_fd_sc_hs__and2_2_1/a_118_74#
+ osc_core_1/sky130_fd_sc_hs__nand2_4_93/a_27_74# osc_core_1/sky130_fd_sc_hs__einvp_1_5/a_44_549#
+ osc_core_1/sky130_fd_sc_hs__nand2_1_9/a_117_74# osc_core_1/sky130_fd_sc_hs__and4_2_3/a_335_74#
+ osc_core_1/sky130_fd_sc_hs__a21oi_1_49/Y osc_core_1/sky130_fd_sc_hs__einvp_1_5/a_310_392#
+ osc_core_1/sky130_fd_sc_hs__einvp_8_5/a_27_368# osc_core_1/sky130_fd_sc_hs__inv_16_9/Y
+ osc_core_1/sky130_fd_sc_hs__nand2_4_45/Y osc_core_1/sky130_fd_sc_hs__a21oi_1_43/a_29_368#
+ osc_core_1/sky130_fd_sc_hs__nand2_2_77/Y osc_core_1/sky130_fd_sc_hs__clkbuf_2_3/A
+ osc_core_1/sky130_fd_sc_hs__nand2_4_9/a_27_74# osc_core_1/sky130_fd_sc_hs__nand2_8_25/a_27_74#
+ osc_core_1/sky130_fd_sc_hs__inv_16_1/Y osc_core_1/sky130_fd_sc_hs__einvp_4_17/a_473_323#
+ osc_core_1/sky130_fd_sc_hs__nand2_2_53/a_27_74# osc_core_1/sky130_fd_sc_hs__inv_16_13/Y
+ osc_core_1/sky130_fd_sc_hs__nand2_4_47/a_27_74# osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_78/a_289_74#
+ osc_core_1/sky130_fd_sc_hs__inv_8_3/A osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_14/a_289_74#
+ osc_core_1/sky130_fd_sc_hs__inv_8_9/A osc_core_1/sky130_fd_sc_hs__nand2_4_75/Y osc_core_1/sky130_fd_sc_hs__nand2_4_61/a_27_74#
+ osc_core_1/sky130_fd_sc_hs__nand2_4_110/Y osc_core_1/sky130_fd_sc_hs__inv_4_9/Y
+ osc_core_1/sky130_fd_sc_hs__einvp_1_9/a_44_549# osc_core_1/sky130_fd_sc_hs__inv_4_7/Y
+ osc_core_1/sky130_fd_sc_hs__einvp_8_8/a_27_368# osc_core_1/sky130_fd_sc_hs__inv_4_23/Y
+ osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_78/a_405_138# osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_45/a_28_74#
+ osc_core_1/sky130_fd_sc_hs__nand2_2_77/a_27_74# osc_core_1/sky130_fd_sc_hs__nand2_2_23/Y
+ osc_core_1/sky130_fd_sc_hs__einvp_8_9/a_27_368# osc_core_1/sky130_fd_sc_hs__clkbuf_4_3/X
+ osc_core_1/sky130_fd_sc_hs__nand2_4_40/Y osc_core_1/sky130_fd_sc_hs__a21oi_1_13/a_29_368#
+ osc_core_1/sky130_fd_sc_hs__nand2_1_3/B osc_core_1/sky130_fd_sc_hs__nand2_8_1/a_27_74#
+ osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_25/X osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_71/X
+ osc_core_1/sky130_fd_sc_hs__nand2_2_21/a_27_74# osc_core_1/sky130_fd_sc_hs__inv_4_1/Y
+ osc_core_1/sky130_fd_sc_hs__nand2_4_87/a_27_74# osc_core_1/sky130_fd_sc_hs__nand2_4_139/Y
+ osc_core_1/sky130_fd_sc_hs__nand2_4_115/a_27_74# osc_core_1/sky130_fd_sc_hs__dlygate4sd2_1_1/a_28_74#
+ osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_17/a_289_74# osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_5/a_405_138#
+ osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_79/A osc_core_1/sky130_fd_sc_hs__clkbuf_2_14/a_43_192#
+ osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_62/a_289_74# osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_35/X
+ osc_core_1/sky130_fd_sc_hs__nand2_2_53/Y osc_core_1/sky130_fd_sc_hs__nand2_4_31/a_27_74#
+ osc_core_1/sky130_fd_sc_hs__nand2_8_19/a_27_74# osc_core_1/sky130_fd_sc_hs__einvp_8_14/a_27_368#
+ osc_core_1/sky130_fd_sc_hs__inv_4_25/Y osc_core_1/sky130_fd_sc_hs__inv_8_1/A osc_core_1/sky130_fd_sc_hs__inv_4_15/Y
+ osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_15/a_28_74# osc_core_1/sky130_fd_sc_hs__nand2_2_47/a_27_74#
+ osc_core_1/sky130_fd_sc_hs__and2_2_3/X osc_core_1/sky130_fd_sc_hs__nand2_2_15/Y
+ osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_3/a_289_74# osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_63/A
+ osc_core_1/sky130_fd_sc_hs__a21oi_1_17/a_29_368# osc_core_1/sky130_fd_sc_hs__nand2_8_33/a_27_74#
+ osc_core_1/sky130_fd_sc_hs__einvp_8_9/a_802_323# osc_core_1/sky130_fd_sc_hs__inv_16_5/Y
+ osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_65/X osc_core_1/sky130_fd_sc_hs__nand2_2_85/Y
+ osc_core_1/sky130_fd_sc_hs__nand2_2_61/a_27_74# osc_core_1/sky130_fd_sc_hs__einvp_2_1/a_263_323#
+ osc_core_1/sky130_fd_sc_hs__nand2_4_155/a_27_74# osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_57/X
+ osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_21/a_405_138# osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_59/a_405_138#
+ osc_core_1/sky130_fd_sc_hs__a21oi_1_47/a_117_74# osc_core_1/sky130_fd_sc_hs__nand2_4_13/Y
+ osc_core_1/sky130_fd_sc_hs__nand2_4_151/Y osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_39/a_28_74#
+ osc_core_1/sky130_fd_sc_hs__nand2_2_61/B osc_core_1/sky130_fd_sc_hs__inv_4_11/Y
+ osc_core_1/sky130_fd_sc_hs__nand2_2_102/a_27_74# osc_core_1/sky130_fd_sc_hs__einvp_2_13/a_27_368#
+ osc_core_1/sky130_fd_sc_hs__einvp_8_15/a_802_323# osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_65/a_289_74#
+ osc_core_1/sky130_fd_sc_hs__nand2_4_71/a_27_74# osc_core_1/sky130_fd_sc_hs__einvp_8_19/a_27_368#
+ osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_53/a_28_74# osc_core_1/sky130_fd_sc_hs__nand2_2_88/a_27_74#
+ osc_core_1/sky130_fd_sc_hs__nand2_2_15/a_27_74# osc_core_1/sky130_fd_sc_hs__nand2_2_5/a_27_74#
+ osc_core_1/sky130_fd_sc_hs__and4_2_3/C osc_core_1/sky130_fd_sc_hs__a21oi_1_45/Y
+ osc_core_1/sky130_fd_sc_hs__nand2_4_110/a_27_74# osc_core_1/sky130_fd_sc_hs__inv_16_7/Y
+ osc_core_1/sky130_fd_sc_hs__einvp_4_5/a_27_368# osc_core_1/sky130_fd_sc_hs__nand2_2_99/B
+ osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_49/a_405_138# osc_core_1/sky130_fd_sc_hs__a21oi_1_33/a_29_368#
+ osc_core_1/sky130_fd_sc_hs__clkbuf_2_1/A osc_core_1/sky130_fd_sc_hs__nand2_2_5/B
+ osc_core_1/sky130_fd_sc_hs__nand2_2_31/a_27_74# osc_core_1/sky130_fd_sc_hs__nand2_4_25/a_27_74#
+ osc_core_1/sky130_fd_sc_hs__inv_4_36/Y osc_core_1/sky130_fd_sc_hs__nand2_2_9/B osc_core_1/sky130_fd_sc_hs__inv_4_39/Y
+ osc_core_1/sky130_fd_sc_hs__nand2_2_9/Y osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_78/a_28_74#
+ osc_core_1/sky130_fd_sc_hs__dfrtp_4_3/a_313_74# osc_core_1/sky130_fd_sc_hs__nand2_2_39/Y
+ osc_core_1/sky130_fd_sc_hs__and4_2_1/a_143_74# osc_core_1/sky130_fd_sc_hs__inv_8_7/A
+ osc_core_1/sky130_fd_sc_hs__nand2_8_27/a_27_74# osc_core_1/sky130_fd_sc_hs__nand2_4_73/Y
+ osc_core_1/sky130_fd_sc_hs__buf_4_1/a_86_260# osc_core_1/sky130_fd_sc_hs__inv_4_33/Y
+ osc_core_1/sky130_fd_sc_hs__dfrtp_4_3/a_494_366# osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_23/a_28_74#
+ osc_core_1/sky130_fd_sc_hs__clkbuf_4_3/a_83_270# osc_core_1/sky130_fd_sc_hs__einvp_1_19/a_310_392#
+ osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_49/X osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_39/a_405_138#
+ osc_core_1/sky130_fd_sc_hs__clkbuf_2_9/a_43_192# osc_core_1/sky130_fd_sc_hs__nand2_8_43/a_27_74#
+ osc_core_1/sky130_fd_sc_hs__nand2_4_35/Y osc_core_1/sky130_fd_sc_hs__einvp_4_9/a_27_368#
+ osc_core_1/sky130_fd_sc_hs__nand2_2_69/Y osc_core_1/sky130_fd_sc_hs__a21oi_1_35/a_29_368#
+ osc_core_1/sky130_fd_sc_hs__nand2_1_1/B osc_core_1/sky130_fd_sc_hs__nand2_2_71/a_27_74#
+ osc_core_1/sky130_fd_sc_hs__inv_4_29/Y osc_core_1/sky130_fd_sc_hs__nand2_4_65/a_27_74#
+ osc_core_1/sky130_fd_sc_hs__nand2_2_43/B osc_core_1/sky130_fd_sc_hs__dfrtp_4_1/a_1647_81#
+ osc_core_1/sky130_fd_sc_hs__nand2_4_137/Y osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_47/a_28_74#
+ osc_core_1/sky130_fd_sc_hs__and4_2_5/a_143_74# osc_core_1/sky130_fd_sc_hs__a21oi_1_32/a_117_74#
+ osc_core_1/sky130_fd_sc_hs__einvp_2_5/a_27_368# osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_45/A
+ osc_core_1/sky130_fd_sc_hs__nand2_2_97/B osc_core_1/sky130_fd_sc_hs__inv_8_5/A osc_core_1/sky130_fd_sc_hs__nand2_2_51/Y
+ osc_core_1/sky130_fd_sc_hs__dfrtp_4_1/a_890_138# osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_29/a_405_138#
+ osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_69/a_405_138# osc_core_1/sky130_fd_sc_hs__nand2_2_97/a_27_74#
+ osc_core_1/sky130_fd_sc_hs__nand2_2_25/a_27_74# osc_core_1/sky130_fd_sc_hs__nand2_2_99/Y
+ osc_core_1/sky130_fd_sc_hs__nand2_4_19/a_27_74# osc_core_1/sky130_fd_sc_hs__nand2_4_117/a_27_74#
+ osc_core_1/sky130_fd_sc_hs__inv_16_9/A osc_core_1/sky130_fd_sc_hs__nand2_4_29/Y
+ osc_core_1/sky130_fd_sc_hs__einvp_8_19/a_27_74# osc_core_1/sky130_fd_sc_hs__nand2_2_85/B
+ osc_core_1/sky130_fd_sc_hs__einvp_2_19/a_263_323# osc_core_1/sky130_fd_sc_hs__dfrtp_4_3/D
+ osc_core_1/sky130_fd_sc_hs__nand2_2_83/Y osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_17/a_28_74#
+ osc_core_1/sky130_fd_sc_hs__einvp_4_7/a_473_323# osc_core_1/sky130_fd_sc_hs__nand2_4_11/Y
+ osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_20/a_405_138# osc_core_1/sky130_fd_sc_hs__a21oi_1_37/a_117_74#
+ osc_core_1/sky130_fd_sc_hs__einvp_2_9/a_27_368# osc_core_1/sky130_fd_sc_hs__nand2_8_37/a_27_74#
+ osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_56/a_289_74# osc_core_1/sky130_fd_sc_hs__inv_4_31/Y
+ osc_core_1/sky130_fd_sc_hs__inv_1_9/Y osc_core_1/sky130_fd_sc_hs__nand2_2_65/a_27_74#
+ osc_core_1/sky130_fd_sc_hs__inv_16_31/A osc_core_1/sky130_fd_sc_hs__einvp_4_7/a_27_74#
+ osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_9/A osc_core_1/sky130_fd_sc_hs__and2_2_1/B
+ osc_core_1/sky130_fd_sc_hs__nand2_4_159/Y osc_core_1/sky130_fd_sc_hs__einvp_1_3/a_318_74#
+ osc_core_1/sky130_fd_sc_hs__nand2_2_71/B osc_core_1/sky130_fd_sc_hs__inv_4_19/Y
+ osc_core_1/sky130_fd_sc_hs__einvp_2_15/a_36_74# osc_core_1/sky130_fd_sc_hs__nand2_2_108/Y
+ osc_core_1/sky130_fd_sc_hs__buf_4_1/X osc_core_1/sky130_fd_sc_hs__nand2_2_73/Y osc_core_1/sky130_fd_sc_hs__einvp_1_3/a_310_392#
+ osc_core_1/sky130_fd_sc_hs__nand2_4_89/Y osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_47/a_405_138#
+ osc_core_1/sky130_fd_sc_hs__nand2_2_19/a_27_74# osc_core_1/sky130_fd_sc_hs__nand2_2_9/a_27_74#
+ osc_core_1/sky130_fd_sc_hs__nand2_2_57/B osc_core_1/sky130_fd_sc_hs__einvp_4_15/a_473_323#
+ osc_core_1/sky130_fd_sc_hs__nand2_2_37/Y osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_59/a_289_74#
+ osc_core_1/sky130_fd_sc_hs__einvp_1_11/a_44_549# osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_71/a_28_74#
+ osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_25/a_289_74# osc_core_1/sky130_fd_sc_hs__clkbuf_2_9/A
+ osc_core_1/sky130_fd_sc_hs__nand2_4_99/a_27_74# osc_core_1/sky130_fd_sc_hs__nand2_4_27/a_27_74#
+ osc_core_1/sky130_fd_sc_hs__nand2_4_71/Y osc_core_1/sky130_fd_sc_hs__dlygate4sd2_1_1/X
+ osc_core_1/sky130_fd_sc_hs__nand2_4_106/Y osc_core_1/sky130_fd_sc_hs__nand2_4_127/a_27_74#
+ osc_core_1/sky130_fd_sc_hs__a21oi_1_1/a_117_74# osc_core_1/sky130_fd_sc_hs__and4_2_5/D
+ osc_core_1/sky130_fd_sc_hs__nand2_4_5/a_27_74# osc_core_1/sky130_fd_sc_hs__einvp_1_7/a_318_74#
+ osc_core_1/sky130_fd_sc_hs__einvp_8_9/a_27_74# osc_core_1/sky130_fd_sc_hs__conb_1_1/LO
+ osc_core_1/sky130_fd_sc_hs__nand2_2_67/Y osc_core_1/sky130_fd_sc_hs__einvp_4_11/a_27_368#
+ osc_core_1/sky130_fd_sc_hs__inv_4_37/Y osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_25/a_28_74#
+ osc_core_1/sky130_fd_sc_hs__einvp_8_2/a_27_368# osc_core_1/sky130_fd_sc_hs__nand3_4_3/a_27_82#
+ osc_core_1/sky130_fd_sc_hs__dfrtp_4_3/a_2010_409# osc_core_1/sky130_fd_sc_hs__einvp_1_15/a_44_549#
+ osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_41/a_28_74# osc_core_1/sky130_fd_sc_hs__nand2_2_73/a_27_74#
+ osc_core_1/sky130_fd_sc_hs__a21oi_1_23/a_117_74# osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_75/a_289_74#
+ osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_3/a_405_138# osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_78/X
+ osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_41/a_289_74# osc_core_1/sky130_fd_sc_hs__a21oi_1_5/a_117_74#
+ osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_68/a_405_138# osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_59/X
+ osc_core_1/sky130_fd_sc_hs__nand2_2_13/Y osc_core_1/sky130_fd_sc_hs__nand2_4_83/a_27_74#
+ osc_core_1/sky130_fd_sc_hs__inv_4_21/Y osc_core_1/sky130_fd_sc_hs__nand2_2_59/Y
+ osc_core_1/sky130_fd_sc_hs__einvp_4_15/a_27_368# osc_core_1/sky130_fd_sc_hs__einvp_4_19/a_27_74#
+ osc_core_1/sky130_fd_sc_hs__nand2_8_7/a_27_74# osc_core_1/sky130_fd_sc_hs__a21oi_1_29/a_29_368#
+ osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_62/X osc_core_1/sky130_fd_sc_hs__nand2_2_99/a_27_74#
+ osc_core_1/sky130_fd_sc_hs__einvp_8_7/a_802_323# osc_core_1/sky130_fd_sc_hs__a21oi_1_42/a_29_368#
+ osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_1/a_28_74# osc_core_1/sky130_fd_sc_hs__nand2_8_15/a_27_74#
+ osc_core_1/sky130_fd_sc_hs__dfrtp_4_1/a_37_78# osc_core_1/sky130_fd_sc_hs__einvp_2_9/a_263_323#
+ osc_core_1/sky130_fd_sc_hs__einvp_1_19/a_44_549# osc_core_1/sky130_fd_sc_hs__nand2_2_88/B
+ osc_core_1/sky130_fd_sc_hs__nand2_2_43/Y osc_core_1/sky130_fd_sc_hs__nand3_4_3/a_456_82#
+ osc_core_1/sky130_fd_sc_hs__and4_2_5/a_56_74# osc_core_1/sky130_fd_sc_hs__nand2_4_57/Y
+ osc_core_1/sky130_fd_sc_hs__nand2_4_39/a_27_74# osc_core_1/sky130_fd_sc_hs__inv_1_7/Y
+ osc_core_1/sky130_fd_sc_hs__nand2_4_135/a_27_74# osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_45/a_289_74#
+ osc_core_1/sky130_fd_sc_hs__a21oi_1_9/a_117_74# osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_21/a_28_74#
+ osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_7/A osc_core_1/sky130_fd_sc_hs__and2_2_1/A
+ osc_core_1/sky130_fd_sc_hs__dfrtp_4_1/a_2010_409# osc_core_1/sky130_fd_sc_hs__einvp_4_1/a_27_74#
+ osc_core_1/sky130_fd_sc_hs__nand2_4_51/a_27_74# osc_core_1/sky130_fd_sc_hs__clkbuf_4_1/A
+ osc_core_1/sky130_fd_sc_hs__nand2_4_151/a_27_74# osc_core_1/sky130_fd_sc_hs__einvp_4_19/a_27_368#
+ osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_35/a_28_74# osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_53/X
+ osc_core_1/sky130_fd_sc_hs__nand2_4_87/Y osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_7/X
+ osc_core_1/sky130_fd_sc_hs__a21oi_1_45/a_29_368# osc_core_1/sky130_fd_sc_hs__nand2_1_5/B
+ osc_core_1/sky130_fd_sc_hs__nand2_2_108/a_27_74# osc_core_1/sky130_fd_sc_hs__nand2_2_79/B
+ osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_1/A osc_core_1/sky130_fd_sc_hs__nand2_2_35/Y
+ osc_core_1/sky130_fd_sc_hs__nand2_2_85/a_27_74# osc_core_1/sky130_fd_sc_hs__nand2_2_13/a_27_74#
+ osc_core_1/sky130_fd_sc_hs__einvp_4_13/a_473_323# osc_core_1/sky130_fd_sc_hs__nand2_4_77/a_27_74#
+ osc_core_1/sky130_fd_sc_hs__nand2_2_1/a_27_74# osc_core_1/sky130_fd_sc_hs__nand2_4_106/a_27_74#
+ osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_49/a_289_74# osc_core_1/sky130_fd_sc_hs__nand2_4_102/Y
+ osc_core_1/sky130_fd_sc_hs__a21oi_1_43/a_117_74# osc_core_1/sky130_fd_sc_hs__bufbuf_8_1/X
+ osc_core_1/sky130_fd_sc_hs__nand2_4_21/a_27_74# osc_core_1/sky130_fd_sc_hs__dfrtp_4_1/a_494_366#
+ osc_core_1/sky130_fd_sc_hs__einvp_8_15/a_27_368# osc_core_1/sky130_fd_sc_hs__einvp_1_17/a_310_392#
+ osc_core_1/sky130_fd_sc_hs__and2_2_3/a_31_74# osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_37/a_405_138#
+ osc_core_1/sky130_fd_sc_hs__nand2_2_65/Y osc_core_1/sky130_fd_sc_hs__nand2_2_37/a_27_74#
+ osc_core_1/sky130_fd_sc_hs__and4_2_1/a_221_74# osc_core_1/sky130_fd_sc_hs__a21oi_1_49/a_29_368#
+ osc_core_1/sky130_fd_sc_hs__clkbuf_2_1/a_43_192# osc_core_1/sky130_fd_sc_hs__einvp_4_1/a_27_368#
+ osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_75/A osc_core_1/sky130_fd_sc_hs__nand2_4_145/a_27_74#
+ osc_core_1/sky130_fd_sc_hs__nand2_4_61/Y osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_21/a_289_74#
+ osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_29/a_28_74# osc_core_1/sky130_fd_sc_hs__a21oi_1_13/a_117_74#
+ osc_core_1/sky130_fd_sc_hs__nand2_2_96/Y osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_31/a_289_74#
+ osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_27/a_405_138# osc_core_1/sky130_fd_sc_hs__nand2_4_60/a_27_74#
+ osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_37/A osc_core_1/sky130_fd_sc_hs__nand2_8_49/a_27_74#
+ osc_core_1/sky130_fd_sc_hs__nand2_4_25/Y osc_core_1/sky130_fd_sc_hs__and4_2_5/a_221_74#
+ osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_7/a_289_74# osc_core_1/sky130_fd_sc_hs__clkbuf_2_5/a_43_192#
+ osc_core_1/sky130_fd_sc_hs__nand2_2_93/a_27_74# osc_core_1/sky130_fd_sc_hs__nand2_4_85/a_27_74#
+ osc_core_1/sky130_fd_sc_hs__nand2_4_15/a_27_74# osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_68/A
+ osc_core_1/sky130_fd_sc_hs__einvp_4_5/a_473_323# osc_core_1/sky130_fd_sc_hs__nand2_4_55/Y
+ osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_17/a_405_138# osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_57/a_405_138#
+ osc_core_1/sky130_fd_sc_hs__inv_1_9/A osc_core_1/sky130_fd_sc_hs__a21oi_1_17/a_117_74#
+ osc_core_1/sky130_fd_sc_hs__nand2_2_89/Y osc_core_1/sky130_fd_sc_hs__einvp_2_17/a_27_368#
+ osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_51/X osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_69/a_289_74#
+ osc_core_1/sky130_fd_sc_hs__einvp_8_8/a_802_323# osc_core_1/sky130_fd_sc_hs__and4_2_3/A
+ osc_core_1/sky130_fd_sc_hs__einvp_8_14/a_27_74# osc_core_1/sky130_fd_sc_hs__dfrtp_4_3/a_699_463#
+ osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_35/a_289_74# osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_3/a_28_74#
+ osc_core_1/sky130_fd_sc_hs__einvp_2_1/a_27_368# osc_core_1/sky130_fd_sc_hs__and4_2_5/C
+ osc_core_1/sky130_fd_sc_hs__nand2_8_17/a_27_74# osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_14/a_28_74#
+ osc_core_1/sky130_fd_sc_hs__conb_1_1/a_21_290# osc_core_1/sky130_fd_sc_hs__nand2_4_139/a_27_74#
+ osc_core_1/sky130_fd_sc_hs__inv_1_1/Y osc_core_1/sky130_fd_sc_hs__clkbuf_2_8/a_43_192#
+ osc_core_1/sky130_fd_sc_hs__einvp_1_1/a_310_392# osc_core_1/sky130_fd_sc_hs__nand2_2_3/Y
+ osc_core_1/sky130_fd_sc_hs__nand2_4_55/a_27_74# osc_core_1/sky130_fd_sc_hs__nand2_2_33/Y
+ osc_core_1/sky130_fd_sc_hs__and4_2_3/a_143_74# osc_core_1/sky130_fd_sc_hs__and4_2_3/B
+ osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_39/a_289_74# osc_core_1/sky130_fd_sc_hs__a21oi_1_33/a_117_74#
+ osc_core_1/sky130_fd_sc_hs__buf_4_1/A osc_core_1/sky130_fd_sc_hs__clkbuf_4_5/a_83_270#
+ osc_core_1/sky130_fd_sc_hs__nand2_2_63/Y osc_core_1/sky130_fd_sc_hs__clkbuf_4_3/A
+ osc_core_1/sky130_fd_sc_hs__a21oi_1_39/a_29_368# osc_core_1/sky130_fd_sc_hs__nand2_4_131/Y
+ osc_core_1/sky130_fd_sc_hs__nand2_4_95/a_27_74# osc_core_1/sky130_fd_sc_hs__nand2_4_123/a_27_74#
+ osc_core_1/sky130_fd_sc_hs__clkbuf_4_5/X osc_core_1/sky130_fd_sc_hs__nand2_4_1/a_27_74#
+ osc_core_1/sky130_fd_sc_hs__clkbuf_1_1/A osc_core_1/sky130_fd_sc_hs__einvp_1_13/a_318_74#
+ osc_core_1/sky130_fd_sc_hs__einvp_8_5/a_27_74# osc_core_1/sky130_fd_sc_hs__a21oi_1_35/a_117_74#
+ osc_core_1/sky130_fd_sc_hs__nand2_1_9/Y osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_53/a_289_74#
+ osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_25/a_405_138# osc_core_1/sky130_fd_sc_hs__nand2_2_55/a_27_74#
+ osc_core_1/sky130_fd_sc_hs__nand2_4_23/Y osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_65/a_405_138#
+ osc_core_1/sky130_fd_sc_hs__nand2_4_49/a_27_74# osc_core_1/sky130_fd_sc_hs__nand2_4_147/a_27_74#
+ osc_core_1/sky130_fd_sc_hs__nand2_8_41/a_27_74# osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_3/A
+ osc_core_1/sky130_fd_sc_hs__and2_2_3/A osc_core_1/sky130_fd_sc_hs__nand2_2_7/B osc_core_1/sky130_fd_sc_hs__nand2_2_19/Y
+ osc_core_1/sky130_fd_sc_hs__einvp_2_17/a_263_323# osc_core_1/sky130_fd_sc_hs__einvp_8_5/a_802_323#
+ osc_core_1/sky130_fd_sc_hs__a21oi_1_21/a_29_368# osc_core_1/sky130_fd_sc_hs__nand2_2_79/a_27_74#
+ osc_core_1/sky130_fd_sc_hs__nand2_4_53/Y osc_core_1/sky130_fd_sc_hs__clkbuf_2_8/A
+ osc_core_1/sky130_fd_sc_hs__and4_2_3/D osc_core_1/sky130_fd_sc_hs__a21oi_1_3/a_29_368#
+ osc_core_1/sky130_fd_sc_hs__einvp_1_17/a_318_74# osc_core_1/sky130_fd_sc_hs__dlygate4sd2_1_1/A
+ osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_56/a_405_138# osc_core_1/sky130_fd_sc_hs__clkbuf_1_1/a_27_74#
+ osc_core_1/sky130_fd_sc_hs__einvp_4_15/a_27_74# osc_core_1/sky130_fd_sc_hs__nand2_8_3/a_27_74#
+ osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_63/a_28_74# osc_core_1/sky130_fd_sc_hs__nand2_2_96/a_27_74#
+ osc_core_1/sky130_fd_sc_hs__nand2_4_89/a_27_74# osc_core_1/sky130_fd_sc_hs__inv_4_13/Y
+ osc_core_1/sky130_fd_sc_hs__nand2_2_49/Y osc_core_1/sky130_fd_sc_hs__einvp_2_1/a_36_74#
+ osc_core_1/sky130_fd_sc_hs__nand2_8_11/a_27_74# osc_core_1/sky130_fd_sc_hs__nand2_2_102/Y
+ osc_core_1/sky130_fd_sc_hs__and2_2_3/B osc_core_1/sky130_fd_sc_hs__dfrtp_4_3/a_124_78#
+ osc_core_1/sky130_fd_sc_hs__nand2_4_83/Y osc_core_1/sky130_fd_sc_hs__and4_2_1/a_56_74#
+ osc_core_1/sky130_fd_sc_hs__nand2_4_33/a_27_74# osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_7/a_28_74#
+ osc_core_1/sky130_fd_sc_hs__nand2_1_3/a_117_74# osc_core_1/sky130_fd_sc_hs__a21oi_1_25/a_29_368#
+ osc_core_1/sky130_fd_sc_hs__nand2_2_31/Y osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_45/a_405_138#
+ osc_core_1/sky130_fd_sc_hs__nand2_2_49/a_27_74# osc_core_1/sky130_fd_sc_hs__a21oi_1_7/a_29_368#
+ osc_core_1/sky130_fd_sc_hs__nand2_2_78/Y osc_core_1/sky130_fd_sc_hs__dlygate4sd2_1_1/a_288_74#
+ osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_31/a_28_74# osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_29/a_289_74#
+ osc_core_1/sky130_fd_sc_hs__clkbuf_2_7/X osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_74/a_289_74#
+ osc_core_1/sky130_fd_sc_hs__nand2_4_157/a_27_74# osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_43/X
+ osc_core_1/sky130_fd_sc_hs__nand2_4_111/Y osc_core_1/sky130_fd_sc_hs__einvp_1_15/a_310_392#
+ osc_core_1/sky130_fd_sc_hs__nand2_4_73/a_27_74# osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_35/a_405_138#
+ osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_75/a_405_138# osc_core_1/sky130_fd_sc_hs__einvp_1_3/a_44_549#
+ osc_core_1/sky130_fd_sc_hs__einvp_4_13/a_27_368# osc_core_1/sky130_fd_sc_hs__nand2_1_7/a_117_74#
+ osc_core_1/sky130_fd_sc_hs__a21oi_1_28/a_29_368# osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_57/a_28_74#
+ osc_core_1/sky130_fd_sc_hs__nand2_4_9/Y osc_core_1/sky130_fd_sc_hs__nand2_2_7/a_27_74#
+ osc_core_1/sky130_fd_sc_hs__dfrtp_4_3/a_1827_81# osc_core_1/sky130_fd_sc_hs__nand2_2_92/Y
+ osc_core_1/sky130_fd_sc_hs__nand2_1_7/Y osc_core_1/sky130_fd_sc_hs__nand2_2_33/a_27_74#
+ osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_33/A osc_core_1/sky130_fd_sc_hs__nand2_2_65/B
+ osc_core_1/sky130_fd_sc_hs__nand2_4_21/Y osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_1/a_405_138#
+ osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_11/a_289_74# osc_core_1/sky130_fd_sc_hs__nand2_4_69/Y
+ osc_core_1/sky130_fd_sc_hs__and2_2_3/a_118_74# osc_core_1/sky130_fd_sc_hs__and4_2_1/X
+ osc_core_1/sky130_fd_sc_hs__nand2_4_41/a_27_74# osc_core_1/sky130_fd_sc_hs__einvp_1_7/a_44_549#
+ osc_core_1/sky130_fd_sc_hs__nand2_4_141/a_27_74# osc_core_1/sky130_fd_sc_hs__nand2_4_121/Y
+ osc_core_1/sky130_fd_sc_hs__nand2_2_17/Y osc_core_1/sky130_fd_sc_hs__einvp_8_7/a_27_368#
+ osc_core_1/sky130_fd_sc_hs__einvp_2_15/a_263_323# osc_core_1/sky130_fd_sc_hs__a21oi_1_11/a_29_368#
+ osc_core_1/sky130_fd_sc_hs__nand2_8_45/a_27_74# osc_core_1/sky130_fd_sc_hs__einvp_2_7/a_263_323#
+ osc_core_1/sky130_fd_sc_hs__nand2_4_99/Y osc_core_1/sky130_fd_sc_hs__nand2_4_67/a_27_74#
+ osc_core_1/sky130_fd_sc_hs__a21oi_1_29/a_117_74# osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_3/X
+ osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_53/a_405_138# osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_47/a_289_74#
+ osc_core_1/sky130_fd_sc_hs__nand2_2_73/B osc_core_1/sky130_fd_sc_hs__dfrtp_4_1/a_699_463#
+ osc_core_1/sky130_fd_sc_hs__a21oi_1_42/a_117_74# osc_core_1/sky130_fd_sc_hs__nand2_2_47/Y
+ osc_core_1/sky130_fd_sc_hs__nand2_4_11/a_27_74# osc_core_1/sky130_fd_sc_hs__nand2_4_81/Y
+ osc_core_1/sky130_fd_sc_hs__nand2_4_115/Y osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_65/a_28_74#
+ osc_core_1/sky130_fd_sc_hs__nand2_2_27/a_27_74# osc_core_1/sky130_fd_sc_hs__einvp_8_8/a_27_74#
+ osc_core_1/sky130_fd_sc_hs__nand2_4_119/a_27_74# osc_core_1/sky130_fd_sc_hs__nand2_4_43/Y
+ osc_core_1/sky130_fd_sc_hs__einvp_2_3/a_36_74# osc_core_1/sky130_fd_sc_hs__a21oi_1_15/a_29_368#
+ osc_core_1/sky130_fd_sc_hs__nand2_8_13/a_27_74# osc_core_1/sky130_fd_sc_hs__and4_2_3/a_56_74#
+ osc_core_1/sky130_fd_sc_hs__nand2_2_43/a_27_74# osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_20/A
+ osc_core_1/sky130_fd_sc_hs__nand2_4_35/a_27_74# osc_core_1/sky130_fd_sc_hs__nand2_2_37/B
+ osc_core_1/sky130_fd_sc_hs__einvp_4_11/a_473_323# osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_9/X
+ osc_core_1/sky130_fd_sc_hs__and4_2_5/B osc_core_1/sky130_fd_sc_hs__nand2_4_145/Y
+ osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_20/a_289_74# osc_core_1/sky130_fd_sc_hs__a21oi_1_45/a_117_74#
+ osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_20/a_28_74# osc_core_1/sky130_fd_sc_hs__clkbuf_2_17/a_43_192#
+ osc_core_1/sky130_fd_sc_hs__nand3_4_3/C osc_core_1/sky130_fd_sc_hs__dfrtp_4_3/a_789_463#
+ osc_core_1/sky130_fd_sc_hs__einvp_8_17/a_27_368# osc_core_1/sky130_fd_sc_hs__nand2_8_39/a_27_74#
+ osc_core_1/sky130_fd_sc_hs__bufbuf_8_1/a_221_368# osc_core_1/sky130_fd_sc_hs__and4_2_3/a_221_74#
+ osc_core_1/sky130_fd_sc_hs__nand2_2_67/a_27_74# osc_core_1/sky130_fd_sc_hs__einvp_4_9/a_27_74#
+ osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_74/a_405_138# osc_core_1/sky130_fd_sc_hs__nand2_2_21/Y
+ osc_core_1/sky130_fd_sc_hs__nand2_4_159/a_27_74# osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_5/a_289_74#
+ osc_core_1/sky130_fd_sc_hs__nand2_4_39/Y osc_core_1/sky130_fd_sc_hs__nand2_4_7/Y
+ osc_core_1/sky130_fd_sc_hs__a21oi_1_19/a_29_368# osc_core_1/sky130_fd_sc_hs__nand2_2_105/a_27_74#
+ osc_core_1/sky130_fd_sc_hs__nand2_2_12/a_27_74# osc_core_1/sky130_fd_sc_hs__nand2_2_84/a_27_74#
+ osc_core_1/sky130_fd_sc_hs__nand2_1_5/Y osc_core_1/sky130_fd_sc_hs__nand2_4_103/a_27_74#
+ osc_core_1/sky130_fd_sc_hs__a21oi_1_49/a_117_74# osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_59/a_28_74#
+ osc_core_1/sky130_fd_sc_hs__einvp_2_15/a_27_368# osc_core_1/sky130_fd_sc_hs__dfrtp_4_1/a_313_74#
+ osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_68/a_289_74# osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_79/X
+ osc_core_1/sky130_fd_sc_hs__inv_1_7/A osc_core_1/sky130_fd_sc_hs__nand2_4_91/a_27_74#
+ osc_core_1/sky130_fd_sc_hs__nand2_4_67/Y osc_core_1/sky130_fd_sc_hs__inv_4_27/Y
+ osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_75/a_28_74# osc_core_1/sky130_fd_sc_hs__clkbuf_4_1/a_83_270#
+ osc_core_1/sky130_fd_sc_hs__einvp_8_3/a_27_74# osc_core_1/sky130_fd_sc_hs__nand2_4_129/a_27_74#
+ osc_core_1/sky130_fd_sc_hs__nand2_8_23/a_27_74# osc_core_1/sky130_fd_sc_hs__nand2_4_7/a_27_74#
+ osc_core_1/sky130_fd_sc_hs__einvp_4_7/a_27_368# osc_core_1/sky130_fd_sc_hs__nand2_2_51/a_27_74#
+ osc_core_1/sky130_fd_sc_hs__dfrtp_4_3/a_834_355# osc_core_1/sky130_fd_sc_hs__nand2_4_45/a_27_74#
+ osc_core_1/sky130_fd_sc_hs__nand2_2_84/Y osc_core_1/sky130_fd_sc_hs__nand2_4_97/Y
+ osc_core_1/sky130_fd_sc_hs__einvp_2_5/a_263_323# osc_core_1/sky130_fd_sc_hs__einvp_4_3/a_473_323#
+ osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_15/a_405_138# osc_core_1/sky130_fd_sc_hs__dfrtp_4_3/a_1627_493#
+ osc_core_1/sky130_fd_sc_hs__einvp_2_19/a_27_368# osc_core_1/sky130_fd_sc_hs__einvp_8_19/a_802_323#
+ osc_core_1/sky130_fd_sc_hs__nand2_2_45/Y osc_core_1/sky130_fd_sc_hs__einvp_2_3/a_27_368#
+ osc_core_1/sky130_fd_sc_hs__dfrtp_4_3/a_812_138# osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_43/a_28_74#
+ osc_core_1/sky130_fd_sc_hs__nand2_4_113/Y osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_53/A
+ osc_core_1/sky130_fd_sc_hs__einvp_4_11/a_27_74# osc_core_1/sky130_fd_sc_hs__nand2_4_41/Y
+ osc_core_1/sky130_fd_sc_hs__nand2_2_92/a_27_74# osc_core_1/sky130_fd_sc_hs__nand2_2_109/Y
+ osc_core_1/sky130_fd_sc_hs__einvp_1_9/a_310_392# osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_43/a_405_138#
+ osc_core_1/sky130_fd_sc_hs__nand2_4_113/a_27_74# osc_core_1/sky130_fd_sc_hs__clkbuf_2_1/X
+ osc_core_1/sky130_fd_sc_hs__nand2_8_9/a_27_74# osc_core_1/sky130_fd_sc_hs__nand2_2_35/B
+ osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_69/a_28_74# osc_core_1/sky130_fd_sc_hs__nand2_2_7/Y
+ osc_core_1/sky130_fd_sc_hs__nand2_4_143/Y osc_core_1/sky130_fd_sc_hs__einvp_8_15/a_27_74#
+ osc_core_1/sky130_fd_sc_hs__einvp_2_7/a_36_74# osc_core_1/sky130_fd_sc_hs__dfrtp_4_3/a_37_78#
+ osc_core_1/sky130_fd_sc_hs__nand2_4_107/Y osc_core_1/sky130_fd_sc_hs__nand2_2_45/a_27_74#
+ osc_core_1/sky130_fd_sc_hs__einvp_1_13/a_310_392# osc_core_1/sky130_fd_sc_hs__dfrtp_4_1/a_1627_493#
+ osc_core_1/sky130_fd_sc_hs__einvp_1_1/a_318_74# osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_33/a_405_138#
+ osc_core_1/sky130_fd_sc_hs__nand2_4_5/Y osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_71/a_405_138#
+ osc_core_1/sky130_fd_sc_hs__einvp_4_3/a_27_74# osc_core_1/sky130_fd_sc_hs__nand2_4_153/a_27_74#
+ osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_37/a_28_74# osc_core_1/sky130_fd_sc_hs__nand2_1_3/Y
+ osc_core_1/sky130_fd_sc_hs__nand2_4_135/Y osc_core_1/sky130_fd_sc_hs__dfrtp_4_1/a_1827_81#
+ osc_core_1/sky130_fd_sc_hs__a21oi_1_39/a_117_74# osc_core_1/sky130_fd_sc_hs__einvp_2_11/a_36_74#
+ osc_core_1/sky130_fd_sc_hs__inv_1_5/A osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_51/a_28_74#
+ osc_core_1/sky130_fd_sc_hs__nand2_4_65/Y osc_core_1/sky130_fd_sc_hs__nand2_4_79/a_27_74#
+ osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_23/a_405_138# osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_63/a_405_138#
+ osc_core_1/sky130_fd_sc_hs__einvp_1_5/a_318_74# osc_core_1/sky130_fd_sc_hs__nand2_4_27/Y
+ osc_core_1/sky130_fd_sc_hs__nand2_4_23/a_27_74# osc_core_1/sky130_fd_sc_hs__nand2_4_121/a_27_74#
+ osc_core_1/sky130_fd_sc_hs__einvp_2_13/a_263_323# osc_core_1/sky130_fd_sc_hs__nand2_4_129/Y
+ osc_core_1/sky130_fd_sc_hs__nand2_2_39/a_27_74# osc_core_1/sky130_fd_sc_hs__nand2_4_95/Y
+ osc_core_1/sky130_fd_sc_hs__clkbuf_2_17/A osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_14/a_405_138#
+ osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_51/a_405_138# osc_core_1/sky130_fd_sc_hs__einvp_1_13/a_44_549#
+ osc_core_1/sky130_fd_sc_hs__a21oi_1_21/a_117_74# osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_71/a_289_74#
+ osc_core_1/sky130_fd_sc_hs__a21oi_1_3/a_117_74# osc_core_1/sky130_fd_sc_hs__einvp_1_9/a_318_74#
+ osc_core_1/sky130_fd_sc_hs__conb_1_1/a_165_290# osc_core_1/sky130_fd_sc_hs__nand2_4_63/a_27_74#
+ osc_core_1/sky130_fd_sc_hs__nand2_2_105/Y osc_core_1/sky130_fd_sc_hs__and4_2_1/a_335_74#
+ osc_core_1/sky130_fd_sc_hs__nand2_2_78/a_27_74# osc_core_1/sky130_fd_sc_hs__nand2_2_5/Y
+ osc_core_1/sky130_fd_sc_hs__nand2_4_141/Y osc_core_1/sky130_fd_sc_hs__dfrtp_4_3/a_1678_395#
+ osc_core_1/sky130_fd_sc_hs__einvp_1_17/a_44_549# osc_core_1/sky130_fd_sc_hs__einvp_4_13/a_27_74#
+ osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_62/a_28_74# osc_core_1/sky130_fd_sc_hs__nand2_2_23/a_27_74#
+ osc_core_1/sky130_fd_sc_hs__nand3_4_1/a_456_82# osc_core_1/sky130_fd_sc_hs__a21oi_1_25/a_117_74#
+ osc_core_1/sky130_fd_sc_hs__nand2_4_17/a_27_74# osc_core_1/sky130_fd_sc_hs__nand2_4_103/Y
+ osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_43/a_289_74# osc_core_1/sky130_fd_sc_hs__dfrtp_4_1/a_789_463#
+ osc_core_1/sky130_fd_sc_hs__a21oi_1_7/a_117_74# osc_core_1/sky130_fd_sc_hs__einvp_8_17/a_27_74#
+ osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_5/a_28_74# osc_core_1/sky130_fd_sc_hs__nand2_4_3/Y
+ osc_core_1/sky130_fd_sc_hs__nand2_4_33/Y osc_core_1/sky130_fd_sc_hs__einvp_2_9/a_36_74#
+ osc_core_1/sky130_fd_sc_hs__einvp_4_17/a_27_368# osc_core_1/sky130_fd_sc_hs__nand2_4_131/a_27_74#
+ osc_core_1/sky130_fd_sc_hs__and4_2_5/a_335_74# osc_core_1/sky130_fd_sc_hs__nand2_1_1/Y
+ osc_core_1/sky130_fd_sc_hs__clkbuf_4_5/A osc_core_1/sky130_fd_sc_hs__nand2_4_133/Y
+ osc_core_1/sky130_fd_sc_hs__nand2_8_35/a_27_74# osc_core_1/sky130_fd_sc_hs__nand2_2_29/Y
+ osc_core_1/sky130_fd_sc_hs__dlygate4sd2_1_1/a_405_138# osc_core_1/sky130_fd_sc_hs__nand2_2_63/a_27_74#
+ osc_core_1/sky130_fd_sc_hs__a21oi_1_28/a_117_74# osc_core_1/sky130_fd_sc_hs__einvp_4_5/a_27_74#
+ osc_core_1/sky130_fd_sc_hs__nand2_4_57/a_27_74# osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_79/a_289_74#
+ osc_core_1/sky130_fd_sc_hs__nand2_4_63/Y osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_9/a_405_138#
+ osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_15/a_289_74# osc_core_1/sky130_fd_sc_hs__nand2_2_97/Y
+ osc_core_1/sky130_fd_sc_hs__nand2_2_103/a_27_74# osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_62/a_405_138#
+ osc_core_1/sky130_fd_sc_hs__nand2_2_12/Y osc_core_1/sky130_fd_sc_hs__einvp_2_13/a_36_74#
+ osc_core_1/sky130_fd_sc_hs__dfrtp_4_1/a_1678_395# osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_56/a_28_74#
+ osc_core_1/sky130_fd_sc_hs__bufbuf_8_1/a_334_368# osc_core_1/sky130_fd_sc_hs__nand2_2_17/a_27_74#
+ osc_core_1/sky130_fd_sc_hs__nand2_2_89/a_27_74# osc_core_1/sky130_fd_sc_hs__nand2_4_111/a_27_74#
+ osc_core_1/sky130_fd_sc_hs__a21oi_1_47/a_29_368# osc_core_1/sky130_fd_sc_hs__nand2_4_127/Y
+ osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_1/a_289_74# osc_core_1/sky130_fd_sc_hs__nand2_4_93/Y
+ osc_core_1/sky130_fd_sc_hs__einvp_8_3/a_802_323# osc_core_1/sky130_fd_sc_hs__dfrtp_4_1/a_834_355#
+ osc_core_1/sky130_fd_sc_hs__einvp_2_3/a_263_323# osc_core_1/sky130_fd_sc_hs__einvp_4_1/a_473_323#
+ osc_core_1/sky130_fd_sc_hs__nand2_4_97/a_27_74# osc_core_1/sky130_fd_sc_hs__nand2_2_42/Y
+ osc_core_1/sky130_fd_sc_hs__nand2_4_125/a_27_74# osc_core_1/sky130_fd_sc_hs__nand2_4_3/a_27_74#
+ osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_79/a_28_74# osc_core_1/sky130_fd_sc_hs__einvp_8_17/a_802_323#
+ osc_core_1/sky130_fd_sc_hs__a21oi_1_11/a_117_74# osc_core_1/sky130_fd_sc_hs__and4_2_5/A
+ osc_core_1/sky130_fd_sc_hs__einvp_2_11/a_27_368# osc_core_1/sky130_fd_sc_hs__clkbuf_2_15/a_43_192#
+ osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_63/a_289_74# osc_core_1/sky130_fd_sc_hs__dfrtp_4_1/a_812_138#
+ osc_core_1/sky130_fd_sc_hs__einvp_8_7/a_27_74# osc_core_1/sky130_fd_sc_hs__nand2_4_157/Y
+ osc_core_1/sky130_fd_sc_hs__nand2_4_19/Y osc_core_1/sky130_fd_sc_hs__nand2_8_29/a_27_74#
+ osc_core_1/sky130_fd_sc_hs__nand2_2_57/a_27_74# osc_core_1/sky130_fd_sc_hs__nand3_4_1/a_27_82#
+ osc_core_1/sky130_fd_sc_hs__nand2_2_71/Y osc_core_1/sky130_fd_sc_hs__nand2_4_149/a_27_74#
+ osc_core_1/sky130_fd_sc_hs__nand2_4_119/Y osc_core_1/sky130_fd_sc_hs__nand2_4_85/Y
+ osc_core_1/sky130_fd_sc_hs__clkbuf_2_3/a_43_192# osc_core_1/sky130_fd_sc_hs__einvp_1_7/a_310_392#
+ osc_core_1/sky130_fd_sc_hs__einvp_4_3/a_27_368# osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_41/a_405_138#
+ osc_core_1/sky130_fd_sc_hs__dfrtp_4_3/a_1350_392# osc_core_1/sky130_fd_sc_hs__nand2_4_49/Y
+ osc_core_1/sky130_fd_sc_hs__einvp_4_19/a_473_323# osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_49/a_28_74#
+ osc_core_1/sky130_fd_sc_hs__a21oi_1_15/a_117_74# osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_33/a_289_74#
+ osc_core_1/sky130_fd_sc_hs__nand2_4_81/a_27_74# osc_core_1/sky130_fd_sc_hs__nand2_4_149/Y
+ osc_core_1/sky130_fd_sc_hs__einvp_4_17/a_27_74# osc_core_1/sky130_fd_sc_hs__nand2_8_5/a_27_74#
+ osc_core_1/sky130_fd_sc_hs__nand2_4_1/Y osc_core_1/sky130_fd_sc_hs__nand2_4_31/Y
+ osc_core_1/sky130_fd_sc_hs__einvp_1_11/a_310_392# osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_31/a_405_138#
+ osc_core_1/sky130_fd_sc_hs__nand2_4_79/Y osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_9/a_289_74#
+ osc_core_1/sky130_fd_sc_hs__clkbuf_2_7/a_43_192# osc_core_1/sky130_fd_sc_hs__a21oi_1_32/a_29_368#
+ osc_core_1/sky130_fd_sc_hs__nand2_2_42/a_27_74# osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_9/a_28_74#
+ osc_core_1/sky130_fd_sc_hs__nand2_2_27/Y osc_core_1/sky130_fd_sc_hs__nand2_4_133/a_27_74#
+ osc_core_1/sky130_fd_sc_hs__nand2_1_7/B osc_core_1/sky130_fd_sc_hs__nand2_4_60/Y
+ osc_core_1/sky130_fd_sc_hs__a21oi_1_19/a_117_74# osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_37/a_289_74#
+ osc_core_1/sky130_fd_sc_hs__dfrtp_4_1/a_1350_392# osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_33/a_28_74#
+ osc_core_1/sky130_fd_sc_hs__nand2_2_57/Y osc_core_1/sky130_fd_sc_hs__nand2_4_125/Y
+ osc_core_1/sky130_fd_sc_hs__nand2_4_91/Y osc_core_1/sky130_fd_sc_hs__a21oi_1_37/a_29_368#
+ osc_core_1/sky130_fd_sc_hs__nand2_2_83/a_27_74# osc_core_1/sky130_fd_sc_hs__nand2_4_75/a_27_74#
+ osc_core_1/sky130_fd_sc_hs__einvp_8_2/a_802_323# osc_core_1/sky130_fd_sc_hs__einvp_2_17/a_36_74#
+ osc_core_1/sky130_fd_sc_hs__nand2_4_102/a_27_74# osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_11/a_405_138#
+ osc_core_1/sky130_fd_sc_hs__einvp_1_11/a_318_74# osc_core_1/sky130_fd_sc_hs__nand2_2_88/Y
+ osc_core_1/sky130_fd_sc_hs__einvp_2_7/a_27_368# osc_core_1/sky130_fd_sc_hs__and2_2_1/a_31_74#
+ osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_51/a_289_74# osc_core_1/sky130_fd_sc_hs__nand2_4_17/Y
+ osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_74/a_28_74# osc_core_1/sky130_fd_sc_hs__nand2_4_155/Y
+ osc_core_1/sky130_fd_sc_hs__nand2_2_35/a_27_74# osc_core_1/sky130_fd_sc_hs__nand2_4_29/a_27_74#
+ osc_core_1/sky130_fd_sc_hs__einvp_8_2/a_27_74# osc_core_1/sky130_fd_sc_hs__nand2_2_103/Y
+ osc_core_1/sky130_fd_sc_hs__nand2_8_21/a_27_74# osc_core_1/sky130_fd_sc_hs__nand2_4_117/Y
+ osc_core_1/sky130_fd_sc_hs__nand2_2_1/Y osc_core_1/sky130_fd_sc_hs__nand2_4_43/a_27_74#
+ osc_core_1/sky130_fd_sc_hs__nand2_4_143/a_27_74# osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_27/a_28_74#
+ osc_core_1/sky130_fd_sc_hs__nand2_4_47/Y osc_core_1/sky130_fd_sc_hs__nand2_2_59/a_27_74#
+ osc_core_1/sky130_fd_sc_hs__einvp_1_15/a_318_74# osc_core_1/sky130_fd_sc_hs__a21oi_1_1/a_29_368#
+ osc_core_1/sky130_fd_sc_hs__nand2_2_79/Y osc_core_1/sky130_fd_sc_hs__nand2_8_47/a_27_74#
+ osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_57/a_289_74# osc_core_1/sky130_fd_sc_hs__bufbuf_8_1/a_27_112#
+ osc_core_1/sky130_fd_sc_hs__nand2_4_147/Y osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_23/a_289_74#
+ osc_core_1/sky130_fd_sc_hs__nand2_4_69/a_27_74# osc_core_1/sky130_fd_sc_hs__nand2_2_61/Y
+ osc_core_1/sky130_fd_sc_hs__nand2_4_77/Y osc_core_1/sky130_fd_sc_hs__dfrtp_4_1/a_124_78#
+ osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_79/a_405_138# osc_core_1/sky130_fd_sc_hs__nand2_4_13/a_27_74#
+ osc_core_1/sky130_fd_sc_hs__nand2_2_25/Y osc_core_1/sky130_fd_sc_hs__nand2_1_1/a_117_74#
+ osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_68/a_28_74# osc_core_1/sky130_fd_sc_hs__a21oi_1_23/a_29_368#
+ osc_core_1/sky130_fd_sc_hs__nand2_2_29/a_27_74# osc_core_1/sky130_fd_sc_hs__einvp_1_19/a_318_74#
+ osc_core_1/sky130_fd_sc_hs__a21oi_1_5/a_29_368# osc_core_1/sky130_fd_sc_hs__dfrtp_4_3/a_1647_81#
+ osc_core
Xsky130_fd_sc_hs__nand2_1_3 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__or2b_4_3/A sky130_fd_sc_hs__or4_2_1/D
+ sky130_fd_sc_hs__nor2_4_3/Y sky130_fd_sc_hs__nand2_1_3/a_117_74# sky130_fd_sc_hs__nand2_1
Xsky130_fd_sc_hs__einvp_2_140 DVSS: DVDD: DVDD: DVSS: dout_p sky130_fd_sc_hs__einvp_2_99/A
+ sky130_fd_sc_hs__dlrtp_1_143/Q sky130_fd_sc_hs__einvp_2_141/a_263_323# sky130_fd_sc_hs__einvp_2_141/a_36_74#
+ sky130_fd_sc_hs__einvp_2_141/a_27_368# sky130_fd_sc_hs__einvp_2
Xsky130_fd_sc_hs__einvp_2_151 DVSS: DVDD: DVDD: DVSS: dout_p sky130_fd_sc_hs__einvp_2_99/A
+ sky130_fd_sc_hs__buf_2_155/X sky130_fd_sc_hs__einvp_2_151/a_263_323# sky130_fd_sc_hs__einvp_2_151/a_36_74#
+ sky130_fd_sc_hs__einvp_2_151/a_27_368# sky130_fd_sc_hs__einvp_2
Xsky130_fd_sc_hs__clkbuf_16_12 DVSS: DVDD: DVDD: DVSS: osc_core_1/pi1_l[1] sky130_fd_sc_hs__clkbuf_4_19/X
+ sky130_fd_sc_hs__clkbuf_16_13/a_114_74# sky130_fd_sc_hs__clkbuf_16
Xsky130_fd_sc_hs__clkbuf_16_23 DVSS: DVDD: DVDD: DVSS: osc_core_1/pi1_l[0] sky130_fd_sc_hs__clkbuf_8_5/X
+ sky130_fd_sc_hs__clkbuf_16_23/a_114_74# sky130_fd_sc_hs__clkbuf_16
Xsky130_fd_sc_hs__clkbuf_16_34 DVSS: DVDD: DVDD: DVSS: osc_core_1/pi3_l[1] sky130_fd_sc_hs__clkbuf_8_9/X
+ sky130_fd_sc_hs__clkbuf_16_35/a_114_74# sky130_fd_sc_hs__clkbuf_16
Xsky130_fd_sc_hs__clkbuf_16_45 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__dlrtp_1_9/GATE
+ sky130_fd_sc_hs__clkbuf_2_3/A sky130_fd_sc_hs__clkbuf_16_45/a_114_74# sky130_fd_sc_hs__clkbuf_16
Xsky130_fd_sc_hs__clkbuf_16_56 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__buf_2_3/A
+ sky130_fd_sc_hs__einvp_8_3/Z sky130_fd_sc_hs__clkbuf_16_57/a_114_74# sky130_fd_sc_hs__clkbuf_16
Xsky130_fd_sc_hs__clkbuf_16_67 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__nand2_2_9/B
+ sky130_fd_sc_hs__or2b_2_5/A sky130_fd_sc_hs__clkbuf_16_67/a_114_74# sky130_fd_sc_hs__clkbuf_16
Xsky130_fd_sc_hs__clkbuf_16_78 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__nor4_2_1/B
+ sky130_fd_sc_hs__clkbuf_8_81/X sky130_fd_sc_hs__clkbuf_16_79/a_114_74# sky130_fd_sc_hs__clkbuf_16
Xsky130_fd_sc_hs__clkbuf_16_89 DVSS: DVDD: DVDD: DVSS: qr_4t1_mux_top_1/clk_IB qr_4t1_mux_top_3/clk_IB
+ sky130_fd_sc_hs__clkbuf_16_89/a_114_74# sky130_fd_sc_hs__clkbuf_16
Xsky130_fd_sc_hs__clkbuf_16_100 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__clkbuf_8_71/A
+ sky130_fd_sc_hs__clkbuf_8_95/X sky130_fd_sc_hs__clkbuf_16_101/a_114_74# sky130_fd_sc_hs__clkbuf_16
Xsky130_fd_sc_hs__clkbuf_16_111 DVSS: DVDD: DVDD: DVSS: prbs_generator_syn_31/rst
+ prbs_generator_syn_27/rst sky130_fd_sc_hs__clkbuf_16_111/a_114_74# sky130_fd_sc_hs__clkbuf_16
Xsky130_fd_sc_hs__clkbuf_16_122 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__clkbuf_8_59/A
+ sky130_fd_sc_hs__clkbuf_8_99/X sky130_fd_sc_hs__clkbuf_16_123/a_114_74# sky130_fd_sc_hs__clkbuf_16
Xsky130_fd_sc_hs__clkbuf_16_133 DVSS: DVDD: DVDD: DVSS: osc_core_1/pi5_l[0] pi5_con[0]
+ sky130_fd_sc_hs__clkbuf_16_133/a_114_74# sky130_fd_sc_hs__clkbuf_16
Xsky130_fd_sc_hs__nand2_2_19 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__buf_8_3/A sky130_fd_sc_hs__nor2_4_1/B
+ sky130_fd_sc_hs__or2b_2_1/A sky130_fd_sc_hs__nand2_2_19/a_27_74# sky130_fd_sc_hs__nand2_2
Xprbs_generator_syn_8 prbs_generator_syn_9/clk prbs_generator_syn_9/rst prbs_generator_syn_9/cke
+ sky130_fd_sc_hs__conb_1_85/LO sky130_fd_sc_hs__conb_1_85/LO sky130_fd_sc_hs__conb_1_85/HI
+ sky130_fd_sc_hs__conb_1_85/HI sky130_fd_sc_hs__conb_1_85/HI prbs_generator_syn_11/eqn[9]
+ sky130_fd_sc_hs__conb_1_85/LO sky130_fd_sc_hs__conb_1_85/HI sky130_fd_sc_hs__conb_1_85/HI
+ sky130_fd_sc_hs__conb_1_85/HI sky130_fd_sc_hs__conb_1_85/HI prbs_generator_syn_9/cke
+ prbs_generator_syn_9/cke prbs_generator_syn_9/eqn[31] prbs_generator_syn_9/cke prbs_generator_syn_9/cke
+ prbs_generator_syn_9/cke prbs_generator_syn_9/cke prbs_generator_syn_9/eqn[1] prbs_generator_syn_9/eqn[1]
+ prbs_generator_syn_9/eqn[1] prbs_generator_syn_9/eqn[1] prbs_generator_syn_9/eqn[1]
+ prbs_generator_syn_9/eqn[2] sky130_fd_sc_hs__conb_1_83/LO sky130_fd_sc_hs__conb_1_83/HI
+ sky130_fd_sc_hs__conb_1_83/LO sky130_fd_sc_hs__conb_1_83/HI sky130_fd_sc_hs__conb_1_83/HI
+ sky130_fd_sc_hs__conb_1_83/LO sky130_fd_sc_hs__conb_1_83/LO sky130_fd_sc_hs__conb_1_83/HI
+ prbs_generator_syn_9/eqn[31] prbs_generator_syn_9/eqn[30] prbs_generator_syn_9/eqn[30]
+ prbs_generator_syn_9/eqn[28] prbs_generator_syn_9/eqn[28] prbs_generator_syn_9/eqn[28]
+ prbs_generator_syn_9/eqn[28] prbs_generator_syn_9/eqn[28] prbs_generator_syn_9/eqn[28]
+ prbs_generator_syn_9/eqn[22] prbs_generator_syn_9/eqn[22] prbs_generator_syn_9/eqn[20]
+ prbs_generator_syn_9/eqn[22] prbs_generator_syn_9/eqn[22] prbs_generator_syn_9/eqn[22]
+ prbs_generator_syn_9/eqn[16] prbs_generator_syn_9/eqn[16] prbs_generator_syn_9/eqn[16]
+ prbs_generator_syn_3/eqn[4] prbs_generator_syn_9/eqn[16] prbs_generator_syn_9/eqn[16]
+ prbs_generator_syn_9/eqn[16] prbs_generator_syn_9/eqn[9] prbs_generator_syn_9/eqn[9]
+ prbs_generator_syn_9/eqn[9] prbs_generator_syn_9/eqn[9] prbs_generator_syn_9/eqn[9]
+ prbs_generator_syn_9/eqn[9] prbs_generator_syn_9/eqn[9] prbs_generator_syn_9/eqn[2]
+ prbs_generator_syn_9/eqn[1] prbs_generator_syn_9/eqn[2] prbs_generator_syn_9/inj_err
+ prbs_generator_syn_9/eqn[31] prbs_generator_syn_9/eqn[31] prbs_generator_syn_9/out
+ DVSS: DVDD: prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_1/a_293_74# prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_15/X
+ prbs_generator_syn_9/sky130_fd_sc_hs__nand2_1_35/B prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_51/Y
+ prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_9/A prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_9/CLK
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_47/a_27_74# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_37/a_1226_296#
+ prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_3/B prbs_generator_syn_9/sky130_fd_sc_hs__nor2b_1_7/a_27_112#
+ prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_29/B prbs_generator_syn_9/sky130_fd_sc_hs__sdlclkp_2_1/a_580_74#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_1/a_1141_508# prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_5/Y
+ prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_41/a_230_79# prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_61/a_138_385#
+ prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_43/a_132_392# prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_3/a_222_392#
+ prbs_generator_syn_9/sky130_fd_sc_hs__nor2b_1_9/a_27_112# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_61/a_27_74#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_35/a_206_368# prbs_generator_syn_9/sky130_fd_sc_hs__nand2_2_3/Y
+ prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_25/B prbs_generator_syn_9/sky130_fd_sc_hs__nand2_1_11/a_117_74#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_67/a_651_503# prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_45/X
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_39/a_696_458# prbs_generator_syn_9/sky130_fd_sc_hs__sdlclkp_2_1/a_1198_74#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_45/a_1034_424# prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_17/a_222_392#
+ prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_55/a_222_392# prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_53/Y
+ prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_35/A prbs_generator_syn_9/m3_13600_1651#
+ prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_59/a_52_123# prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_5/a_293_74#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_35/a_1226_296# prbs_generator_syn_9/sky130_fd_sc_hs__nand2_1_51/B
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_5/a_651_503# prbs_generator_syn_9/sky130_fd_sc_hs__nand2_1_21/B
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_8/a_27_74# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_15/a_27_74#
+ prbs_generator_syn_9/sky130_fd_sc_hs__and2b_2_1/X prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_13/X
+ prbs_generator_syn_9/sky130_fd_sc_hs__nand2_2_3/a_27_74# prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_50/a_138_385#
+ prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_33/a_132_392# prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_1/a_376_368#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_25/a_206_368# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_35/a_437_503#
+ prbs_generator_syn_9/sky130_fd_sc_hs__sdlclkp_2_1/a_708_451# prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_45/a_230_79#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_29/a_696_458# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_32/a_27_74#
+ prbs_generator_syn_9/sky130_fd_sc_hs__nor2b_1_4/Y prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_59/a_293_74#
+ prbs_generator_syn_9/sky130_fd_sc_hs__nand2_1_47/a_117_74# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_73/a_735_102#
+ prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_21/a_112_119# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_23/a_1141_508#
+ prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_25/a_293_74# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_7/Q
+ prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_3/a_112_119# prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_35/B
+ prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_51/X prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_53/a_1178_124#
+ prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_23/a_132_392# prbs_generator_syn_9/sky130_fd_sc_hs__nand2_1_3/B
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_15/a_206_368# prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_63/a_132_392#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_55/a_27_74# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_25/a_437_503#
+ prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_41/a_52_123# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_47/a_651_503#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_73/a_1141_508# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_19/a_696_458#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_57/a_696_458# prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_7/X
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_43/a_1034_424# prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_55/A
+ prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_11/a_112_119# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_21/a_1141_508#
+ prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_35/a_222_392# prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_49/a_230_79#
+ prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_67/Y prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_71/a_27_74#
+ prbs_generator_syn_9/sky130_fd_sc_hs__nand2_1_33/B prbs_generator_syn_9/sky130_fd_sc_hs__conb_1_1/LO
+ prbs_generator_syn_9/sky130_fd_sc_hs__nand2_1_19/a_117_74# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_51/a_1178_124#
+ prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_33/X prbs_generator_syn_9/sky130_fd_sc_hs__nand2_1_29/B
+ prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_41/Y prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_53/a_132_392#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_45/a_206_368# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_15/a_437_503#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_37/a_651_503# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_39/a_544_485#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_53/a_735_102# prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_45/a_52_123#
+ prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_1/B prbs_generator_syn_9/sky130_fd_sc_hs__nand2_2_3/B
+ prbs_generator_syn_9/sky130_fd_sc_hs__clkbuf_16_1/A prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_21/X
+ prbs_generator_syn_9/sky130_fd_sc_hs__nand2_1_25/B prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_39/a_376_368#
+ prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_63/X prbs_generator_syn_9/m3_13600_3481#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_69/a_1178_124# prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_21/a_138_385#
+ prbs_generator_syn_9/sky130_fd_sc_hs__nor2b_1_8/Y prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_19/a_1178_124#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_49/a_27_74# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_45/a_437_503#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_27/a_651_503# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_71/a_1141_508#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_65/a_651_503# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_29/a_544_485#
+ prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_3/a_138_385# prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_55/X
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_43/a_735_102# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_41/a_1034_424#
+ prbs_generator_syn_9/sky130_fd_sc_hs__nand2_1_9/B prbs_generator_syn_9/sky130_fd_sc_hs__nor2b_1_9/Y
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_59/a_1034_424# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_39/a_1141_508#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_33/a_1226_296# prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_49/a_52_123#
+ prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_47/Y prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_43/Y
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_4/a_651_503# prbs_generator_syn_9/sky130_fd_sc_hs__nand2_1_49/B
+ prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_19/A prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_11/a_138_385#
+ prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_5/X prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_63/a_206_368#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_17/a_651_503# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_19/a_544_485#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_55/a_651_503# prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_9/Y
+ prbs_generator_syn_9/sky130_fd_sc_hs__nand2_1_17/B prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_57/a_544_485#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_67/a_696_458# prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_35/X
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_19/a_27_74# prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_45/a_222_392#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_32/a_1226_296# prbs_generator_syn_9/sky130_fd_sc_hs__nand2_1_43/B
+ prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_25/A prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_1/a_206_368#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_49/a_1226_296# prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_1/a_112_119#
+ prbs_generator_syn_9/sky130_fd_sc_hs__or2_1_1/X prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_59/a_376_368#
+ prbs_generator_syn_9/sky130_fd_sc_hs__nand2_1_19/B prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_5/a_696_458#
+ prbs_generator_syn_9/sky130_fd_sc_hs__nor2b_1_1/Y prbs_generator_syn_9/sky130_fd_sc_hs__nor2b_1_5/a_278_368#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_17/a_1178_124# prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_39/X
+ prbs_generator_syn_9/m3_13600_5433# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_63/a_437_503#
+ prbs_generator_syn_9/sky130_fd_sc_hs__nand2_2_5/B prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_23/a_735_102#
+ prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_53/A prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_61/a_735_102#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_57/a_1034_424# prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_63/B
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_37/a_1141_508# prbs_generator_syn_9/sky130_fd_sc_hs__nand2_1_47/B
+ prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_29/X prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_65/Y
+ prbs_generator_syn_9/m3_13600_4701# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_1/a_437_503#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_67/a_1178_124# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_9/a_735_102#
+ prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_13/a_132_392# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_15/a_1178_124#
+ prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_15/A prbs_generator_syn_9/sky130_fd_sc_hs__nand2_1_1/B
+ prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_43/B prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_35/a_651_503#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_8/D prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_29/A
+ prbs_generator_syn_9/sky130_fd_sc_hs__nand2_1_7/B prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_13/a_735_102#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_47/a_696_458# prbs_generator_syn_9/sky130_fd_sc_hs__nand2_1_31/B
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_51/a_735_102# prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_59/X
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_35/a_1141_508# prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_25/a_222_392#
+ prbs_generator_syn_9/sky130_fd_sc_hs__sdlclkp_2_1/a_288_48# prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_55/B
+ prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_17/B prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_43/A
+ prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_7/A prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_65/a_1178_124#
+ prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_59/Y prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_41/X
+ prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_21/a_230_79# prbs_generator_syn_9/sky130_fd_sc_hs__nand2_1_57/a_117_74#
+ prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_1/a_222_392# prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_19/B
+ prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_35/a_293_74# prbs_generator_syn_9/sky130_fd_sc_hs__nand2_1_23/a_117_74#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_73/a_206_368# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_25/a_651_503#
+ prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_1/a_138_385# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_37/a_696_458#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_67/a_544_485# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_43/a_27_74#
+ prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_9/X prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_55/a_1034_424#
+ prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_39/a_112_119# prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_15/a_222_392#
+ prbs_generator_syn_9/sky130_fd_sc_hs__conb_1_1/HI prbs_generator_syn_9/sky130_fd_sc_hs__nand2_1_23/B
+ prbs_generator_syn_9/sky130_fd_sc_hs__nand2_1_53/B prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_9/a_1178_124#
+ prbs_generator_syn_9/sky130_fd_sc_hs__nor2b_1_4/A prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_47/a_1226_296#
+ prbs_generator_syn_9/m3_13600_11045# prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_17/X
+ prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_29/a_376_368# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_5/a_544_485#
+ prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_3/X prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_31/a_132_392#
+ prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_61/A prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_15/a_651_503#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_73/a_437_503# prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_25/a_230_79#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_27/a_696_458# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_65/a_696_458#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_33/a_735_102# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_71/a_735_102#
+ prbs_generator_syn_9/m3_13600_7263# prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_43/a_222_392#
+ prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_50/Y prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_8/a_1178_124#
+ prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_53/B prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_19/a_376_368#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_63/a_1178_124# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_4/a_696_458#
+ prbs_generator_syn_9/sky130_fd_sc_hs__nor2b_1_4/a_278_368# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_13/a_1178_124#
+ prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_61/a_132_392# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_53/a_206_368#
+ prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_21/a_52_123# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_45/a_651_503#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_17/a_696_458# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_47/a_544_485#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_55/a_696_458# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_21/a_735_102#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_37/a_27_74# prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_61/B
+ prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_61/X prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_59/a_112_119#
+ prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_31/A prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_33/a_222_392#
+ prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_29/a_230_79# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_45/a_1226_296#
+ prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_9/a_132_392# prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_5/A
+ prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_57/Y prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_31/X
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_51/a_27_74# prbs_generator_syn_9/sky130_fd_sc_hs__nor2b_1_8/a_27_112#
+ prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_47/a_376_368# prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_53/a_293_74#
+ prbs_generator_syn_9/sky130_fd_sc_hs__nand2_1_43/a_117_74# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_8/a_735_102#
+ prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_21/a_293_74# prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_39/a_138_385#
+ prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_63/Y prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_51/a_132_392#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_43/a_206_368# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_53/a_437_503#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_37/a_544_485# prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_57/X
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_53/a_1034_424# prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_25/a_52_123#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_33/a_1141_508# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_63/Q
+ prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_23/a_222_392# prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_63/a_222_392#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_7/a_1178_124# prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_53/X
+ prbs_generator_syn_9/sky130_fd_sc_hs__nand2_2_5/Y prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_61/a_1178_124#
+ prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_1/a_230_79# prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_43/a_230_79#
+ prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_11/a_230_79# prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_41/a_132_392#
+ prbs_generator_syn_9/sky130_fd_sc_hs__nand2_1_13/a_117_74# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_43/a_437_503#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_27/a_544_485# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_63/a_651_503#
+ prbs_generator_syn_9/sky130_fd_sc_hs__nand2_1_7/a_117_74# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_35/a_696_458#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_65/a_544_485# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_51/a_1034_424#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_41/a_735_102# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_32/a_1141_508#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_49/a_1141_508# prbs_generator_syn_9/sky130_fd_sc_hs__nand2_1_55/B
+ prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_53/a_222_392# prbs_generator_syn_9/sky130_fd_sc_hs__sdlclkp_2_1/a_114_112#
+ prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_9/a_293_74# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_43/a_1226_296#
+ prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_29/a_52_123# prbs_generator_syn_9/sky130_fd_sc_hs__nand2_1_37/B
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_1/a_651_503# prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_27/a_376_368#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_4/a_544_485# prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_67/a_376_368#
+ prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_27/X prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_1/X
+ prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_59/a_138_385# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_29/a_1178_124#
+ prbs_generator_syn_9/m3_13600_2871# prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_5/a_230_79#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_23/a_206_368# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_61/a_206_368#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_17/a_544_485# prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_15/a_230_79#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_25/a_696_458# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_55/a_544_485#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_32/a_735_102# prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_29/a_293_74#
+ prbs_generator_syn_9/sky130_fd_sc_hs__nand2_1_17/a_117_74# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_69/a_1034_424#
+ prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_29/a_112_119# prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_37/X
+ prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_31/B prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_19/a_1034_424#
+ prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_33/A prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_9/a_206_368#
+ prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_57/a_376_368# prbs_generator_syn_9/sky130_fd_sc_hs__sdlclkp_2_1/a_706_317#
+ prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_11/B prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_1/a_52_123#
+ prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_39/B prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_21/a_132_392#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_13/a_206_368# prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_43/a_52_123#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_51/a_206_368# prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_47/X
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_23/a_437_503# prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_11/a_52_123#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_61/a_437_503# prbs_generator_syn_9/sky130_fd_sc_hs__nor2b_1_7/Y
+ prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_51/A prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_15/a_696_458#
+ prbs_generator_syn_9/sky130_fd_sc_hs__nor2b_1_5/Y prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_9/a_230_79#
+ prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_25/X prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_19/a_112_119#
+ prbs_generator_syn_9/sky130_fd_sc_hs__nand2_1_45/B prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_5/a_1178_124#
+ prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_19/a_230_79# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_41/a_1226_296#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_59/a_1226_296# prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_63/a_230_79#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_51/Q prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_7/a_132_392#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_9/a_437_503# prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_46/a_376_368#
+ prbs_generator_syn_9/sky130_fd_sc_hs__nand2_1_33/a_117_74# prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_11/a_293_74#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_27/a_1178_124# prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_11/a_132_392#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_13/a_437_503# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_51/a_437_503#
+ prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_5/a_52_123# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_35/a_544_485#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_73/a_651_503# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_45/a_696_458#
+ prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_15/a_52_123# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_47/a_1141_508#
+ prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_47/a_112_119# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_4/a_1178_124#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_17/a_1034_424# prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_23/B
+ prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_37/a_376_368# prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_15/B
+ prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_7/Y prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_29/a_138_385#
+ prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_33/a_230_79# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_25/a_1178_124#
+ prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_47/a_293_74# prbs_generator_syn_9/sky130_fd_sc_hs__nand2_1_37/a_117_74#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_33/a_206_368# prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_15/a_293_74#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_71/a_206_368# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_25/a_544_485#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_67/a_1034_424# prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_13/a_222_392#
+ prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_9/a_52_123# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_15/a_1034_424#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_57/a_1226_296# prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_19/a_52_123#
+ prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_23/X prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_63/a_52_123#
+ prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_19/a_138_385# prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_9/a_376_368#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_21/a_206_368# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_33/a_437_503#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_71/a_437_503# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_53/a_651_503#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_15/a_544_485# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_63/a_696_458#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_65/a_1034_424# prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_19/a_293_74#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_45/a_1141_508# prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_27/a_112_119#
+ prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_67/a_112_119# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_1/a_1178_124#
+ prbs_generator_syn_9/sky130_fd_sc_hs__conb_1_1/a_21_290# prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_63/a_293_74#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_8/a_206_368# prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_17/a_376_368#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_63/a_27_74# prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_21/A
+ prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_55/a_376_368# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_1/a_696_458#
+ prbs_generator_syn_9/sky130_fd_sc_hs__nor2b_1_1/a_278_368# prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_47/a_138_385#
+ prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_33/a_52_123# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_9/a_1034_424#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_21/a_437_503# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_1/a_27_74#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_43/a_651_503# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_1/Q
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_45/a_544_485# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_69/a_735_102#
+ prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_57/a_112_119# prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_31/a_222_392#
+ prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_13/A prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_55/a_1226_296#
+ prbs_generator_syn_9/sky130_fd_sc_hs__nand2_2_5/a_27_74# prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_53/a_230_79#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_8/a_437_503# prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_67/a_293_74#
+ prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_33/a_293_74# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_7/a_735_102#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_23/a_1178_124# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_41/a_206_368#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_8/a_1034_424# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_63/a_1034_424#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_59/a_735_102# prbs_generator_syn_9/sky130_fd_sc_hs__nand2_1_5/B
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_43/a_1141_508# prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_46/a_112_119#
+ prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_61/a_222_392# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_13/a_1034_424#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_73/a_1178_124# prbs_generator_syn_9/sky130_fd_sc_hs__nand2_1_27/B
+ prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_13/B prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_57/a_27_74#
+ prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_57/a_230_79# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_21/a_1178_124#
+ prbs_generator_syn_9/sky130_fd_sc_hs__nor2b_1_1/a_27_112# prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_27/a_138_385#
+ prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_23/a_230_79# prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_67/a_138_385#
+ prbs_generator_syn_9/sky130_fd_sc_hs__nand2_1_41/B prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_9/a_222_392#
+ prbs_generator_syn_9/sky130_fd_sc_hs__nand2_1_27/a_117_74# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_32/a_206_368#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_23/a_651_503# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_41/a_437_503#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_73/a_27_74# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_61/a_651_503#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_63/a_544_485# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_49/a_735_102#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_73/a_696_458# prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_37/a_112_119#
+ prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_51/a_222_392# prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_43/X
+ prbs_generator_syn_9/sky130_fd_sc_hs__nand2_2_1/B prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_9/a_651_503#
+ prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_53/a_52_123# prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_49/X
+ prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_25/a_376_368# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_1/a_544_485#
+ prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_65/a_376_368# prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_57/a_138_385#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_27/a_27_74# prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_39/a_132_392#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_7/a_1034_424# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_13/a_651_503#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_32/a_437_503# prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_27/a_230_79#
+ prbs_generator_syn_9/m3_13600_12265# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_51/a_651_503#
+ prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_59/B prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_47/A
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_61/a_1034_424# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_41/a_1141_508#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_59/a_1141_508# prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_41/a_222_392#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_53/a_1226_296# prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_3/A
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_71/a_1178_124# prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_9/a_112_119#
+ prbs_generator_syn_9/sky130_fd_sc_hs__nand2_1_3/a_117_74# prbs_generator_syn_9/m3_13600_8483#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_39/a_1178_124# prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_57/a_52_123#
+ prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_46/a_138_385# prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_23/a_52_123#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_67/a_27_74# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_53/a_696_458#
+ prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_17/a_112_119# prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_11/A
+ prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_55/a_112_119# prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_1/A
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_51/a_1226_296# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_29/a_1034_424#
+ prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_59/A prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_23/A
+ prbs_generator_syn_9/sky130_fd_sc_hs__nand2_1_39/B prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_5/a_27_74#
+ prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_57/a_293_74# prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_37/a_138_385#
+ prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_59/a_132_392# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_33/a_651_503#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_71/a_651_503# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_43/a_696_458#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_73/a_544_485# prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_27/a_52_123#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_57/a_1141_508# prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_21/a_222_392#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_35/a_27_74# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_69/a_1226_296#
+ prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_37/B prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_19/a_1226_296#
+ prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_35/a_376_368# prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_47/a_230_79#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_37/a_1178_124# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_5/a_1034_424#
+ prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_49/a_132_392# prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_7/a_222_392#
+ prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_27/a_293_74# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_21/a_651_503#
+ prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_9/a_138_385# prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_11/a_222_392#
+ prbs_generator_syn_9/m3_13600_14095# prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_50/A
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_27/a_1034_424# prbs_generator_syn_9/sky130_fd_sc_hs__nand2_1_13/B
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_8/a_651_503# prbs_generator_syn_9/m3_13600_9703#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_35/a_1178_124# prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_17/a_138_385#
+ prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_55/a_138_385# prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_7/a_230_79#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_4/a_1034_424# prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_7/a_376_368#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_69/a_206_368# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_23/a_696_458#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_53/a_544_485# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_39/a_735_102#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_61/a_696_458# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_55/a_1141_508#
+ prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_25/a_112_119# prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_65/a_112_119#
+ prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_43/a_293_74# prbs_generator_syn_9/sky130_fd_sc_hs__nand2_1_57/B
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_25/a_1034_424# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_7/a_206_368#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_17/a_1226_296# prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_15/a_376_368#
+ prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_53/a_376_368# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_9/a_696_458#
+ prbs_generator_syn_9/m3_13600_431# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_45/a_27_74#
+ prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_47/a_52_123# prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_29/a_132_392#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_59/a_206_368# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_69/a_437_503#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_41/a_651_503# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_43/a_544_485#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_13/a_696_458# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_29/a_735_102#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_51/a_696_458# prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_61/Y
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_67/a_1226_296# prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_5/a_132_392#
+ prbs_generator_syn_9/sky130_fd_sc_hs__and2b_2_1/a_198_48# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_7/a_437_503#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_15/a_1226_296# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_69/a_27_74#
+ prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_46/a_293_74# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_1/a_1034_424#
+ prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_19/a_132_392# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_49/a_206_368#
+ prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_7/a_52_123# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_59/a_437_503#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_32/a_651_503# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_7/a_27_74#
+ prbs_generator_syn_9/sky130_fd_sc_hs__nand2_2_1/a_27_74# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_19/a_735_102#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_57/a_735_102# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_65/a_1226_296#
+ prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_37/A prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_33/a_376_368#
+ prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_37/a_230_79# prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_25/a_138_385#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_39/a_27_74# prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_65/a_138_385#
+ prbs_generator_syn_9/sky130_fd_sc_hs__nor2b_1_9/a_278_368# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_49/a_437_503#
+ prbs_generator_syn_9/sky130_fd_sc_hs__and2b_2_1/a_505_74# prbs_generator_syn_9/sky130_fd_sc_hs__nand2_1_51/a_117_74#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_23/a_544_485# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_33/a_696_458#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_61/a_544_485# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_9/a_1226_296#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_53/a_1141_508# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_71/a_696_458#
+ prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_35/a_112_119# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_23/a_1034_424#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_9/a_544_485# prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_63/a_376_368#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_33/a_1178_124# prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_5/a_376_368#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_13/a_544_485# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_73/a_1034_424#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_21/a_696_458# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_51/a_544_485#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_8/a_1226_296# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_51/a_1141_508#
+ prbs_generator_syn_9/sky130_fd_sc_hs__nand2_1_55/a_117_74# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_21/a_1034_424#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_63/a_1226_296# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_23/a_27_74#
+ prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_7/a_112_119# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_13/a_1226_296#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_8/a_696_458# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_32/a_1178_124#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_49/a_1178_124# prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_37/a_52_123#
+ prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_27/a_132_392# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_71/Q
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_67/a_735_102# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_69/a_1141_508#
+ prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_15/a_112_119# prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_53/a_112_119#
+ prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_39/a_222_392# prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_55/a_230_79#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_19/a_1141_508# prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_37/a_293_74#
+ prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_43/a_376_368# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_5/a_735_102#
+ prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_35/a_138_385# prbs_generator_syn_9/sky130_fd_sc_hs__sdlclkp_2_1/a_114_424#
+ prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_57/a_132_392# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_71/a_1034_424#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_7/a_1226_296# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_33/a_544_485#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_41/a_696_458# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_71/a_544_485#
+ prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_21/B prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_61/a_1226_296#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_39/a_1034_424# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_17/a_27_74#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_9/a_27_74# prbs_generator_syn_9/sky130_fd_sc_hs__nor2b_1_5/a_27_112#
+ prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_47/a_132_392# prbs_generator_syn_9/sky130_fd_sc_hs__nor2b_1_8/a_278_368#
+ prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_9/B prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_39/a_206_368#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_33/a_27_74# prbs_generator_syn_9/sky130_fd_sc_hs__nand2_1_41/a_117_74#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_69/a_651_503# prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_51/a_293_74#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_21/a_544_485# prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_7/a_138_385#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_32/a_696_458# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_47/a_735_102#
+ prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_33/a_112_119# prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_59/a_222_392#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_17/a_1141_508# prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_55/a_52_123#
+ prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_3/a_293_74# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_7/a_651_503#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_29/a_1226_296# prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_23/a_376_368#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_8/a_544_485# prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_47/B
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_47/a_1178_124# prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_15/a_138_385#
+ prbs_generator_syn_9/sky130_fd_sc_hs__sdlclkp_2_1/a_1195_374# prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_53/a_138_385#
+ prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_37/a_132_392# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_29/a_206_368#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_39/a_437_503# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_59/a_651_503#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_37/a_735_102# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_67/a_1141_508#
+ prbs_generator_syn_9/sky130_fd_sc_hs__and2b_2_1/a_27_74# prbs_generator_syn_9/sky130_fd_sc_hs__conb_1_1/a_165_290#
+ prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_55/a_293_74# prbs_generator_syn_9/sky130_fd_sc_hs__nand2_1_45/a_117_74#
+ prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_63/a_112_119# prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_49/a_222_392#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_37/a_1034_424# prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_23/a_293_74#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_15/a_1141_508# prbs_generator_syn_9/sky130_fd_sc_hs__nand2_1_5/a_117_74#
+ prbs_generator_syn_9/m3_13600_13485# prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_5/a_112_119#
+ prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_13/a_376_368# prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_51/a_376_368#
+ prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_7/a_293_74# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_19/a_206_368#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_57/a_206_368# prbs_generator_syn_9/sky130_fd_sc_hs__sdlclkp_2_1/a_318_74#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_29/a_437_503# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_49/a_651_503#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_25/a_27_74# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_5/a_1226_296#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_41/a_544_485# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_27/a_735_102#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_65/a_1141_508# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_65/a_735_102#
+ prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_3/a_230_79# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_35/a_1034_424#
+ prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_13/a_230_79# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_41/a_27_74#
+ prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_3/a_132_392# prbs_generator_syn_9/sky130_fd_sc_hs__nand2_1_49/a_117_74#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_27/a_1226_296# prbs_generator_syn_9/sky130_fd_sc_hs__nand2_1_15/a_117_74#
+ prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_41/a_376_368# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_45/a_1178_124#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_4/a_735_102# prbs_generator_syn_9/sky130_fd_sc_hs__nand2_1_9/a_117_74#
+ prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_33/a_138_385# prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_17/a_132_392#
+ prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_55/a_132_392# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_9/a_1141_508#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_19/a_437_503# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_57/a_437_503#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_4/a_1226_296# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_32/a_544_485#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_17/a_735_102# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_55/a_735_102#
+ prbs_generator_syn_9/m3_13600_2261# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_65/a_27_74#
+ prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_29/a_222_392# prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_43/a_112_119#
+ prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_19/X prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_25/a_1226_296#
+ prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_31/a_376_368# prbs_generator_syn_9/sky130_fd_sc_hs__or2_1_1/a_63_368#
+ prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_17/a_230_79# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_4/a_27_74#
+ prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_61/a_230_79# prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_63/a_138_385#
+ prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_5/a_222_392# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_8/a_1141_508#
+ prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_41/a_293_74# prbs_generator_syn_9/sky130_fd_sc_hs__nand2_1_31/a_117_74#
+ prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_5/a_138_385# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_63/a_1141_508#
+ prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_19/a_222_392# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_13/a_1141_508#
+ prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_3/a_52_123# prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_13/a_52_123#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_43/a_1178_124# prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_61/a_376_368#
+ prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_35/a_132_392# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_67/a_206_368#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_1/a_1226_296# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_69/a_696_458#
+ prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_31/a_230_79# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_35/a_735_102#
+ prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_23/a_112_119# prbs_generator_syn_9/sky130_fd_sc_hs__nand2_1_35/a_117_74#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_59/a_27_74# prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_13/a_293_74#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_5/a_206_368# prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_50/a_376_368#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_7/a_696_458# prbs_generator_syn_9/sky130_fd_sc_hs__nor2b_1_7/a_278_368#
+ prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_17/a_52_123# prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_43/a_138_385#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_7/a_1141_508# prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_61/a_52_123#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_67/a_437_503# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_61/a_1141_508#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_25/a_735_102# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_59/a_696_458#
+ prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_13/a_112_119# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_33/a_1034_424#
+ prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_51/a_112_119# prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_35/a_230_79#
+ prbs_generator_syn_9/m3_13600_4091# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_23/a_1226_296#
+ prbs_generator_syn_9/sky130_fd_sc_hs__nand2_1_39/a_117_74# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_29/a_27_74#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_5/a_437_503# prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_17/a_293_74#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_41/a_1178_124# prbs_generator_syn_9/sky130_fd_sc_hs__or2_1_1/a_152_368#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_59/a_1178_124# prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_61/a_293_74#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_47/a_206_368# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_39/a_651_503#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_49/a_696_458# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_15/a_735_102#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_32/a_1034_424# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_73/a_1226_296#
+ prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_27/a_222_392# prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_41/a_112_119#
+ prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_31/a_52_123# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_49/a_1034_424#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_29/a_1141_508# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_21/a_1226_296#
+ prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_39/a_230_79# prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_23/a_138_385#
+ prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_51/a_230_79# prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_45/a_132_392#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_37/a_206_368# prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_65/a_293_74#
+ prbs_generator_syn_9/sky130_fd_sc_hs__nand2_1_53/a_117_74# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_47/a_437_503#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_29/a_651_503# prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_31/a_293_74#
+ prbs_generator_syn_9/sky130_fd_sc_hs__nand2_1_21/a_117_74# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_69/a_544_485#
+ prbs_generator_syn_9/sky130_fd_sc_hs__clkbuf_16_1/a_114_74# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_45/a_735_102#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_13/a_27_74# prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_31/a_112_119#
+ prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_57/a_222_392# prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_35/a_52_123#
+ prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_21/a_376_368# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_7/a_544_485#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_57/a_1178_124# prbs_generator_syn_9/m3_13600_6043#
+ prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_13/a_138_385# prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_51/a_138_385#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_5/a_1141_508# prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_3/a_376_368#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_27/a_206_368# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_65/a_206_368#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_37/a_437_503# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_19/a_651_503#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_57/a_651_503# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_59/a_544_485#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_71/a_1226_296# prbs_generator_syn_9/sky130_fd_sc_hs__nand2_1_25/a_117_74#
+ prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_61/a_112_119# prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_47/a_222_392#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_27/a_1141_508# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_53/a_27_74#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_4/a_206_368# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_39/a_1226_296#
+ prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_11/a_376_368# prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_39/a_52_123#
+ prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_41/a_138_385# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_4/a_1141_508#
+ prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_25/a_132_392# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_17/a_206_368#
+ prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_41/A prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_55/a_206_368#
+ prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_51/a_52_123# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_27/a_437_503#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_65/a_437_503# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_49/a_544_485#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_63/a_735_102# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_47/a_1034_424#
+ prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_50/a_112_119# prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_37/a_222_392#
+ prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_59/a_230_79# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_25/a_1141_508#
+ prbs_generator_syn_9/sky130_fd_sc_hs__nor2b_1_4/a_27_112# prbs_generator_syn_9/sky130_fd_sc_hs__sdlclkp_2_1/a_685_81#
+ prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_1/a_132_392# prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_39/a_293_74#
+ prbs_generator_syn_9/sky130_fd_sc_hs__nand2_1_29/a_117_74# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_4/a_437_503#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_55/a_1178_124# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_21/a_27_74#
+ prbs_generator_syn_9/m3_13600_12875# prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_50/a_293_74#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_1/a_735_102# prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_31/a_138_385#
+ prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_15/a_132_392# prbs_generator_syn_9/sky130_fd_sc_hs__nand2_1_1/a_117_74#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_17/a_437_503# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_55/a_437_503#
+ prbs_generator_syn
Xsky130_fd_sc_hs__clkbuf_4_100 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__clkbuf_4_109/X
+ fine_freq_track_1/fftl_en sky130_fd_sc_hs__clkbuf_4_101/a_83_270# sky130_fd_sc_hs__clkbuf_4
Xsky130_fd_sc_hs__clkbuf_4_111 DVSS: DVDD: DVDD: DVSS: inj_en osc_core_1/inj_en sky130_fd_sc_hs__clkbuf_4_111/a_83_270#
+ sky130_fd_sc_hs__clkbuf_4
Xsky130_fd_sc_hs__clkbuf_4_122 DVSS: DVDD: DVDD: DVSS: CTL_BUF_N[5] sky130_fd_sc_hs__clkbuf_4_123/X
+ sky130_fd_sc_hs__clkbuf_4_123/a_83_270# sky130_fd_sc_hs__clkbuf_4
Xsky130_fd_sc_hs__clkbuf_4_133 DVSS: DVDD: DVDD: DVSS: inj_error sky130_fd_sc_hs__clkbuf_8_91/A
+ sky130_fd_sc_hs__clkbuf_4_133/a_83_270# sky130_fd_sc_hs__clkbuf_4
Xsky130_fd_sc_hs__o21ai_2_2 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__inv_4_13/Y sky130_fd_sc_hs__o21ai_2_3/A2
+ sky130_fd_sc_hs__nand2_2_9/B sky130_fd_sc_hs__buf_2_41/A sky130_fd_sc_hs__o21ai_2_3/a_116_368#
+ sky130_fd_sc_hs__o21ai_2_3/a_27_74# sky130_fd_sc_hs__o21ai_2
Xsky130_fd_sc_hs__clkdlyinv5sd2_1_7 DVSS: DVDD: DVSS: DVDD: dout_n sky130_fd_sc_hs__and2_2_1/A
+ sky130_fd_sc_hs__clkdlyinv5sd2_1_7/a_28_74# sky130_fd_sc_hs__clkdlyinv5sd2_1_7/a_682_74#
+ sky130_fd_sc_hs__clkdlyinv5sd2_1_7/a_549_74# sky130_fd_sc_hs__clkdlyinv5sd2_1_7/a_288_74#
+ sky130_fd_sc_hs__clkdlyinv5sd2_1
Xsky130_fd_sc_hs__clkbuf_4_40 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__clkbuf_4_47/X
+ sky130_fd_sc_hs__clkbuf_4_41/X sky130_fd_sc_hs__clkbuf_4_41/a_83_270# sky130_fd_sc_hs__clkbuf_4
Xsky130_fd_sc_hs__clkbuf_4_51 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__clkbuf_4_51/A
+ sky130_fd_sc_hs__clkbuf_8_29/A sky130_fd_sc_hs__clkbuf_4_51/a_83_270# sky130_fd_sc_hs__clkbuf_4
Xsky130_fd_sc_hs__clkbuf_4_62 DVSS: DVDD: DVDD: DVSS: fine_control_avg_window_select[2]
+ sky130_fd_sc_hs__clkbuf_4_63/X sky130_fd_sc_hs__clkbuf_4_63/a_83_270# sky130_fd_sc_hs__clkbuf_4
Xsky130_fd_sc_hs__clkbuf_4_73 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__or2b_4_5/X
+ sky130_fd_sc_hs__o21ai_2_3/A2 sky130_fd_sc_hs__clkbuf_4_73/a_83_270# sky130_fd_sc_hs__clkbuf_4
Xsky130_fd_sc_hs__clkbuf_4_84 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__buf_2_131/X
+ sky130_fd_sc_hs__inv_4_23/A sky130_fd_sc_hs__clkbuf_4_85/a_83_270# sky130_fd_sc_hs__clkbuf_4
Xsky130_fd_sc_hs__clkbuf_4_95 DVSS: DVDD: DVDD: DVSS: div_ratio_half[2] sky130_fd_sc_hs__clkbuf_4_95/X
+ sky130_fd_sc_hs__clkbuf_4_95/a_83_270# sky130_fd_sc_hs__clkbuf_4
Xsky130_fd_sc_hs__clkinv_8_10 DVSS: DVDD: DVDD: DVSS: prbs_generator_syn_5/out hr_16t4_mux_top_3/din[7]
+ sky130_fd_sc_hs__clkinv_8
Xqr_4t1_mux_top_3 qr_4t1_mux_top_3/clk_Q hr_16t4_mux_top_3/clk qr_4t1_mux_top_3/clk_I
+ qr_4t1_mux_top_3/clk_IB qr_4t1_mux_top_3/din[3] qr_4t1_mux_top_3/din[2] qr_4t1_mux_top_3/din[1]
+ qr_4t1_mux_top_3/din[0] qr_4t1_mux_top_3/rst qr_4t1_mux_top_3/din_3_dummy qr_4t1_mux_top_3/din_3_dummy
+ qr_4t1_mux_top_3/din_3_dummy qr_4t1_mux_top_3/din_3_dummy dout_n qr_4t1_mux_top_3/mux_out_dummy
+ DVSS: DVDD: qr_4t1_mux_top_3/sky130_fd_sc_hs__dfxtp_2_1/a_1172_124# qr_4t1_mux_top_3/sky130_fd_sc_hs__dfxtp_2_3/a_1217_314#
+ qr_4t1_mux_top_3/sky130_fd_sc_hs__dfxtp_4_1/a_1141_508# qr_4t1_mux_top_3/sky130_fd_sc_hs__dfxtp_2_3/a_695_459#
+ qr_4t1_mux_top_3/sky130_fd_sc_hs__dfxtp_4_3/a_651_503# qr_4t1_mux_top_3/sky130_fd_sc_hs__dfxtp_2_1/a_538_429#
+ qr_4t1_mux_top_3/sky130_fd_sc_hs__mux4_1_1/A0 qr_4t1_mux_top_3/sky130_fd_sc_hs__mux4_1_1/a_264_74#
+ qr_4t1_mux_top_3/sky130_fd_sc_hs__dfxtp_2_1/a_1217_314# qr_4t1_mux_top_3/sky130_fd_sc_hs__mux4_1_1/a_1338_125#
+ qr_4t1_mux_top_3/sky130_fd_sc_hs__mux4_4_1/a_758_306# qr_4t1_mux_top_3/sky130_fd_sc_hs__mux4_1_1/A2
+ qr_4t1_mux_top_3/sky130_fd_sc_hs__dfxtp_2_7/a_206_368# qr_4t1_mux_top_3/sky130_fd_sc_hs__dfxtp_2_5/a_431_508#
+ qr_4t1_mux_top_3/sky130_fd_sc_hs__mux4_1_1/A1 qr_4t1_mux_top_3/sky130_fd_sc_hs__dfxtp_2_7/D
+ qr_4t1_mux_top_3/sky130_fd_sc_hs__dfxtp_4_1/a_206_368# qr_4t1_mux_top_3/sky130_fd_sc_hs__dfxtp_2_7/a_708_101#
+ qr_4t1_mux_top_3/sky130_fd_sc_hs__dfxtp_4_3/a_696_458# qr_4t1_mux_top_3/sky130_fd_sc_hs__dfxtp_2_9/a_644_504#
+ qr_4t1_mux_top_3/sky130_fd_sc_hs__mux4_1_1/X qr_4t1_mux_top_3/sky130_fd_sc_hs__dfxtp_2_11/a_206_368#
+ qr_4t1_mux_top_3/sky130_fd_sc_hs__dfxtp_4_1/a_437_503# qr_4t1_mux_top_3/sky130_fd_sc_hs__clkbuf_1_1/a_27_74#
+ qr_4t1_mux_top_3/sky130_fd_sc_hs__dfxtp_2_3/a_431_508# qr_4t1_mux_top_3/sky130_fd_sc_hs__dfxtp_4_3/a_544_485#
+ qr_4t1_mux_top_3/sky130_fd_sc_hs__dfxtp_2_9/a_538_429# qr_4t1_mux_top_3/sky130_fd_sc_hs__dfxtp_2_11/a_708_101#
+ qr_4t1_mux_top_3/sky130_fd_sc_hs__dfxtp_2_11/a_1125_508# qr_4t1_mux_top_3/sky130_fd_sc_hs__mux4_1_1/a_27_74#
+ qr_4t1_mux_top_3/sky130_fd_sc_hs__mux4_1_1/a_342_74# qr_4t1_mux_top_3/sky130_fd_sc_hs__dfxtp_2_11/a_27_74#
+ qr_4t1_mux_top_3/sky130_fd_sc_hs__dfxtp_2_1/a_695_459# qr_4t1_mux_top_3/sky130_fd_sc_hs__dfxtp_4_1/a_651_503#
+ qr_4t1_mux_top_3/sky130_fd_sc_hs__dfxtp_4_1/D qr_4t1_mux_top_3/sky130_fd_sc_hs__dfxtp_2_7/a_644_504#
+ qr_4t1_mux_top_3/sky130_fd_sc_hs__dfxtp_4_3/a_1178_124# qr_4t1_mux_top_3/sky130_fd_sc_hs__clkbuf_2_1/a_43_192#
+ qr_4t1_mux_top_3/sky130_fd_sc_hs__dfxtp_2_5/a_206_368# qr_4t1_mux_top_3/sky130_fd_sc_hs__clkbuf_1_5/X
+ qr_4t1_mux_top_3/sky130_fd_sc_hs__dfxtp_2_9/a_1125_508# qr_4t1_mux_top_3/sky130_fd_sc_hs__clkbuf_2_3/X
+ qr_4t1_mux_top_3/sky130_fd_sc_hs__dfxtp_2_7/a_538_429# qr_4t1_mux_top_3/sky130_fd_sc_hs__dfxtp_2_9/Q
+ qr_4t1_mux_top_3/sky130_fd_sc_hs__dfxtp_4_1/a_1178_124# qr_4t1_mux_top_3/sky130_fd_sc_hs__dfxtp_2_11/a_644_504#
+ qr_4t1_mux_top_3/sky130_fd_sc_hs__dfxtp_4_1/a_696_458# qr_4t1_mux_top_3/sky130_fd_sc_hs__dfxtp_2_5/a_27_74#
+ qr_4t1_mux_top_3/sky130_fd_sc_hs__dfxtp_2_5/a_708_101# qr_4t1_mux_top_3/sky130_fd_sc_hs__dfxtp_4_1/a_27_74#
+ qr_4t1_mux_top_3/sky130_fd_sc_hs__mux4_4_1/a_1285_377# qr_4t1_mux_top_3/sky130_fd_sc_hs__dfxtp_2_7/a_1125_508#
+ qr_4t1_mux_top_3/sky130_fd_sc_hs__mux4_1_1/a_537_341# qr_4t1_mux_top_3/sky130_fd_sc_hs__mux4_1_1/a_255_341#
+ qr_4t1_mux_top_3/sky130_fd_sc_hs__mux4_4_1/A0 qr_4t1_mux_top_3/sky130_fd_sc_hs__clkbuf_1_3/X
+ qr_4t1_mux_top_3/sky130_fd_sc_hs__mux4_1_1/A3 qr_4t1_mux_top_3/sky130_fd_sc_hs__dfxtp_2_11/a_538_429#
+ qr_4t1_mux_top_3/sky130_fd_sc_hs__dfxtp_2_3/a_206_368# qr_4t1_mux_top_3/sky130_fd_sc_hs__dfxtp_2_1/a_431_508#
+ qr_4t1_mux_top_3/sky130_fd_sc_hs__clkbuf_1_1/X qr_4t1_mux_top_3/sky130_fd_sc_hs__dfxtp_2_9/a_695_459#
+ qr_4t1_mux_top_3/sky130_fd_sc_hs__dfxtp_4_1/a_544_485# qr_4t1_mux_top_3/sky130_fd_sc_hs__dfxtp_2_5/a_1125_508#
+ qr_4t1_mux_top_3/sky130_fd_sc_hs__mux4_4_1/A2 qr_4t1_mux_top_3/sky130_fd_sc_hs__dfxtp_2_7/a_27_74#
+ qr_4t1_mux_top_3/sky130_fd_sc_hs__dfxtp_2_3/a_708_101# qr_4t1_mux_top_3/sky130_fd_sc_hs__dfxtp_2_3/a_1125_508#
+ qr_4t1_mux_top_3/sky130_fd_sc_hs__dfxtp_4_3/a_27_74# qr_4t1_mux_top_3/sky130_fd_sc_hs__dfxtp_2_11/a_1019_424#
+ qr_4t1_mux_top_3/sky130_fd_sc_hs__mux4_1_1/a_450_74# qr_4t1_mux_top_3/sky130_fd_sc_hs__dfxtp_4_3/a_1034_424#
+ qr_4t1_mux_top_3/sky130_fd_sc_hs__clkbuf_1_3/a_27_74# qr_4t1_mux_top_3/sky130_fd_sc_hs__dfxtp_2_1/a_1125_508#
+ qr_4t1_mux_top_3/sky130_fd_sc_hs__mux4_4_1/a_114_126# qr_4t1_mux_top_3/sky130_fd_sc_hs__dfxtp_2_1/a_27_74#
+ qr_4t1_mux_top_3/sky130_fd_sc_hs__dfxtp_2_5/a_644_504# qr_4t1_mux_top_3/sky130_fd_sc_hs__dfxtp_4_1/a_1034_424#
+ qr_4t1_mux_top_3/sky130_fd_sc_hs__dfxtp_2_11/a_1172_124# qr_4t1_mux_top_3/sky130_fd_sc_hs__mux4_4_1/a_1450_121#
+ qr_4t1_mux_top_3/sky130_fd_sc_hs__dfxtp_2_9/a_431_508# qr_4t1_mux_top_3/sky130_fd_sc_hs__dfxtp_2_7/a_695_459#
+ qr_4t1_mux_top_3/sky130_fd_sc_hs__mux4_4_1/a_1191_121# qr_4t1_mux_top_3/sky130_fd_sc_hs__mux4_1_1/a_768_74#
+ qr_4t1_mux_top_3/sky130_fd_sc_hs__dfxtp_2_5/a_538_429# qr_4t1_mux_top_3/sky130_fd_sc_hs__dfxtp_2_9/a_1019_424#
+ qr_4t1_mux_top_3/sky130_fd_sc_hs__mux4_1_1/a_1396_99# qr_4t1_mux_top_3/sky130_fd_sc_hs__dfxtp_2_3/a_644_504#
+ qr_4t1_mux_top_3/sky130_fd_sc_hs__mux4_1_1/a_1065_387# qr_4t1_mux_top_3/sky130_fd_sc_hs__dfxtp_4_3/a_735_102#
+ qr_4t1_mux_top_3/sky130_fd_sc_hs__dfxtp_2_3/a_27_74# qr_4t1_mux_top_3/sky130_fd_sc_hs__dfxtp_2_11/a_695_459#
+ qr_4t1_mux_top_3/sky130_fd_sc_hs__dfxtp_2_11/a_1217_314# qr_4t1_mux_top_3/sky130_fd_sc_hs__dfxtp_2_7/a_1019_424#
+ qr_4t1_mux_top_3/sky130_fd_sc_hs__dfxtp_2_1/a_206_368# qr_4t1_mux_top_3/sky130_fd_sc_hs__mux4_4_1/a_1278_121#
+ qr_4t1_mux_top_3/sky130_fd_sc_hs__dfxtp_2_3/a_538_429# qr_4t1_mux_top_3/sky130_fd_sc_hs__dfxtp_4_3/a_1226_296#
+ qr_4t1_mux_top_3/sky130_fd_sc_hs__dfxtp_2_1/a_708_101# qr_4t1_mux_top_3/sky130_fd_sc_hs__dfxtp_2_9/a_1172_124#
+ qr_4t1_mux_top_3/sky130_fd_sc_hs__mux4_4_1/a_509_392# qr_4t1_mux_top_3/sky130_fd_sc_hs__dfxtp_2_5/a_1019_424#
+ qr_4t1_mux_top_3/sky130_fd_sc_hs__dfxtp_2_3/a_1019_424# qr_4t1_mux_top_3/sky130_fd_sc_hs__dfxtp_2_7/a_431_508#
+ qr_4t1_mux_top_3/sky130_fd_sc_hs__dfxtp_2_7/a_1172_124# qr_4t1_mux_top_3/sky130_fd_sc_hs__dfxtp_4_1/a_1226_296#
+ qr_4t1_mux_top_3/sky130_fd_sc_hs__mux4_4_1/a_1465_377# qr_4t1_mux_top_3/sky130_fd_sc_hs__mux4_1_1/a_846_74#
+ qr_4t1_mux_top_3/sky130_fd_sc_hs__mux4_4_1/a_2199_74# qr_4t1_mux_top_3/sky130_fd_sc_hs__dfxtp_2_9/a_1217_314#
+ qr_4t1_mux_top_3/sky130_fd_sc_hs__dfxtp_4_3/a_206_368# qr_4t1_mux_top_3/sky130_fd_sc_hs__clkbuf_2_3/a_43_192#
+ qr_4t1_mux_top_3/sky130_fd_sc_hs__mux4_4_1/a_296_392# qr_4t1_mux_top_3/sky130_fd_sc_hs__dfxtp_2_1/a_1019_424#
+ qr_4t1_mux_top_3/sky130_fd_sc_hs__dfxtp_4_3/a_437_503# qr_4t1_mux_top_3/sky130_fd_sc_hs__dfxtp_2_11/a_431_508#
+ qr_4t1_mux_top_3/sky130_fd_sc_hs__dfxtp_2_5/a_1172_124# qr_4t1_mux_top_3/sky130_fd_sc_hs__dfxtp_2_9/a_27_74#
+ qr_4t1_mux_top_3/sky130_fd_sc_hs__dfxtp_2_7/a_1217_314# qr_4t1_mux_top_3/sky130_fd_sc_hs__dfxtp_2_9/a_206_368#
+ qr_4t1_mux_top_3/sky130_fd_sc_hs__dfxtp_2_3/a_1172_124# qr_4t1_mux_top_3/sky130_fd_sc_hs__dfxtp_2_5/a_695_459#
+ qr_4t1_mux_top_3/sky130_fd_sc_hs__mux4_4_1/a_2489_347# qr_4t1_mux_top_3/sky130_fd_sc_hs__mux4_1_1/a_763_341#
+ qr_4t1_mux_top_3/sky130_fd_sc_hs__dfxtp_4_3/a_1141_508# qr_4t1_mux_top_3/sky130_fd_sc_hs__mux4_4_1/a_299_126#
+ qr_4t1_mux_top_3/sky130_fd_sc_hs__dfxtp_2_9/a_708_101# qr_4t1_mux_top_3/sky130_fd_sc_hs__mux4_4_1/a_116_392#
+ qr_4t1_mux_top_3/sky130_fd_sc_hs__dfxtp_2_1/a_644_504# qr_4t1_mux_top_3/sky130_fd_sc_hs__mux4_1_1/a_979_74#
+ qr_4t1_mux_top_3/sky130_fd_sc_hs__dfxtp_2_5/a_1217_314# qr_4t1_mux_top_3/sky130_fd_sc_hs__dfxtp_4_1/a_735_102#
+ qr_4t1_mux_top_3/sky130_fd_sc_hs__clkbuf_1_5/a_27_74# qr_4t1_mux_top
Xsky130_fd_sc_hs__inv_4_19 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__inv_4_19/Y sky130_fd_sc_hs__inv_4_19/A
+ sky130_fd_sc_hs__inv_4
Xsky130_fd_sc_hs__conb_1_130 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__conb_1_131/LO
+ sky130_fd_sc_hs__conb_1_131/HI sky130_fd_sc_hs__conb_1_131/a_165_290# sky130_fd_sc_hs__conb_1_131/a_21_290#
+ sky130_fd_sc_hs__conb_1
Xsky130_fd_sc_hs__conb_1_141 DVSS: DVDD: DVDD: DVSS: prbs_generator_syn_15/eqn[30]
+ sky130_fd_sc_hs__conb_1_141/HI sky130_fd_sc_hs__conb_1_141/a_165_290# sky130_fd_sc_hs__conb_1_141/a_21_290#
+ sky130_fd_sc_hs__conb_1
Xsky130_fd_sc_hs__conb_1_152 DVSS: DVDD: DVDD: DVSS: prbs_generator_syn_17/eqn[9]
+ sky130_fd_sc_hs__conb_1_153/HI sky130_fd_sc_hs__conb_1_153/a_165_290# sky130_fd_sc_hs__conb_1_153/a_21_290#
+ sky130_fd_sc_hs__conb_1
Xsky130_fd_sc_hs__conb_1_163 DVSS: DVDD: DVDD: DVSS: prbs_generator_syn_17/eqn[2]
+ prbs_generator_syn_17/eqn[1] sky130_fd_sc_hs__conb_1_163/a_165_290# sky130_fd_sc_hs__conb_1_163/a_21_290#
+ sky130_fd_sc_hs__conb_1
Xsky130_fd_sc_hs__conb_1_174 DVSS: DVDD: DVDD: DVSS: prbs_generator_syn_23/eqn[9]
+ sky130_fd_sc_hs__conb_1_175/HI sky130_fd_sc_hs__conb_1_175/a_165_290# sky130_fd_sc_hs__conb_1_175/a_21_290#
+ sky130_fd_sc_hs__conb_1
Xsky130_fd_sc_hs__conb_1_185 DVSS: DVDD: DVDD: DVSS: prbs_generator_syn_29/eqn[9]
+ sky130_fd_sc_hs__conb_1_185/HI sky130_fd_sc_hs__conb_1_185/a_165_290# sky130_fd_sc_hs__conb_1_185/a_21_290#
+ sky130_fd_sc_hs__conb_1
Xsky130_fd_sc_hs__conb_1_196 DVSS: DVDD: DVDD: DVSS: prbs_generator_syn_19/eqn[22]
+ prbs_generator_syn_19/eqn[20] sky130_fd_sc_hs__conb_1_197/a_165_290# sky130_fd_sc_hs__conb_1_197/a_21_290#
+ sky130_fd_sc_hs__conb_1
Xosc_core_1 osc_core_1/glob_en osc_core_1/delay_con_lsb[4] osc_core_1/delay_con_lsb[3]
+ osc_core_1/delay_con_lsb[2] osc_core_1/delay_con_lsb[1] osc_core_1/delay_con_lsb[0]
+ osc_core_1/delay_con_msb[7] osc_core_1/delay_con_msb[6] osc_core_1/delay_con_msb[5]
+ osc_core_1/delay_con_msb[4] osc_core_1/delay_con_msb[3] osc_core_1/delay_con_msb[2]
+ osc_core_1/delay_con_msb[1] osc_core_1/delay_con_msb[0] osc_core_1/con_perb_5[3]
+ osc_core_1/con_perb_5[2] osc_core_1/con_perb_5[1] osc_core_1/con_perb_5[0] osc_core_1/con_perb_5[3]
+ osc_core_1/con_perb_5[2] osc_core_1/con_perb_5[1] osc_core_1/con_perb_5[0] osc_core_1/con_perb_5[3]
+ osc_core_1/con_perb_5[2] osc_core_1/con_perb_5[1] osc_core_1/con_perb_5[0] osc_core_1/con_perb_5[3]
+ osc_core_1/con_perb_5[2] osc_core_1/con_perb_5[1] osc_core_1/con_perb_5[0] osc_core_1/con_perb_5[3]
+ osc_core_1/con_perb_5[2] osc_core_1/con_perb_5[1] osc_core_1/con_perb_5[0] osc_core_1/ref_clk
+ osc_core_1/pi1_l[3] osc_core_1/pi1_l[2] osc_core_1/pi1_l[1] osc_core_1/pi1_l[0]
+ osc_core_1/pi1_r[3] osc_core_1/pi1_r[2] osc_core_1/pi1_r[1] osc_core_1/pi1_r[0]
+ osc_core_1/pi2_l[3] osc_core_1/pi2_l[2] osc_core_1/pi2_l[1] osc_core_1/pi2_l[0]
+ osc_core_1/pi2_r[3] osc_core_1/pi2_r[2] osc_core_1/pi2_r[1] osc_core_1/pi2_r[0]
+ osc_core_1/pi3_l[3] osc_core_1/pi3_l[2] osc_core_1/pi3_l[1] osc_core_1/pi3_l[0]
+ osc_core_1/pi3_r[3] osc_core_1/pi3_r[2] osc_core_1/pi3_r[1] osc_core_1/pi3_r[0]
+ osc_core_1/pi4_l[3] osc_core_1/pi4_l[2] osc_core_1/pi4_l[1] osc_core_1/pi4_l[0]
+ osc_core_1/pi4_r[3] osc_core_1/pi4_r[2] osc_core_1/pi4_r[1] osc_core_1/pi4_r[0]
+ osc_core_1/pi5_l[3] osc_core_1/pi5_l[2] osc_core_1/pi5_l[1] osc_core_1/pi5_l[0]
+ osc_core_1/pi5_r[3] osc_core_1/pi5_r[2] osc_core_1/pi5_r[1] osc_core_1/pi5_r[0]
+ osc_core_1/osc_000 osc_core_1/osc_036 osc_core_1/osc_072 osc_core_1/osc_108 osc_core_1/osc_144
+ osc_core_1/inj_en osc_core_1/inj_out osc_core_1/osc_hold osc_core_1/p1 osc_core_1/p2
+ osc_core_1/p3 osc_core_1/p4 osc_core_1/p5 DVSS: AVDD osc_core_1/sky130_fd_sc_hs__einvp_2_5/a_36_74#
+ osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_75/X osc_core_1/sky130_fd_sc_hs__nand2_2_93/Y
+ osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_1/X osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_11/a_28_74#
+ osc_core_1/sky130_fd_sc_hs__inv_4_5/Y osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_27/a_289_74#
+ osc_core_1/sky130_fd_sc_hs__nand2_8_9/B osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_7/a_405_138#
+ osc_core_1/sky130_fd_sc_hs__nand2_4_40/a_27_74# osc_core_1/sky130_fd_sc_hs__dfrtp_4_3/a_890_138#
+ osc_core_1/sky130_fd_sc_hs__nand2_1_9/B osc_core_1/sky130_fd_sc_hs__nand2_4_137/a_27_74#
+ osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_56/A osc_core_1/sky130_fd_sc_hs__inv_4_17/Y
+ osc_core_1/sky130_fd_sc_hs__nand2_2_55/Y osc_core_1/sky130_fd_sc_hs__nand2_8_31/a_27_74#
+ osc_core_1/sky130_fd_sc_hs__nand2_4_53/a_27_74# osc_core_1/sky130_fd_sc_hs__nand2_4_123/Y
+ osc_core_1/sky130_fd_sc_hs__einvp_1_1/a_44_549# osc_core_1/sky130_fd_sc_hs__nand2_1_5/a_117_74#
+ osc_core_1/sky130_fd_sc_hs__inv_4_3/Y osc_core_1/sky130_fd_sc_hs__nand2_2_69/a_27_74#
+ osc_core_1/sky130_fd_sc_hs__einvp_2_11/a_263_323# osc_core_1/sky130_fd_sc_hs__einvp_8_3/a_27_368#
+ osc_core_1/sky130_fd_sc_hs__nand2_2_84/B osc_core_1/sky130_fd_sc_hs__a21oi_1_9/a_29_368#
+ osc_core_1/sky130_fd_sc_hs__nand2_4_51/Y osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_68/X
+ osc_core_1/sky130_fd_sc_hs__einvp_4_9/a_473_323# osc_core_1/sky130_fd_sc_hs__nand2_2_109/a_27_74#
+ osc_core_1/sky130_fd_sc_hs__inv_16_3/Y osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_31/X
+ osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_5/A osc_core_1/sky130_fd_sc_hs__nand2_2_45/B
+ osc_core_1/sky130_fd_sc_hs__nand2_2_3/a_27_74# osc_core_1/sky130_fd_sc_hs__einvp_8_14/a_802_323#
+ osc_core_1/sky130_fd_sc_hs__einvp_2_19/a_36_74# osc_core_1/sky130_fd_sc_hs__nand2_4_15/Y
+ osc_core_1/sky130_fd_sc_hs__nand2_4_153/Y osc_core_1/sky130_fd_sc_hs__nand2_4_107/a_27_74#
+ osc_core_1/sky130_fd_sc_hs__and4_2_3/X osc_core_1/sky130_fd_sc_hs__and2_2_1/a_118_74#
+ osc_core_1/sky130_fd_sc_hs__nand2_4_93/a_27_74# osc_core_1/sky130_fd_sc_hs__einvp_1_5/a_44_549#
+ osc_core_1/sky130_fd_sc_hs__nand2_1_9/a_117_74# osc_core_1/sky130_fd_sc_hs__and4_2_3/a_335_74#
+ osc_core_1/sky130_fd_sc_hs__a21oi_1_49/Y osc_core_1/sky130_fd_sc_hs__einvp_1_5/a_310_392#
+ osc_core_1/sky130_fd_sc_hs__einvp_8_5/a_27_368# osc_core_1/sky130_fd_sc_hs__inv_16_9/Y
+ osc_core_1/sky130_fd_sc_hs__nand2_4_45/Y osc_core_1/sky130_fd_sc_hs__a21oi_1_43/a_29_368#
+ osc_core_1/sky130_fd_sc_hs__nand2_2_77/Y osc_core_1/sky130_fd_sc_hs__clkbuf_2_3/A
+ osc_core_1/sky130_fd_sc_hs__nand2_4_9/a_27_74# osc_core_1/sky130_fd_sc_hs__nand2_8_25/a_27_74#
+ osc_core_1/sky130_fd_sc_hs__inv_16_1/Y osc_core_1/sky130_fd_sc_hs__einvp_4_17/a_473_323#
+ osc_core_1/sky130_fd_sc_hs__nand2_2_53/a_27_74# osc_core_1/sky130_fd_sc_hs__inv_16_13/Y
+ osc_core_1/sky130_fd_sc_hs__nand2_4_47/a_27_74# osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_78/a_289_74#
+ osc_core_1/sky130_fd_sc_hs__inv_8_3/A osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_14/a_289_74#
+ osc_core_1/sky130_fd_sc_hs__inv_8_9/A osc_core_1/sky130_fd_sc_hs__nand2_4_75/Y osc_core_1/sky130_fd_sc_hs__nand2_4_61/a_27_74#
+ osc_core_1/sky130_fd_sc_hs__nand2_4_110/Y osc_core_1/sky130_fd_sc_hs__inv_4_9/Y
+ osc_core_1/sky130_fd_sc_hs__einvp_1_9/a_44_549# osc_core_1/sky130_fd_sc_hs__inv_4_7/Y
+ osc_core_1/sky130_fd_sc_hs__einvp_8_8/a_27_368# osc_core_1/sky130_fd_sc_hs__inv_4_23/Y
+ osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_78/a_405_138# osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_45/a_28_74#
+ osc_core_1/sky130_fd_sc_hs__nand2_2_77/a_27_74# osc_core_1/sky130_fd_sc_hs__nand2_2_23/Y
+ osc_core_1/sky130_fd_sc_hs__einvp_8_9/a_27_368# osc_core_1/sky130_fd_sc_hs__clkbuf_4_3/X
+ osc_core_1/sky130_fd_sc_hs__nand2_4_40/Y osc_core_1/sky130_fd_sc_hs__a21oi_1_13/a_29_368#
+ osc_core_1/sky130_fd_sc_hs__nand2_1_3/B osc_core_1/sky130_fd_sc_hs__nand2_8_1/a_27_74#
+ osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_25/X osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_71/X
+ osc_core_1/sky130_fd_sc_hs__nand2_2_21/a_27_74# osc_core_1/sky130_fd_sc_hs__inv_4_1/Y
+ osc_core_1/sky130_fd_sc_hs__nand2_4_87/a_27_74# osc_core_1/sky130_fd_sc_hs__nand2_4_139/Y
+ osc_core_1/sky130_fd_sc_hs__nand2_4_115/a_27_74# osc_core_1/sky130_fd_sc_hs__dlygate4sd2_1_1/a_28_74#
+ osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_17/a_289_74# osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_5/a_405_138#
+ osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_79/A osc_core_1/sky130_fd_sc_hs__clkbuf_2_14/a_43_192#
+ osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_62/a_289_74# osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_35/X
+ osc_core_1/sky130_fd_sc_hs__nand2_2_53/Y osc_core_1/sky130_fd_sc_hs__nand2_4_31/a_27_74#
+ osc_core_1/sky130_fd_sc_hs__nand2_8_19/a_27_74# osc_core_1/sky130_fd_sc_hs__einvp_8_14/a_27_368#
+ osc_core_1/sky130_fd_sc_hs__inv_4_25/Y osc_core_1/sky130_fd_sc_hs__inv_8_1/A osc_core_1/sky130_fd_sc_hs__inv_4_15/Y
+ osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_15/a_28_74# osc_core_1/sky130_fd_sc_hs__nand2_2_47/a_27_74#
+ osc_core_1/sky130_fd_sc_hs__and2_2_3/X osc_core_1/sky130_fd_sc_hs__nand2_2_15/Y
+ osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_3/a_289_74# osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_63/A
+ osc_core_1/sky130_fd_sc_hs__a21oi_1_17/a_29_368# osc_core_1/sky130_fd_sc_hs__nand2_8_33/a_27_74#
+ osc_core_1/sky130_fd_sc_hs__einvp_8_9/a_802_323# osc_core_1/sky130_fd_sc_hs__inv_16_5/Y
+ osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_65/X osc_core_1/sky130_fd_sc_hs__nand2_2_85/Y
+ osc_core_1/sky130_fd_sc_hs__nand2_2_61/a_27_74# osc_core_1/sky130_fd_sc_hs__einvp_2_1/a_263_323#
+ osc_core_1/sky130_fd_sc_hs__nand2_4_155/a_27_74# osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_57/X
+ osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_21/a_405_138# osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_59/a_405_138#
+ osc_core_1/sky130_fd_sc_hs__a21oi_1_47/a_117_74# osc_core_1/sky130_fd_sc_hs__nand2_4_13/Y
+ osc_core_1/sky130_fd_sc_hs__nand2_4_151/Y osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_39/a_28_74#
+ osc_core_1/sky130_fd_sc_hs__nand2_2_61/B osc_core_1/sky130_fd_sc_hs__inv_4_11/Y
+ osc_core_1/sky130_fd_sc_hs__nand2_2_102/a_27_74# osc_core_1/sky130_fd_sc_hs__einvp_2_13/a_27_368#
+ osc_core_1/sky130_fd_sc_hs__einvp_8_15/a_802_323# osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_65/a_289_74#
+ osc_core_1/sky130_fd_sc_hs__nand2_4_71/a_27_74# osc_core_1/sky130_fd_sc_hs__einvp_8_19/a_27_368#
+ osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_53/a_28_74# osc_core_1/sky130_fd_sc_hs__nand2_2_88/a_27_74#
+ osc_core_1/sky130_fd_sc_hs__nand2_2_15/a_27_74# osc_core_1/sky130_fd_sc_hs__nand2_2_5/a_27_74#
+ osc_core_1/sky130_fd_sc_hs__and4_2_3/C osc_core_1/sky130_fd_sc_hs__a21oi_1_45/Y
+ osc_core_1/sky130_fd_sc_hs__nand2_4_110/a_27_74# osc_core_1/sky130_fd_sc_hs__inv_16_7/Y
+ osc_core_1/sky130_fd_sc_hs__einvp_4_5/a_27_368# osc_core_1/sky130_fd_sc_hs__nand2_2_99/B
+ osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_49/a_405_138# osc_core_1/sky130_fd_sc_hs__a21oi_1_33/a_29_368#
+ osc_core_1/sky130_fd_sc_hs__clkbuf_2_1/A osc_core_1/sky130_fd_sc_hs__nand2_2_5/B
+ osc_core_1/sky130_fd_sc_hs__nand2_2_31/a_27_74# osc_core_1/sky130_fd_sc_hs__nand2_4_25/a_27_74#
+ osc_core_1/sky130_fd_sc_hs__inv_4_36/Y osc_core_1/sky130_fd_sc_hs__nand2_2_9/B osc_core_1/sky130_fd_sc_hs__inv_4_39/Y
+ osc_core_1/sky130_fd_sc_hs__nand2_2_9/Y osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_78/a_28_74#
+ osc_core_1/sky130_fd_sc_hs__dfrtp_4_3/a_313_74# osc_core_1/sky130_fd_sc_hs__nand2_2_39/Y
+ osc_core_1/sky130_fd_sc_hs__and4_2_1/a_143_74# osc_core_1/sky130_fd_sc_hs__inv_8_7/A
+ osc_core_1/sky130_fd_sc_hs__nand2_8_27/a_27_74# osc_core_1/sky130_fd_sc_hs__nand2_4_73/Y
+ osc_core_1/sky130_fd_sc_hs__buf_4_1/a_86_260# osc_core_1/sky130_fd_sc_hs__inv_4_33/Y
+ osc_core_1/sky130_fd_sc_hs__dfrtp_4_3/a_494_366# osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_23/a_28_74#
+ osc_core_1/sky130_fd_sc_hs__clkbuf_4_3/a_83_270# osc_core_1/sky130_fd_sc_hs__einvp_1_19/a_310_392#
+ osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_49/X osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_39/a_405_138#
+ osc_core_1/sky130_fd_sc_hs__clkbuf_2_9/a_43_192# osc_core_1/sky130_fd_sc_hs__nand2_8_43/a_27_74#
+ osc_core_1/sky130_fd_sc_hs__nand2_4_35/Y osc_core_1/sky130_fd_sc_hs__einvp_4_9/a_27_368#
+ osc_core_1/sky130_fd_sc_hs__nand2_2_69/Y osc_core_1/sky130_fd_sc_hs__a21oi_1_35/a_29_368#
+ osc_core_1/sky130_fd_sc_hs__nand2_1_1/B osc_core_1/sky130_fd_sc_hs__nand2_2_71/a_27_74#
+ osc_core_1/sky130_fd_sc_hs__inv_4_29/Y osc_core_1/sky130_fd_sc_hs__nand2_4_65/a_27_74#
+ osc_core_1/sky130_fd_sc_hs__nand2_2_43/B osc_core_1/sky130_fd_sc_hs__dfrtp_4_1/a_1647_81#
+ osc_core_1/sky130_fd_sc_hs__nand2_4_137/Y osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_47/a_28_74#
+ osc_core_1/sky130_fd_sc_hs__and4_2_5/a_143_74# osc_core_1/sky130_fd_sc_hs__a21oi_1_32/a_117_74#
+ osc_core_1/sky130_fd_sc_hs__einvp_2_5/a_27_368# osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_45/A
+ osc_core_1/sky130_fd_sc_hs__nand2_2_97/B osc_core_1/sky130_fd_sc_hs__inv_8_5/A osc_core_1/sky130_fd_sc_hs__nand2_2_51/Y
+ osc_core_1/sky130_fd_sc_hs__dfrtp_4_1/a_890_138# osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_29/a_405_138#
+ osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_69/a_405_138# osc_core_1/sky130_fd_sc_hs__nand2_2_97/a_27_74#
+ osc_core_1/sky130_fd_sc_hs__nand2_2_25/a_27_74# osc_core_1/sky130_fd_sc_hs__nand2_2_99/Y
+ osc_core_1/sky130_fd_sc_hs__nand2_4_19/a_27_74# osc_core_1/sky130_fd_sc_hs__nand2_4_117/a_27_74#
+ osc_core_1/sky130_fd_sc_hs__inv_16_9/A osc_core_1/sky130_fd_sc_hs__nand2_4_29/Y
+ osc_core_1/sky130_fd_sc_hs__einvp_8_19/a_27_74# osc_core_1/sky130_fd_sc_hs__nand2_2_85/B
+ osc_core_1/sky130_fd_sc_hs__einvp_2_19/a_263_323# osc_core_1/sky130_fd_sc_hs__dfrtp_4_3/D
+ osc_core_1/sky130_fd_sc_hs__nand2_2_83/Y osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_17/a_28_74#
+ osc_core_1/sky130_fd_sc_hs__einvp_4_7/a_473_323# osc_core_1/sky130_fd_sc_hs__nand2_4_11/Y
+ osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_20/a_405_138# osc_core_1/sky130_fd_sc_hs__a21oi_1_37/a_117_74#
+ osc_core_1/sky130_fd_sc_hs__einvp_2_9/a_27_368# osc_core_1/sky130_fd_sc_hs__nand2_8_37/a_27_74#
+ osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_56/a_289_74# osc_core_1/sky130_fd_sc_hs__inv_4_31/Y
+ osc_core_1/sky130_fd_sc_hs__inv_1_9/Y osc_core_1/sky130_fd_sc_hs__nand2_2_65/a_27_74#
+ osc_core_1/sky130_fd_sc_hs__inv_16_31/A osc_core_1/sky130_fd_sc_hs__einvp_4_7/a_27_74#
+ osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_9/A osc_core_1/sky130_fd_sc_hs__and2_2_1/B
+ osc_core_1/sky130_fd_sc_hs__nand2_4_159/Y osc_core_1/sky130_fd_sc_hs__einvp_1_3/a_318_74#
+ osc_core_1/sky130_fd_sc_hs__nand2_2_71/B osc_core_1/sky130_fd_sc_hs__inv_4_19/Y
+ osc_core_1/sky130_fd_sc_hs__einvp_2_15/a_36_74# osc_core_1/sky130_fd_sc_hs__nand2_2_108/Y
+ osc_core_1/sky130_fd_sc_hs__buf_4_1/X osc_core_1/sky130_fd_sc_hs__nand2_2_73/Y osc_core_1/sky130_fd_sc_hs__einvp_1_3/a_310_392#
+ osc_core_1/sky130_fd_sc_hs__nand2_4_89/Y osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_47/a_405_138#
+ osc_core_1/sky130_fd_sc_hs__nand2_2_19/a_27_74# osc_core_1/sky130_fd_sc_hs__nand2_2_9/a_27_74#
+ osc_core_1/sky130_fd_sc_hs__nand2_2_57/B osc_core_1/sky130_fd_sc_hs__einvp_4_15/a_473_323#
+ osc_core_1/sky130_fd_sc_hs__nand2_2_37/Y osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_59/a_289_74#
+ osc_core_1/sky130_fd_sc_hs__einvp_1_11/a_44_549# osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_71/a_28_74#
+ osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_25/a_289_74# osc_core_1/sky130_fd_sc_hs__clkbuf_2_9/A
+ osc_core_1/sky130_fd_sc_hs__nand2_4_99/a_27_74# osc_core_1/sky130_fd_sc_hs__nand2_4_27/a_27_74#
+ osc_core_1/sky130_fd_sc_hs__nand2_4_71/Y osc_core_1/sky130_fd_sc_hs__dlygate4sd2_1_1/X
+ osc_core_1/sky130_fd_sc_hs__nand2_4_106/Y osc_core_1/sky130_fd_sc_hs__nand2_4_127/a_27_74#
+ osc_core_1/sky130_fd_sc_hs__a21oi_1_1/a_117_74# osc_core_1/sky130_fd_sc_hs__and4_2_5/D
+ osc_core_1/sky130_fd_sc_hs__nand2_4_5/a_27_74# osc_core_1/sky130_fd_sc_hs__einvp_1_7/a_318_74#
+ osc_core_1/sky130_fd_sc_hs__einvp_8_9/a_27_74# osc_core_1/sky130_fd_sc_hs__conb_1_1/LO
+ osc_core_1/sky130_fd_sc_hs__nand2_2_67/Y osc_core_1/sky130_fd_sc_hs__einvp_4_11/a_27_368#
+ osc_core_1/sky130_fd_sc_hs__inv_4_37/Y osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_25/a_28_74#
+ osc_core_1/sky130_fd_sc_hs__einvp_8_2/a_27_368# osc_core_1/sky130_fd_sc_hs__nand3_4_3/a_27_82#
+ osc_core_1/sky130_fd_sc_hs__dfrtp_4_3/a_2010_409# osc_core_1/sky130_fd_sc_hs__einvp_1_15/a_44_549#
+ osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_41/a_28_74# osc_core_1/sky130_fd_sc_hs__nand2_2_73/a_27_74#
+ osc_core_1/sky130_fd_sc_hs__a21oi_1_23/a_117_74# osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_75/a_289_74#
+ osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_3/a_405_138# osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_78/X
+ osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_41/a_289_74# osc_core_1/sky130_fd_sc_hs__a21oi_1_5/a_117_74#
+ osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_68/a_405_138# osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_59/X
+ osc_core_1/sky130_fd_sc_hs__nand2_2_13/Y osc_core_1/sky130_fd_sc_hs__nand2_4_83/a_27_74#
+ osc_core_1/sky130_fd_sc_hs__inv_4_21/Y osc_core_1/sky130_fd_sc_hs__nand2_2_59/Y
+ osc_core_1/sky130_fd_sc_hs__einvp_4_15/a_27_368# osc_core_1/sky130_fd_sc_hs__einvp_4_19/a_27_74#
+ osc_core_1/sky130_fd_sc_hs__nand2_8_7/a_27_74# osc_core_1/sky130_fd_sc_hs__a21oi_1_29/a_29_368#
+ osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_62/X osc_core_1/sky130_fd_sc_hs__nand2_2_99/a_27_74#
+ osc_core_1/sky130_fd_sc_hs__einvp_8_7/a_802_323# osc_core_1/sky130_fd_sc_hs__a21oi_1_42/a_29_368#
+ osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_1/a_28_74# osc_core_1/sky130_fd_sc_hs__nand2_8_15/a_27_74#
+ osc_core_1/sky130_fd_sc_hs__dfrtp_4_1/a_37_78# osc_core_1/sky130_fd_sc_hs__einvp_2_9/a_263_323#
+ osc_core_1/sky130_fd_sc_hs__einvp_1_19/a_44_549# osc_core_1/sky130_fd_sc_hs__nand2_2_88/B
+ osc_core_1/sky130_fd_sc_hs__nand2_2_43/Y osc_core_1/sky130_fd_sc_hs__nand3_4_3/a_456_82#
+ osc_core_1/sky130_fd_sc_hs__and4_2_5/a_56_74# osc_core_1/sky130_fd_sc_hs__nand2_4_57/Y
+ osc_core_1/sky130_fd_sc_hs__nand2_4_39/a_27_74# osc_core_1/sky130_fd_sc_hs__inv_1_7/Y
+ osc_core_1/sky130_fd_sc_hs__nand2_4_135/a_27_74# osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_45/a_289_74#
+ osc_core_1/sky130_fd_sc_hs__a21oi_1_9/a_117_74# osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_21/a_28_74#
+ osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_7/A osc_core_1/sky130_fd_sc_hs__and2_2_1/A
+ osc_core_1/sky130_fd_sc_hs__dfrtp_4_1/a_2010_409# osc_core_1/sky130_fd_sc_hs__einvp_4_1/a_27_74#
+ osc_core_1/sky130_fd_sc_hs__nand2_4_51/a_27_74# osc_core_1/sky130_fd_sc_hs__clkbuf_4_1/A
+ osc_core_1/sky130_fd_sc_hs__nand2_4_151/a_27_74# osc_core_1/sky130_fd_sc_hs__einvp_4_19/a_27_368#
+ osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_35/a_28_74# osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_53/X
+ osc_core_1/sky130_fd_sc_hs__nand2_4_87/Y osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_7/X
+ osc_core_1/sky130_fd_sc_hs__a21oi_1_45/a_29_368# osc_core_1/sky130_fd_sc_hs__nand2_1_5/B
+ osc_core_1/sky130_fd_sc_hs__nand2_2_108/a_27_74# osc_core_1/sky130_fd_sc_hs__nand2_2_79/B
+ osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_1/A osc_core_1/sky130_fd_sc_hs__nand2_2_35/Y
+ osc_core_1/sky130_fd_sc_hs__nand2_2_85/a_27_74# osc_core_1/sky130_fd_sc_hs__nand2_2_13/a_27_74#
+ osc_core_1/sky130_fd_sc_hs__einvp_4_13/a_473_323# osc_core_1/sky130_fd_sc_hs__nand2_4_77/a_27_74#
+ osc_core_1/sky130_fd_sc_hs__nand2_2_1/a_27_74# osc_core_1/sky130_fd_sc_hs__nand2_4_106/a_27_74#
+ osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_49/a_289_74# osc_core_1/sky130_fd_sc_hs__nand2_4_102/Y
+ osc_core_1/sky130_fd_sc_hs__a21oi_1_43/a_117_74# osc_core_1/sky130_fd_sc_hs__bufbuf_8_1/X
+ osc_core_1/sky130_fd_sc_hs__nand2_4_21/a_27_74# osc_core_1/sky130_fd_sc_hs__dfrtp_4_1/a_494_366#
+ osc_core_1/sky130_fd_sc_hs__einvp_8_15/a_27_368# osc_core_1/sky130_fd_sc_hs__einvp_1_17/a_310_392#
+ osc_core_1/sky130_fd_sc_hs__and2_2_3/a_31_74# osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_37/a_405_138#
+ osc_core_1/sky130_fd_sc_hs__nand2_2_65/Y osc_core_1/sky130_fd_sc_hs__nand2_2_37/a_27_74#
+ osc_core_1/sky130_fd_sc_hs__and4_2_1/a_221_74# osc_core_1/sky130_fd_sc_hs__a21oi_1_49/a_29_368#
+ osc_core_1/sky130_fd_sc_hs__clkbuf_2_1/a_43_192# osc_core_1/sky130_fd_sc_hs__einvp_4_1/a_27_368#
+ osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_75/A osc_core_1/sky130_fd_sc_hs__nand2_4_145/a_27_74#
+ osc_core_1/sky130_fd_sc_hs__nand2_4_61/Y osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_21/a_289_74#
+ osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_29/a_28_74# osc_core_1/sky130_fd_sc_hs__a21oi_1_13/a_117_74#
+ osc_core_1/sky130_fd_sc_hs__nand2_2_96/Y osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_31/a_289_74#
+ osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_27/a_405_138# osc_core_1/sky130_fd_sc_hs__nand2_4_60/a_27_74#
+ osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_37/A osc_core_1/sky130_fd_sc_hs__nand2_8_49/a_27_74#
+ osc_core_1/sky130_fd_sc_hs__nand2_4_25/Y osc_core_1/sky130_fd_sc_hs__and4_2_5/a_221_74#
+ osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_7/a_289_74# osc_core_1/sky130_fd_sc_hs__clkbuf_2_5/a_43_192#
+ osc_core_1/sky130_fd_sc_hs__nand2_2_93/a_27_74# osc_core_1/sky130_fd_sc_hs__nand2_4_85/a_27_74#
+ osc_core_1/sky130_fd_sc_hs__nand2_4_15/a_27_74# osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_68/A
+ osc_core_1/sky130_fd_sc_hs__einvp_4_5/a_473_323# osc_core_1/sky130_fd_sc_hs__nand2_4_55/Y
+ osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_17/a_405_138# osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_57/a_405_138#
+ osc_core_1/sky130_fd_sc_hs__inv_1_9/A osc_core_1/sky130_fd_sc_hs__a21oi_1_17/a_117_74#
+ osc_core_1/sky130_fd_sc_hs__nand2_2_89/Y osc_core_1/sky130_fd_sc_hs__einvp_2_17/a_27_368#
+ osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_51/X osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_69/a_289_74#
+ osc_core_1/sky130_fd_sc_hs__einvp_8_8/a_802_323# osc_core_1/sky130_fd_sc_hs__and4_2_3/A
+ osc_core_1/sky130_fd_sc_hs__einvp_8_14/a_27_74# osc_core_1/sky130_fd_sc_hs__dfrtp_4_3/a_699_463#
+ osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_35/a_289_74# osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_3/a_28_74#
+ osc_core_1/sky130_fd_sc_hs__einvp_2_1/a_27_368# osc_core_1/sky130_fd_sc_hs__and4_2_5/C
+ osc_core_1/sky130_fd_sc_hs__nand2_8_17/a_27_74# osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_14/a_28_74#
+ osc_core_1/sky130_fd_sc_hs__conb_1_1/a_21_290# osc_core_1/sky130_fd_sc_hs__nand2_4_139/a_27_74#
+ osc_core_1/sky130_fd_sc_hs__inv_1_1/Y osc_core_1/sky130_fd_sc_hs__clkbuf_2_8/a_43_192#
+ osc_core_1/sky130_fd_sc_hs__einvp_1_1/a_310_392# osc_core_1/sky130_fd_sc_hs__nand2_2_3/Y
+ osc_core_1/sky130_fd_sc_hs__nand2_4_55/a_27_74# osc_core_1/sky130_fd_sc_hs__nand2_2_33/Y
+ osc_core_1/sky130_fd_sc_hs__and4_2_3/a_143_74# osc_core_1/sky130_fd_sc_hs__and4_2_3/B
+ osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_39/a_289_74# osc_core_1/sky130_fd_sc_hs__a21oi_1_33/a_117_74#
+ osc_core_1/sky130_fd_sc_hs__buf_4_1/A osc_core_1/sky130_fd_sc_hs__clkbuf_4_5/a_83_270#
+ osc_core_1/sky130_fd_sc_hs__nand2_2_63/Y osc_core_1/sky130_fd_sc_hs__clkbuf_4_3/A
+ osc_core_1/sky130_fd_sc_hs__a21oi_1_39/a_29_368# osc_core_1/sky130_fd_sc_hs__nand2_4_131/Y
+ osc_core_1/sky130_fd_sc_hs__nand2_4_95/a_27_74# osc_core_1/sky130_fd_sc_hs__nand2_4_123/a_27_74#
+ osc_core_1/sky130_fd_sc_hs__clkbuf_4_5/X osc_core_1/sky130_fd_sc_hs__nand2_4_1/a_27_74#
+ osc_core_1/sky130_fd_sc_hs__clkbuf_1_1/A osc_core_1/sky130_fd_sc_hs__einvp_1_13/a_318_74#
+ osc_core_1/sky130_fd_sc_hs__einvp_8_5/a_27_74# osc_core_1/sky130_fd_sc_hs__a21oi_1_35/a_117_74#
+ osc_core_1/sky130_fd_sc_hs__nand2_1_9/Y osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_53/a_289_74#
+ osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_25/a_405_138# osc_core_1/sky130_fd_sc_hs__nand2_2_55/a_27_74#
+ osc_core_1/sky130_fd_sc_hs__nand2_4_23/Y osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_65/a_405_138#
+ osc_core_1/sky130_fd_sc_hs__nand2_4_49/a_27_74# osc_core_1/sky130_fd_sc_hs__nand2_4_147/a_27_74#
+ osc_core_1/sky130_fd_sc_hs__nand2_8_41/a_27_74# osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_3/A
+ osc_core_1/sky130_fd_sc_hs__and2_2_3/A osc_core_1/sky130_fd_sc_hs__nand2_2_7/B osc_core_1/sky130_fd_sc_hs__nand2_2_19/Y
+ osc_core_1/sky130_fd_sc_hs__einvp_2_17/a_263_323# osc_core_1/sky130_fd_sc_hs__einvp_8_5/a_802_323#
+ osc_core_1/sky130_fd_sc_hs__a21oi_1_21/a_29_368# osc_core_1/sky130_fd_sc_hs__nand2_2_79/a_27_74#
+ osc_core_1/sky130_fd_sc_hs__nand2_4_53/Y osc_core_1/sky130_fd_sc_hs__clkbuf_2_8/A
+ osc_core_1/sky130_fd_sc_hs__and4_2_3/D osc_core_1/sky130_fd_sc_hs__a21oi_1_3/a_29_368#
+ osc_core_1/sky130_fd_sc_hs__einvp_1_17/a_318_74# osc_core_1/sky130_fd_sc_hs__dlygate4sd2_1_1/A
+ osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_56/a_405_138# osc_core_1/sky130_fd_sc_hs__clkbuf_1_1/a_27_74#
+ osc_core_1/sky130_fd_sc_hs__einvp_4_15/a_27_74# osc_core_1/sky130_fd_sc_hs__nand2_8_3/a_27_74#
+ osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_63/a_28_74# osc_core_1/sky130_fd_sc_hs__nand2_2_96/a_27_74#
+ osc_core_1/sky130_fd_sc_hs__nand2_4_89/a_27_74# osc_core_1/sky130_fd_sc_hs__inv_4_13/Y
+ osc_core_1/sky130_fd_sc_hs__nand2_2_49/Y osc_core_1/sky130_fd_sc_hs__einvp_2_1/a_36_74#
+ osc_core_1/sky130_fd_sc_hs__nand2_8_11/a_27_74# osc_core_1/sky130_fd_sc_hs__nand2_2_102/Y
+ osc_core_1/sky130_fd_sc_hs__and2_2_3/B osc_core_1/sky130_fd_sc_hs__dfrtp_4_3/a_124_78#
+ osc_core_1/sky130_fd_sc_hs__nand2_4_83/Y osc_core_1/sky130_fd_sc_hs__and4_2_1/a_56_74#
+ osc_core_1/sky130_fd_sc_hs__nand2_4_33/a_27_74# osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_7/a_28_74#
+ osc_core_1/sky130_fd_sc_hs__nand2_1_3/a_117_74# osc_core_1/sky130_fd_sc_hs__a21oi_1_25/a_29_368#
+ osc_core_1/sky130_fd_sc_hs__nand2_2_31/Y osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_45/a_405_138#
+ osc_core_1/sky130_fd_sc_hs__nand2_2_49/a_27_74# osc_core_1/sky130_fd_sc_hs__a21oi_1_7/a_29_368#
+ osc_core_1/sky130_fd_sc_hs__nand2_2_78/Y osc_core_1/sky130_fd_sc_hs__dlygate4sd2_1_1/a_288_74#
+ osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_31/a_28_74# osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_29/a_289_74#
+ osc_core_1/sky130_fd_sc_hs__clkbuf_2_7/X osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_74/a_289_74#
+ osc_core_1/sky130_fd_sc_hs__nand2_4_157/a_27_74# osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_43/X
+ osc_core_1/sky130_fd_sc_hs__nand2_4_111/Y osc_core_1/sky130_fd_sc_hs__einvp_1_15/a_310_392#
+ osc_core_1/sky130_fd_sc_hs__nand2_4_73/a_27_74# osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_35/a_405_138#
+ osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_75/a_405_138# osc_core_1/sky130_fd_sc_hs__einvp_1_3/a_44_549#
+ osc_core_1/sky130_fd_sc_hs__einvp_4_13/a_27_368# osc_core_1/sky130_fd_sc_hs__nand2_1_7/a_117_74#
+ osc_core_1/sky130_fd_sc_hs__a21oi_1_28/a_29_368# osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_57/a_28_74#
+ osc_core_1/sky130_fd_sc_hs__nand2_4_9/Y osc_core_1/sky130_fd_sc_hs__nand2_2_7/a_27_74#
+ osc_core_1/sky130_fd_sc_hs__dfrtp_4_3/a_1827_81# osc_core_1/sky130_fd_sc_hs__nand2_2_92/Y
+ osc_core_1/sky130_fd_sc_hs__nand2_1_7/Y osc_core_1/sky130_fd_sc_hs__nand2_2_33/a_27_74#
+ osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_33/A osc_core_1/sky130_fd_sc_hs__nand2_2_65/B
+ osc_core_1/sky130_fd_sc_hs__nand2_4_21/Y osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_1/a_405_138#
+ osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_11/a_289_74# osc_core_1/sky130_fd_sc_hs__nand2_4_69/Y
+ osc_core_1/sky130_fd_sc_hs__and2_2_3/a_118_74# osc_core_1/sky130_fd_sc_hs__and4_2_1/X
+ osc_core_1/sky130_fd_sc_hs__nand2_4_41/a_27_74# osc_core_1/sky130_fd_sc_hs__einvp_1_7/a_44_549#
+ osc_core_1/sky130_fd_sc_hs__nand2_4_141/a_27_74# osc_core_1/sky130_fd_sc_hs__nand2_4_121/Y
+ osc_core_1/sky130_fd_sc_hs__nand2_2_17/Y osc_core_1/sky130_fd_sc_hs__einvp_8_7/a_27_368#
+ osc_core_1/sky130_fd_sc_hs__einvp_2_15/a_263_323# osc_core_1/sky130_fd_sc_hs__a21oi_1_11/a_29_368#
+ osc_core_1/sky130_fd_sc_hs__nand2_8_45/a_27_74# osc_core_1/sky130_fd_sc_hs__einvp_2_7/a_263_323#
+ osc_core_1/sky130_fd_sc_hs__nand2_4_99/Y osc_core_1/sky130_fd_sc_hs__nand2_4_67/a_27_74#
+ osc_core_1/sky130_fd_sc_hs__a21oi_1_29/a_117_74# osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_3/X
+ osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_53/a_405_138# osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_47/a_289_74#
+ osc_core_1/sky130_fd_sc_hs__nand2_2_73/B osc_core_1/sky130_fd_sc_hs__dfrtp_4_1/a_699_463#
+ osc_core_1/sky130_fd_sc_hs__a21oi_1_42/a_117_74# osc_core_1/sky130_fd_sc_hs__nand2_2_47/Y
+ osc_core_1/sky130_fd_sc_hs__nand2_4_11/a_27_74# osc_core_1/sky130_fd_sc_hs__nand2_4_81/Y
+ osc_core_1/sky130_fd_sc_hs__nand2_4_115/Y osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_65/a_28_74#
+ osc_core_1/sky130_fd_sc_hs__nand2_2_27/a_27_74# osc_core_1/sky130_fd_sc_hs__einvp_8_8/a_27_74#
+ osc_core_1/sky130_fd_sc_hs__nand2_4_119/a_27_74# osc_core_1/sky130_fd_sc_hs__nand2_4_43/Y
+ osc_core_1/sky130_fd_sc_hs__einvp_2_3/a_36_74# osc_core_1/sky130_fd_sc_hs__a21oi_1_15/a_29_368#
+ osc_core_1/sky130_fd_sc_hs__nand2_8_13/a_27_74# osc_core_1/sky130_fd_sc_hs__and4_2_3/a_56_74#
+ osc_core_1/sky130_fd_sc_hs__nand2_2_43/a_27_74# osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_20/A
+ osc_core_1/sky130_fd_sc_hs__nand2_4_35/a_27_74# osc_core_1/sky130_fd_sc_hs__nand2_2_37/B
+ osc_core_1/sky130_fd_sc_hs__einvp_4_11/a_473_323# osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_9/X
+ osc_core_1/sky130_fd_sc_hs__and4_2_5/B osc_core_1/sky130_fd_sc_hs__nand2_4_145/Y
+ osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_20/a_289_74# osc_core_1/sky130_fd_sc_hs__a21oi_1_45/a_117_74#
+ osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_20/a_28_74# osc_core_1/sky130_fd_sc_hs__clkbuf_2_17/a_43_192#
+ osc_core_1/sky130_fd_sc_hs__nand3_4_3/C osc_core_1/sky130_fd_sc_hs__dfrtp_4_3/a_789_463#
+ osc_core_1/sky130_fd_sc_hs__einvp_8_17/a_27_368# osc_core_1/sky130_fd_sc_hs__nand2_8_39/a_27_74#
+ osc_core_1/sky130_fd_sc_hs__bufbuf_8_1/a_221_368# osc_core_1/sky130_fd_sc_hs__and4_2_3/a_221_74#
+ osc_core_1/sky130_fd_sc_hs__nand2_2_67/a_27_74# osc_core_1/sky130_fd_sc_hs__einvp_4_9/a_27_74#
+ osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_74/a_405_138# osc_core_1/sky130_fd_sc_hs__nand2_2_21/Y
+ osc_core_1/sky130_fd_sc_hs__nand2_4_159/a_27_74# osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_5/a_289_74#
+ osc_core_1/sky130_fd_sc_hs__nand2_4_39/Y osc_core_1/sky130_fd_sc_hs__nand2_4_7/Y
+ osc_core_1/sky130_fd_sc_hs__a21oi_1_19/a_29_368# osc_core_1/sky130_fd_sc_hs__nand2_2_105/a_27_74#
+ osc_core_1/sky130_fd_sc_hs__nand2_2_12/a_27_74# osc_core_1/sky130_fd_sc_hs__nand2_2_84/a_27_74#
+ osc_core_1/sky130_fd_sc_hs__nand2_1_5/Y osc_core_1/sky130_fd_sc_hs__nand2_4_103/a_27_74#
+ osc_core_1/sky130_fd_sc_hs__a21oi_1_49/a_117_74# osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_59/a_28_74#
+ osc_core_1/sky130_fd_sc_hs__einvp_2_15/a_27_368# osc_core_1/sky130_fd_sc_hs__dfrtp_4_1/a_313_74#
+ osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_68/a_289_74# osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_79/X
+ osc_core_1/sky130_fd_sc_hs__inv_1_7/A osc_core_1/sky130_fd_sc_hs__nand2_4_91/a_27_74#
+ osc_core_1/sky130_fd_sc_hs__nand2_4_67/Y osc_core_1/sky130_fd_sc_hs__inv_4_27/Y
+ osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_75/a_28_74# osc_core_1/sky130_fd_sc_hs__clkbuf_4_1/a_83_270#
+ osc_core_1/sky130_fd_sc_hs__einvp_8_3/a_27_74# osc_core_1/sky130_fd_sc_hs__nand2_4_129/a_27_74#
+ osc_core_1/sky130_fd_sc_hs__nand2_8_23/a_27_74# osc_core_1/sky130_fd_sc_hs__nand2_4_7/a_27_74#
+ osc_core_1/sky130_fd_sc_hs__einvp_4_7/a_27_368# osc_core_1/sky130_fd_sc_hs__nand2_2_51/a_27_74#
+ osc_core_1/sky130_fd_sc_hs__dfrtp_4_3/a_834_355# osc_core_1/sky130_fd_sc_hs__nand2_4_45/a_27_74#
+ osc_core_1/sky130_fd_sc_hs__nand2_2_84/Y osc_core_1/sky130_fd_sc_hs__nand2_4_97/Y
+ osc_core_1/sky130_fd_sc_hs__einvp_2_5/a_263_323# osc_core_1/sky130_fd_sc_hs__einvp_4_3/a_473_323#
+ osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_15/a_405_138# osc_core_1/sky130_fd_sc_hs__dfrtp_4_3/a_1627_493#
+ osc_core_1/sky130_fd_sc_hs__einvp_2_19/a_27_368# osc_core_1/sky130_fd_sc_hs__einvp_8_19/a_802_323#
+ osc_core_1/sky130_fd_sc_hs__nand2_2_45/Y osc_core_1/sky130_fd_sc_hs__einvp_2_3/a_27_368#
+ osc_core_1/sky130_fd_sc_hs__dfrtp_4_3/a_812_138# osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_43/a_28_74#
+ osc_core_1/sky130_fd_sc_hs__nand2_4_113/Y osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_53/A
+ osc_core_1/sky130_fd_sc_hs__einvp_4_11/a_27_74# osc_core_1/sky130_fd_sc_hs__nand2_4_41/Y
+ osc_core_1/sky130_fd_sc_hs__nand2_2_92/a_27_74# osc_core_1/sky130_fd_sc_hs__nand2_2_109/Y
+ osc_core_1/sky130_fd_sc_hs__einvp_1_9/a_310_392# osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_43/a_405_138#
+ osc_core_1/sky130_fd_sc_hs__nand2_4_113/a_27_74# osc_core_1/sky130_fd_sc_hs__clkbuf_2_1/X
+ osc_core_1/sky130_fd_sc_hs__nand2_8_9/a_27_74# osc_core_1/sky130_fd_sc_hs__nand2_2_35/B
+ osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_69/a_28_74# osc_core_1/sky130_fd_sc_hs__nand2_2_7/Y
+ osc_core_1/sky130_fd_sc_hs__nand2_4_143/Y osc_core_1/sky130_fd_sc_hs__einvp_8_15/a_27_74#
+ osc_core_1/sky130_fd_sc_hs__einvp_2_7/a_36_74# osc_core_1/sky130_fd_sc_hs__dfrtp_4_3/a_37_78#
+ osc_core_1/sky130_fd_sc_hs__nand2_4_107/Y osc_core_1/sky130_fd_sc_hs__nand2_2_45/a_27_74#
+ osc_core_1/sky130_fd_sc_hs__einvp_1_13/a_310_392# osc_core_1/sky130_fd_sc_hs__dfrtp_4_1/a_1627_493#
+ osc_core_1/sky130_fd_sc_hs__einvp_1_1/a_318_74# osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_33/a_405_138#
+ osc_core_1/sky130_fd_sc_hs__nand2_4_5/Y osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_71/a_405_138#
+ osc_core_1/sky130_fd_sc_hs__einvp_4_3/a_27_74# osc_core_1/sky130_fd_sc_hs__nand2_4_153/a_27_74#
+ osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_37/a_28_74# osc_core_1/sky130_fd_sc_hs__nand2_1_3/Y
+ osc_core_1/sky130_fd_sc_hs__nand2_4_135/Y osc_core_1/sky130_fd_sc_hs__dfrtp_4_1/a_1827_81#
+ osc_core_1/sky130_fd_sc_hs__a21oi_1_39/a_117_74# osc_core_1/sky130_fd_sc_hs__einvp_2_11/a_36_74#
+ osc_core_1/sky130_fd_sc_hs__inv_1_5/A osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_51/a_28_74#
+ osc_core_1/sky130_fd_sc_hs__nand2_4_65/Y osc_core_1/sky130_fd_sc_hs__nand2_4_79/a_27_74#
+ osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_23/a_405_138# osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_63/a_405_138#
+ osc_core_1/sky130_fd_sc_hs__einvp_1_5/a_318_74# osc_core_1/sky130_fd_sc_hs__nand2_4_27/Y
+ osc_core_1/sky130_fd_sc_hs__nand2_4_23/a_27_74# osc_core_1/sky130_fd_sc_hs__nand2_4_121/a_27_74#
+ osc_core_1/sky130_fd_sc_hs__einvp_2_13/a_263_323# osc_core_1/sky130_fd_sc_hs__nand2_4_129/Y
+ osc_core_1/sky130_fd_sc_hs__nand2_2_39/a_27_74# osc_core_1/sky130_fd_sc_hs__nand2_4_95/Y
+ osc_core_1/sky130_fd_sc_hs__clkbuf_2_17/A osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_14/a_405_138#
+ osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_51/a_405_138# osc_core_1/sky130_fd_sc_hs__einvp_1_13/a_44_549#
+ osc_core_1/sky130_fd_sc_hs__a21oi_1_21/a_117_74# osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_71/a_289_74#
+ osc_core_1/sky130_fd_sc_hs__a21oi_1_3/a_117_74# osc_core_1/sky130_fd_sc_hs__einvp_1_9/a_318_74#
+ osc_core_1/sky130_fd_sc_hs__conb_1_1/a_165_290# osc_core_1/sky130_fd_sc_hs__nand2_4_63/a_27_74#
+ osc_core_1/sky130_fd_sc_hs__nand2_2_105/Y osc_core_1/sky130_fd_sc_hs__and4_2_1/a_335_74#
+ osc_core_1/sky130_fd_sc_hs__nand2_2_78/a_27_74# osc_core_1/sky130_fd_sc_hs__nand2_2_5/Y
+ osc_core_1/sky130_fd_sc_hs__nand2_4_141/Y osc_core_1/sky130_fd_sc_hs__dfrtp_4_3/a_1678_395#
+ osc_core_1/sky130_fd_sc_hs__einvp_1_17/a_44_549# osc_core_1/sky130_fd_sc_hs__einvp_4_13/a_27_74#
+ osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_62/a_28_74# osc_core_1/sky130_fd_sc_hs__nand2_2_23/a_27_74#
+ osc_core_1/sky130_fd_sc_hs__nand3_4_1/a_456_82# osc_core_1/sky130_fd_sc_hs__a21oi_1_25/a_117_74#
+ osc_core_1/sky130_fd_sc_hs__nand2_4_17/a_27_74# osc_core_1/sky130_fd_sc_hs__nand2_4_103/Y
+ osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_43/a_289_74# osc_core_1/sky130_fd_sc_hs__dfrtp_4_1/a_789_463#
+ osc_core_1/sky130_fd_sc_hs__a21oi_1_7/a_117_74# osc_core_1/sky130_fd_sc_hs__einvp_8_17/a_27_74#
+ osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_5/a_28_74# osc_core_1/sky130_fd_sc_hs__nand2_4_3/Y
+ osc_core_1/sky130_fd_sc_hs__nand2_4_33/Y osc_core_1/sky130_fd_sc_hs__einvp_2_9/a_36_74#
+ osc_core_1/sky130_fd_sc_hs__einvp_4_17/a_27_368# osc_core_1/sky130_fd_sc_hs__nand2_4_131/a_27_74#
+ osc_core_1/sky130_fd_sc_hs__and4_2_5/a_335_74# osc_core_1/sky130_fd_sc_hs__nand2_1_1/Y
+ osc_core_1/sky130_fd_sc_hs__clkbuf_4_5/A osc_core_1/sky130_fd_sc_hs__nand2_4_133/Y
+ osc_core_1/sky130_fd_sc_hs__nand2_8_35/a_27_74# osc_core_1/sky130_fd_sc_hs__nand2_2_29/Y
+ osc_core_1/sky130_fd_sc_hs__dlygate4sd2_1_1/a_405_138# osc_core_1/sky130_fd_sc_hs__nand2_2_63/a_27_74#
+ osc_core_1/sky130_fd_sc_hs__a21oi_1_28/a_117_74# osc_core_1/sky130_fd_sc_hs__einvp_4_5/a_27_74#
+ osc_core_1/sky130_fd_sc_hs__nand2_4_57/a_27_74# osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_79/a_289_74#
+ osc_core_1/sky130_fd_sc_hs__nand2_4_63/Y osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_9/a_405_138#
+ osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_15/a_289_74# osc_core_1/sky130_fd_sc_hs__nand2_2_97/Y
+ osc_core_1/sky130_fd_sc_hs__nand2_2_103/a_27_74# osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_62/a_405_138#
+ osc_core_1/sky130_fd_sc_hs__nand2_2_12/Y osc_core_1/sky130_fd_sc_hs__einvp_2_13/a_36_74#
+ osc_core_1/sky130_fd_sc_hs__dfrtp_4_1/a_1678_395# osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_56/a_28_74#
+ osc_core_1/sky130_fd_sc_hs__bufbuf_8_1/a_334_368# osc_core_1/sky130_fd_sc_hs__nand2_2_17/a_27_74#
+ osc_core_1/sky130_fd_sc_hs__nand2_2_89/a_27_74# osc_core_1/sky130_fd_sc_hs__nand2_4_111/a_27_74#
+ osc_core_1/sky130_fd_sc_hs__a21oi_1_47/a_29_368# osc_core_1/sky130_fd_sc_hs__nand2_4_127/Y
+ osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_1/a_289_74# osc_core_1/sky130_fd_sc_hs__nand2_4_93/Y
+ osc_core_1/sky130_fd_sc_hs__einvp_8_3/a_802_323# osc_core_1/sky130_fd_sc_hs__dfrtp_4_1/a_834_355#
+ osc_core_1/sky130_fd_sc_hs__einvp_2_3/a_263_323# osc_core_1/sky130_fd_sc_hs__einvp_4_1/a_473_323#
+ osc_core_1/sky130_fd_sc_hs__nand2_4_97/a_27_74# osc_core_1/sky130_fd_sc_hs__nand2_2_42/Y
+ osc_core_1/sky130_fd_sc_hs__nand2_4_125/a_27_74# osc_core_1/sky130_fd_sc_hs__nand2_4_3/a_27_74#
+ osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_79/a_28_74# osc_core_1/sky130_fd_sc_hs__einvp_8_17/a_802_323#
+ osc_core_1/sky130_fd_sc_hs__a21oi_1_11/a_117_74# osc_core_1/sky130_fd_sc_hs__and4_2_5/A
+ osc_core_1/sky130_fd_sc_hs__einvp_2_11/a_27_368# osc_core_1/sky130_fd_sc_hs__clkbuf_2_15/a_43_192#
+ osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_63/a_289_74# osc_core_1/sky130_fd_sc_hs__dfrtp_4_1/a_812_138#
+ osc_core_1/sky130_fd_sc_hs__einvp_8_7/a_27_74# osc_core_1/sky130_fd_sc_hs__nand2_4_157/Y
+ osc_core_1/sky130_fd_sc_hs__nand2_4_19/Y osc_core_1/sky130_fd_sc_hs__nand2_8_29/a_27_74#
+ osc_core_1/sky130_fd_sc_hs__nand2_2_57/a_27_74# osc_core_1/sky130_fd_sc_hs__nand3_4_1/a_27_82#
+ osc_core_1/sky130_fd_sc_hs__nand2_2_71/Y osc_core_1/sky130_fd_sc_hs__nand2_4_149/a_27_74#
+ osc_core_1/sky130_fd_sc_hs__nand2_4_119/Y osc_core_1/sky130_fd_sc_hs__nand2_4_85/Y
+ osc_core_1/sky130_fd_sc_hs__clkbuf_2_3/a_43_192# osc_core_1/sky130_fd_sc_hs__einvp_1_7/a_310_392#
+ osc_core_1/sky130_fd_sc_hs__einvp_4_3/a_27_368# osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_41/a_405_138#
+ osc_core_1/sky130_fd_sc_hs__dfrtp_4_3/a_1350_392# osc_core_1/sky130_fd_sc_hs__nand2_4_49/Y
+ osc_core_1/sky130_fd_sc_hs__einvp_4_19/a_473_323# osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_49/a_28_74#
+ osc_core_1/sky130_fd_sc_hs__a21oi_1_15/a_117_74# osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_33/a_289_74#
+ osc_core_1/sky130_fd_sc_hs__nand2_4_81/a_27_74# osc_core_1/sky130_fd_sc_hs__nand2_4_149/Y
+ osc_core_1/sky130_fd_sc_hs__einvp_4_17/a_27_74# osc_core_1/sky130_fd_sc_hs__nand2_8_5/a_27_74#
+ osc_core_1/sky130_fd_sc_hs__nand2_4_1/Y osc_core_1/sky130_fd_sc_hs__nand2_4_31/Y
+ osc_core_1/sky130_fd_sc_hs__einvp_1_11/a_310_392# osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_31/a_405_138#
+ osc_core_1/sky130_fd_sc_hs__nand2_4_79/Y osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_9/a_289_74#
+ osc_core_1/sky130_fd_sc_hs__clkbuf_2_7/a_43_192# osc_core_1/sky130_fd_sc_hs__a21oi_1_32/a_29_368#
+ osc_core_1/sky130_fd_sc_hs__nand2_2_42/a_27_74# osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_9/a_28_74#
+ osc_core_1/sky130_fd_sc_hs__nand2_2_27/Y osc_core_1/sky130_fd_sc_hs__nand2_4_133/a_27_74#
+ osc_core_1/sky130_fd_sc_hs__nand2_1_7/B osc_core_1/sky130_fd_sc_hs__nand2_4_60/Y
+ osc_core_1/sky130_fd_sc_hs__a21oi_1_19/a_117_74# osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_37/a_289_74#
+ osc_core_1/sky130_fd_sc_hs__dfrtp_4_1/a_1350_392# osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_33/a_28_74#
+ osc_core_1/sky130_fd_sc_hs__nand2_2_57/Y osc_core_1/sky130_fd_sc_hs__nand2_4_125/Y
+ osc_core_1/sky130_fd_sc_hs__nand2_4_91/Y osc_core_1/sky130_fd_sc_hs__a21oi_1_37/a_29_368#
+ osc_core_1/sky130_fd_sc_hs__nand2_2_83/a_27_74# osc_core_1/sky130_fd_sc_hs__nand2_4_75/a_27_74#
+ osc_core_1/sky130_fd_sc_hs__einvp_8_2/a_802_323# osc_core_1/sky130_fd_sc_hs__einvp_2_17/a_36_74#
+ osc_core_1/sky130_fd_sc_hs__nand2_4_102/a_27_74# osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_11/a_405_138#
+ osc_core_1/sky130_fd_sc_hs__einvp_1_11/a_318_74# osc_core_1/sky130_fd_sc_hs__nand2_2_88/Y
+ osc_core_1/sky130_fd_sc_hs__einvp_2_7/a_27_368# osc_core_1/sky130_fd_sc_hs__and2_2_1/a_31_74#
+ osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_51/a_289_74# osc_core_1/sky130_fd_sc_hs__nand2_4_17/Y
+ osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_74/a_28_74# osc_core_1/sky130_fd_sc_hs__nand2_4_155/Y
+ osc_core_1/sky130_fd_sc_hs__nand2_2_35/a_27_74# osc_core_1/sky130_fd_sc_hs__nand2_4_29/a_27_74#
+ osc_core_1/sky130_fd_sc_hs__einvp_8_2/a_27_74# osc_core_1/sky130_fd_sc_hs__nand2_2_103/Y
+ osc_core_1/sky130_fd_sc_hs__nand2_8_21/a_27_74# osc_core_1/sky130_fd_sc_hs__nand2_4_117/Y
+ osc_core_1/sky130_fd_sc_hs__nand2_2_1/Y osc_core_1/sky130_fd_sc_hs__nand2_4_43/a_27_74#
+ osc_core_1/sky130_fd_sc_hs__nand2_4_143/a_27_74# osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_27/a_28_74#
+ osc_core_1/sky130_fd_sc_hs__nand2_4_47/Y osc_core_1/sky130_fd_sc_hs__nand2_2_59/a_27_74#
+ osc_core_1/sky130_fd_sc_hs__einvp_1_15/a_318_74# osc_core_1/sky130_fd_sc_hs__a21oi_1_1/a_29_368#
+ osc_core_1/sky130_fd_sc_hs__nand2_2_79/Y osc_core_1/sky130_fd_sc_hs__nand2_8_47/a_27_74#
+ osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_57/a_289_74# osc_core_1/sky130_fd_sc_hs__bufbuf_8_1/a_27_112#
+ osc_core_1/sky130_fd_sc_hs__nand2_4_147/Y osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_23/a_289_74#
+ osc_core_1/sky130_fd_sc_hs__nand2_4_69/a_27_74# osc_core_1/sky130_fd_sc_hs__nand2_2_61/Y
+ osc_core_1/sky130_fd_sc_hs__nand2_4_77/Y osc_core_1/sky130_fd_sc_hs__dfrtp_4_1/a_124_78#
+ osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_79/a_405_138# osc_core_1/sky130_fd_sc_hs__nand2_4_13/a_27_74#
+ osc_core_1/sky130_fd_sc_hs__nand2_2_25/Y osc_core_1/sky130_fd_sc_hs__nand2_1_1/a_117_74#
+ osc_core_1/sky130_fd_sc_hs__dlygate4sd3_1_68/a_28_74# osc_core_1/sky130_fd_sc_hs__a21oi_1_23/a_29_368#
+ osc_core_1/sky130_fd_sc_hs__nand2_2_29/a_27_74# osc_core_1/sky130_fd_sc_hs__einvp_1_19/a_318_74#
+ osc_core_1/sky130_fd_sc_hs__a21oi_1_5/a_29_368# osc_core_1/sky130_fd_sc_hs__dfrtp_4_3/a_1647_81#
+ osc_core
Xsky130_fd_sc_hs__einvp_2_130 DVSS: DVDD: DVDD: DVSS: dout_n sky130_fd_sc_hs__buf_8_1/X
+ sky130_fd_sc_hs__dlrtp_1_127/Q sky130_fd_sc_hs__einvp_2_131/a_263_323# sky130_fd_sc_hs__einvp_2_131/a_36_74#
+ sky130_fd_sc_hs__einvp_2_131/a_27_368# sky130_fd_sc_hs__einvp_2
Xsky130_fd_sc_hs__einvp_2_141 DVSS: DVDD: DVDD: DVSS: dout_p sky130_fd_sc_hs__einvp_2_99/A
+ sky130_fd_sc_hs__dlrtp_1_143/Q sky130_fd_sc_hs__einvp_2_141/a_263_323# sky130_fd_sc_hs__einvp_2_141/a_36_74#
+ sky130_fd_sc_hs__einvp_2_141/a_27_368# sky130_fd_sc_hs__einvp_2
Xsky130_fd_sc_hs__einvp_2_152 DVSS: DVDD: DVDD: DVSS: dout_p sky130_fd_sc_hs__einvp_2_99/A
+ sky130_fd_sc_hs__dlrtp_1_157/Q sky130_fd_sc_hs__einvp_2_153/a_263_323# sky130_fd_sc_hs__einvp_2_153/a_36_74#
+ sky130_fd_sc_hs__einvp_2_153/a_27_368# sky130_fd_sc_hs__einvp_2
Xsky130_fd_sc_hs__clkbuf_16_13 DVSS: DVDD: DVDD: DVSS: osc_core_1/pi1_l[1] sky130_fd_sc_hs__clkbuf_4_19/X
+ sky130_fd_sc_hs__clkbuf_16_13/a_114_74# sky130_fd_sc_hs__clkbuf_16
Xsky130_fd_sc_hs__clkbuf_16_24 DVSS: DVDD: DVDD: DVSS: osc_core_1/pi3_l[3] sky130_fd_sc_hs__clkbuf_8_11/X
+ sky130_fd_sc_hs__clkbuf_16_25/a_114_74# sky130_fd_sc_hs__clkbuf_16
Xsky130_fd_sc_hs__clkbuf_16_35 DVSS: DVDD: DVDD: DVSS: osc_core_1/pi3_l[1] sky130_fd_sc_hs__clkbuf_8_9/X
+ sky130_fd_sc_hs__clkbuf_16_35/a_114_74# sky130_fd_sc_hs__clkbuf_16
Xsky130_fd_sc_hs__clkbuf_16_46 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__buf_8_1/A
+ sky130_fd_sc_hs__nand2_2_1/Y sky130_fd_sc_hs__clkbuf_16_47/a_114_74# sky130_fd_sc_hs__clkbuf_16
Xsky130_fd_sc_hs__clkbuf_16_57 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__buf_2_3/A
+ sky130_fd_sc_hs__einvp_8_3/Z sky130_fd_sc_hs__clkbuf_16_57/a_114_74# sky130_fd_sc_hs__clkbuf_16
Xsky130_fd_sc_hs__clkbuf_16_68 DVSS: DVDD: DVDD: DVSS: qr_4t1_mux_top_1/rst qr_4t1_mux_top_3/rst
+ sky130_fd_sc_hs__clkbuf_16_69/a_114_74# sky130_fd_sc_hs__clkbuf_16
Xsky130_fd_sc_hs__clkbuf_16_79 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__nor4_2_1/B
+ sky130_fd_sc_hs__clkbuf_8_81/X sky130_fd_sc_hs__clkbuf_16_79/a_114_74# sky130_fd_sc_hs__clkbuf_16
Xsky130_fd_sc_hs__clkbuf_16_101 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__clkbuf_8_71/A
+ sky130_fd_sc_hs__clkbuf_8_95/X sky130_fd_sc_hs__clkbuf_16_101/a_114_74# sky130_fd_sc_hs__clkbuf_16
Xsky130_fd_sc_hs__clkbuf_16_112 DVSS: DVDD: DVDD: DVSS: prbs_generator_syn_31/inj_err
+ prbs_generator_syn_27/inj_err sky130_fd_sc_hs__clkbuf_16_113/a_114_74# sky130_fd_sc_hs__clkbuf_16
Xsky130_fd_sc_hs__clkbuf_16_123 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__clkbuf_8_59/A
+ sky130_fd_sc_hs__clkbuf_8_99/X sky130_fd_sc_hs__clkbuf_16_123/a_114_74# sky130_fd_sc_hs__clkbuf_16
Xprbs_generator_syn_9 prbs_generator_syn_9/clk prbs_generator_syn_9/rst prbs_generator_syn_9/cke
+ sky130_fd_sc_hs__conb_1_85/LO sky130_fd_sc_hs__conb_1_85/LO sky130_fd_sc_hs__conb_1_85/HI
+ sky130_fd_sc_hs__conb_1_85/HI sky130_fd_sc_hs__conb_1_85/HI prbs_generator_syn_11/eqn[9]
+ sky130_fd_sc_hs__conb_1_85/LO sky130_fd_sc_hs__conb_1_85/HI sky130_fd_sc_hs__conb_1_85/HI
+ sky130_fd_sc_hs__conb_1_85/HI sky130_fd_sc_hs__conb_1_85/HI prbs_generator_syn_9/cke
+ prbs_generator_syn_9/cke prbs_generator_syn_9/eqn[31] prbs_generator_syn_9/cke prbs_generator_syn_9/cke
+ prbs_generator_syn_9/cke prbs_generator_syn_9/cke prbs_generator_syn_9/eqn[1] prbs_generator_syn_9/eqn[1]
+ prbs_generator_syn_9/eqn[1] prbs_generator_syn_9/eqn[1] prbs_generator_syn_9/eqn[1]
+ prbs_generator_syn_9/eqn[2] sky130_fd_sc_hs__conb_1_83/LO sky130_fd_sc_hs__conb_1_83/HI
+ sky130_fd_sc_hs__conb_1_83/LO sky130_fd_sc_hs__conb_1_83/HI sky130_fd_sc_hs__conb_1_83/HI
+ sky130_fd_sc_hs__conb_1_83/LO sky130_fd_sc_hs__conb_1_83/LO sky130_fd_sc_hs__conb_1_83/HI
+ prbs_generator_syn_9/eqn[31] prbs_generator_syn_9/eqn[30] prbs_generator_syn_9/eqn[30]
+ prbs_generator_syn_9/eqn[28] prbs_generator_syn_9/eqn[28] prbs_generator_syn_9/eqn[28]
+ prbs_generator_syn_9/eqn[28] prbs_generator_syn_9/eqn[28] prbs_generator_syn_9/eqn[28]
+ prbs_generator_syn_9/eqn[22] prbs_generator_syn_9/eqn[22] prbs_generator_syn_9/eqn[20]
+ prbs_generator_syn_9/eqn[22] prbs_generator_syn_9/eqn[22] prbs_generator_syn_9/eqn[22]
+ prbs_generator_syn_9/eqn[16] prbs_generator_syn_9/eqn[16] prbs_generator_syn_9/eqn[16]
+ prbs_generator_syn_3/eqn[4] prbs_generator_syn_9/eqn[16] prbs_generator_syn_9/eqn[16]
+ prbs_generator_syn_9/eqn[16] prbs_generator_syn_9/eqn[9] prbs_generator_syn_9/eqn[9]
+ prbs_generator_syn_9/eqn[9] prbs_generator_syn_9/eqn[9] prbs_generator_syn_9/eqn[9]
+ prbs_generator_syn_9/eqn[9] prbs_generator_syn_9/eqn[9] prbs_generator_syn_9/eqn[2]
+ prbs_generator_syn_9/eqn[1] prbs_generator_syn_9/eqn[2] prbs_generator_syn_9/inj_err
+ prbs_generator_syn_9/eqn[31] prbs_generator_syn_9/eqn[31] prbs_generator_syn_9/out
+ DVSS: DVDD: prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_1/a_293_74# prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_15/X
+ prbs_generator_syn_9/sky130_fd_sc_hs__nand2_1_35/B prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_51/Y
+ prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_9/A prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_9/CLK
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_47/a_27_74# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_37/a_1226_296#
+ prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_3/B prbs_generator_syn_9/sky130_fd_sc_hs__nor2b_1_7/a_27_112#
+ prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_29/B prbs_generator_syn_9/sky130_fd_sc_hs__sdlclkp_2_1/a_580_74#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_1/a_1141_508# prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_5/Y
+ prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_41/a_230_79# prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_61/a_138_385#
+ prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_43/a_132_392# prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_3/a_222_392#
+ prbs_generator_syn_9/sky130_fd_sc_hs__nor2b_1_9/a_27_112# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_61/a_27_74#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_35/a_206_368# prbs_generator_syn_9/sky130_fd_sc_hs__nand2_2_3/Y
+ prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_25/B prbs_generator_syn_9/sky130_fd_sc_hs__nand2_1_11/a_117_74#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_67/a_651_503# prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_45/X
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_39/a_696_458# prbs_generator_syn_9/sky130_fd_sc_hs__sdlclkp_2_1/a_1198_74#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_45/a_1034_424# prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_17/a_222_392#
+ prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_55/a_222_392# prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_53/Y
+ prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_35/A prbs_generator_syn_9/m3_13600_1651#
+ prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_59/a_52_123# prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_5/a_293_74#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_35/a_1226_296# prbs_generator_syn_9/sky130_fd_sc_hs__nand2_1_51/B
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_5/a_651_503# prbs_generator_syn_9/sky130_fd_sc_hs__nand2_1_21/B
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_8/a_27_74# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_15/a_27_74#
+ prbs_generator_syn_9/sky130_fd_sc_hs__and2b_2_1/X prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_13/X
+ prbs_generator_syn_9/sky130_fd_sc_hs__nand2_2_3/a_27_74# prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_50/a_138_385#
+ prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_33/a_132_392# prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_1/a_376_368#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_25/a_206_368# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_35/a_437_503#
+ prbs_generator_syn_9/sky130_fd_sc_hs__sdlclkp_2_1/a_708_451# prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_45/a_230_79#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_29/a_696_458# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_32/a_27_74#
+ prbs_generator_syn_9/sky130_fd_sc_hs__nor2b_1_4/Y prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_59/a_293_74#
+ prbs_generator_syn_9/sky130_fd_sc_hs__nand2_1_47/a_117_74# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_73/a_735_102#
+ prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_21/a_112_119# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_23/a_1141_508#
+ prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_25/a_293_74# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_7/Q
+ prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_3/a_112_119# prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_35/B
+ prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_51/X prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_53/a_1178_124#
+ prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_23/a_132_392# prbs_generator_syn_9/sky130_fd_sc_hs__nand2_1_3/B
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_15/a_206_368# prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_63/a_132_392#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_55/a_27_74# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_25/a_437_503#
+ prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_41/a_52_123# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_47/a_651_503#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_73/a_1141_508# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_19/a_696_458#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_57/a_696_458# prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_7/X
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_43/a_1034_424# prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_55/A
+ prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_11/a_112_119# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_21/a_1141_508#
+ prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_35/a_222_392# prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_49/a_230_79#
+ prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_67/Y prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_71/a_27_74#
+ prbs_generator_syn_9/sky130_fd_sc_hs__nand2_1_33/B prbs_generator_syn_9/sky130_fd_sc_hs__conb_1_1/LO
+ prbs_generator_syn_9/sky130_fd_sc_hs__nand2_1_19/a_117_74# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_51/a_1178_124#
+ prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_33/X prbs_generator_syn_9/sky130_fd_sc_hs__nand2_1_29/B
+ prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_41/Y prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_53/a_132_392#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_45/a_206_368# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_15/a_437_503#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_37/a_651_503# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_39/a_544_485#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_53/a_735_102# prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_45/a_52_123#
+ prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_1/B prbs_generator_syn_9/sky130_fd_sc_hs__nand2_2_3/B
+ prbs_generator_syn_9/sky130_fd_sc_hs__clkbuf_16_1/A prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_21/X
+ prbs_generator_syn_9/sky130_fd_sc_hs__nand2_1_25/B prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_39/a_376_368#
+ prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_63/X prbs_generator_syn_9/m3_13600_3481#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_69/a_1178_124# prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_21/a_138_385#
+ prbs_generator_syn_9/sky130_fd_sc_hs__nor2b_1_8/Y prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_19/a_1178_124#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_49/a_27_74# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_45/a_437_503#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_27/a_651_503# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_71/a_1141_508#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_65/a_651_503# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_29/a_544_485#
+ prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_3/a_138_385# prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_55/X
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_43/a_735_102# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_41/a_1034_424#
+ prbs_generator_syn_9/sky130_fd_sc_hs__nand2_1_9/B prbs_generator_syn_9/sky130_fd_sc_hs__nor2b_1_9/Y
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_59/a_1034_424# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_39/a_1141_508#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_33/a_1226_296# prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_49/a_52_123#
+ prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_47/Y prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_43/Y
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_4/a_651_503# prbs_generator_syn_9/sky130_fd_sc_hs__nand2_1_49/B
+ prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_19/A prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_11/a_138_385#
+ prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_5/X prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_63/a_206_368#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_17/a_651_503# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_19/a_544_485#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_55/a_651_503# prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_9/Y
+ prbs_generator_syn_9/sky130_fd_sc_hs__nand2_1_17/B prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_57/a_544_485#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_67/a_696_458# prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_35/X
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_19/a_27_74# prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_45/a_222_392#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_32/a_1226_296# prbs_generator_syn_9/sky130_fd_sc_hs__nand2_1_43/B
+ prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_25/A prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_1/a_206_368#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_49/a_1226_296# prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_1/a_112_119#
+ prbs_generator_syn_9/sky130_fd_sc_hs__or2_1_1/X prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_59/a_376_368#
+ prbs_generator_syn_9/sky130_fd_sc_hs__nand2_1_19/B prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_5/a_696_458#
+ prbs_generator_syn_9/sky130_fd_sc_hs__nor2b_1_1/Y prbs_generator_syn_9/sky130_fd_sc_hs__nor2b_1_5/a_278_368#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_17/a_1178_124# prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_39/X
+ prbs_generator_syn_9/m3_13600_5433# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_63/a_437_503#
+ prbs_generator_syn_9/sky130_fd_sc_hs__nand2_2_5/B prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_23/a_735_102#
+ prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_53/A prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_61/a_735_102#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_57/a_1034_424# prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_63/B
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_37/a_1141_508# prbs_generator_syn_9/sky130_fd_sc_hs__nand2_1_47/B
+ prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_29/X prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_65/Y
+ prbs_generator_syn_9/m3_13600_4701# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_1/a_437_503#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_67/a_1178_124# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_9/a_735_102#
+ prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_13/a_132_392# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_15/a_1178_124#
+ prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_15/A prbs_generator_syn_9/sky130_fd_sc_hs__nand2_1_1/B
+ prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_43/B prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_35/a_651_503#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_8/D prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_29/A
+ prbs_generator_syn_9/sky130_fd_sc_hs__nand2_1_7/B prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_13/a_735_102#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_47/a_696_458# prbs_generator_syn_9/sky130_fd_sc_hs__nand2_1_31/B
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_51/a_735_102# prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_59/X
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_35/a_1141_508# prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_25/a_222_392#
+ prbs_generator_syn_9/sky130_fd_sc_hs__sdlclkp_2_1/a_288_48# prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_55/B
+ prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_17/B prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_43/A
+ prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_7/A prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_65/a_1178_124#
+ prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_59/Y prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_41/X
+ prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_21/a_230_79# prbs_generator_syn_9/sky130_fd_sc_hs__nand2_1_57/a_117_74#
+ prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_1/a_222_392# prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_19/B
+ prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_35/a_293_74# prbs_generator_syn_9/sky130_fd_sc_hs__nand2_1_23/a_117_74#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_73/a_206_368# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_25/a_651_503#
+ prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_1/a_138_385# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_37/a_696_458#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_67/a_544_485# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_43/a_27_74#
+ prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_9/X prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_55/a_1034_424#
+ prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_39/a_112_119# prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_15/a_222_392#
+ prbs_generator_syn_9/sky130_fd_sc_hs__conb_1_1/HI prbs_generator_syn_9/sky130_fd_sc_hs__nand2_1_23/B
+ prbs_generator_syn_9/sky130_fd_sc_hs__nand2_1_53/B prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_9/a_1178_124#
+ prbs_generator_syn_9/sky130_fd_sc_hs__nor2b_1_4/A prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_47/a_1226_296#
+ prbs_generator_syn_9/m3_13600_11045# prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_17/X
+ prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_29/a_376_368# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_5/a_544_485#
+ prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_3/X prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_31/a_132_392#
+ prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_61/A prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_15/a_651_503#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_73/a_437_503# prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_25/a_230_79#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_27/a_696_458# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_65/a_696_458#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_33/a_735_102# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_71/a_735_102#
+ prbs_generator_syn_9/m3_13600_7263# prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_43/a_222_392#
+ prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_50/Y prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_8/a_1178_124#
+ prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_53/B prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_19/a_376_368#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_63/a_1178_124# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_4/a_696_458#
+ prbs_generator_syn_9/sky130_fd_sc_hs__nor2b_1_4/a_278_368# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_13/a_1178_124#
+ prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_61/a_132_392# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_53/a_206_368#
+ prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_21/a_52_123# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_45/a_651_503#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_17/a_696_458# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_47/a_544_485#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_55/a_696_458# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_21/a_735_102#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_37/a_27_74# prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_61/B
+ prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_61/X prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_59/a_112_119#
+ prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_31/A prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_33/a_222_392#
+ prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_29/a_230_79# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_45/a_1226_296#
+ prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_9/a_132_392# prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_5/A
+ prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_57/Y prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_31/X
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_51/a_27_74# prbs_generator_syn_9/sky130_fd_sc_hs__nor2b_1_8/a_27_112#
+ prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_47/a_376_368# prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_53/a_293_74#
+ prbs_generator_syn_9/sky130_fd_sc_hs__nand2_1_43/a_117_74# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_8/a_735_102#
+ prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_21/a_293_74# prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_39/a_138_385#
+ prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_63/Y prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_51/a_132_392#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_43/a_206_368# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_53/a_437_503#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_37/a_544_485# prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_57/X
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_53/a_1034_424# prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_25/a_52_123#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_33/a_1141_508# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_63/Q
+ prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_23/a_222_392# prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_63/a_222_392#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_7/a_1178_124# prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_53/X
+ prbs_generator_syn_9/sky130_fd_sc_hs__nand2_2_5/Y prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_61/a_1178_124#
+ prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_1/a_230_79# prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_43/a_230_79#
+ prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_11/a_230_79# prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_41/a_132_392#
+ prbs_generator_syn_9/sky130_fd_sc_hs__nand2_1_13/a_117_74# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_43/a_437_503#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_27/a_544_485# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_63/a_651_503#
+ prbs_generator_syn_9/sky130_fd_sc_hs__nand2_1_7/a_117_74# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_35/a_696_458#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_65/a_544_485# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_51/a_1034_424#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_41/a_735_102# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_32/a_1141_508#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_49/a_1141_508# prbs_generator_syn_9/sky130_fd_sc_hs__nand2_1_55/B
+ prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_53/a_222_392# prbs_generator_syn_9/sky130_fd_sc_hs__sdlclkp_2_1/a_114_112#
+ prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_9/a_293_74# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_43/a_1226_296#
+ prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_29/a_52_123# prbs_generator_syn_9/sky130_fd_sc_hs__nand2_1_37/B
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_1/a_651_503# prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_27/a_376_368#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_4/a_544_485# prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_67/a_376_368#
+ prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_27/X prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_1/X
+ prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_59/a_138_385# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_29/a_1178_124#
+ prbs_generator_syn_9/m3_13600_2871# prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_5/a_230_79#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_23/a_206_368# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_61/a_206_368#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_17/a_544_485# prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_15/a_230_79#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_25/a_696_458# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_55/a_544_485#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_32/a_735_102# prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_29/a_293_74#
+ prbs_generator_syn_9/sky130_fd_sc_hs__nand2_1_17/a_117_74# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_69/a_1034_424#
+ prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_29/a_112_119# prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_37/X
+ prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_31/B prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_19/a_1034_424#
+ prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_33/A prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_9/a_206_368#
+ prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_57/a_376_368# prbs_generator_syn_9/sky130_fd_sc_hs__sdlclkp_2_1/a_706_317#
+ prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_11/B prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_1/a_52_123#
+ prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_39/B prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_21/a_132_392#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_13/a_206_368# prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_43/a_52_123#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_51/a_206_368# prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_47/X
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_23/a_437_503# prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_11/a_52_123#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_61/a_437_503# prbs_generator_syn_9/sky130_fd_sc_hs__nor2b_1_7/Y
+ prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_51/A prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_15/a_696_458#
+ prbs_generator_syn_9/sky130_fd_sc_hs__nor2b_1_5/Y prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_9/a_230_79#
+ prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_25/X prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_19/a_112_119#
+ prbs_generator_syn_9/sky130_fd_sc_hs__nand2_1_45/B prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_5/a_1178_124#
+ prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_19/a_230_79# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_41/a_1226_296#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_59/a_1226_296# prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_63/a_230_79#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_51/Q prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_7/a_132_392#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_9/a_437_503# prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_46/a_376_368#
+ prbs_generator_syn_9/sky130_fd_sc_hs__nand2_1_33/a_117_74# prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_11/a_293_74#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_27/a_1178_124# prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_11/a_132_392#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_13/a_437_503# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_51/a_437_503#
+ prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_5/a_52_123# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_35/a_544_485#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_73/a_651_503# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_45/a_696_458#
+ prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_15/a_52_123# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_47/a_1141_508#
+ prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_47/a_112_119# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_4/a_1178_124#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_17/a_1034_424# prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_23/B
+ prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_37/a_376_368# prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_15/B
+ prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_7/Y prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_29/a_138_385#
+ prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_33/a_230_79# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_25/a_1178_124#
+ prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_47/a_293_74# prbs_generator_syn_9/sky130_fd_sc_hs__nand2_1_37/a_117_74#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_33/a_206_368# prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_15/a_293_74#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_71/a_206_368# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_25/a_544_485#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_67/a_1034_424# prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_13/a_222_392#
+ prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_9/a_52_123# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_15/a_1034_424#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_57/a_1226_296# prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_19/a_52_123#
+ prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_23/X prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_63/a_52_123#
+ prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_19/a_138_385# prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_9/a_376_368#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_21/a_206_368# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_33/a_437_503#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_71/a_437_503# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_53/a_651_503#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_15/a_544_485# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_63/a_696_458#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_65/a_1034_424# prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_19/a_293_74#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_45/a_1141_508# prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_27/a_112_119#
+ prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_67/a_112_119# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_1/a_1178_124#
+ prbs_generator_syn_9/sky130_fd_sc_hs__conb_1_1/a_21_290# prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_63/a_293_74#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_8/a_206_368# prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_17/a_376_368#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_63/a_27_74# prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_21/A
+ prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_55/a_376_368# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_1/a_696_458#
+ prbs_generator_syn_9/sky130_fd_sc_hs__nor2b_1_1/a_278_368# prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_47/a_138_385#
+ prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_33/a_52_123# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_9/a_1034_424#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_21/a_437_503# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_1/a_27_74#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_43/a_651_503# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_1/Q
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_45/a_544_485# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_69/a_735_102#
+ prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_57/a_112_119# prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_31/a_222_392#
+ prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_13/A prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_55/a_1226_296#
+ prbs_generator_syn_9/sky130_fd_sc_hs__nand2_2_5/a_27_74# prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_53/a_230_79#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_8/a_437_503# prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_67/a_293_74#
+ prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_33/a_293_74# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_7/a_735_102#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_23/a_1178_124# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_41/a_206_368#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_8/a_1034_424# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_63/a_1034_424#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_59/a_735_102# prbs_generator_syn_9/sky130_fd_sc_hs__nand2_1_5/B
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_43/a_1141_508# prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_46/a_112_119#
+ prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_61/a_222_392# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_13/a_1034_424#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_73/a_1178_124# prbs_generator_syn_9/sky130_fd_sc_hs__nand2_1_27/B
+ prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_13/B prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_57/a_27_74#
+ prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_57/a_230_79# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_21/a_1178_124#
+ prbs_generator_syn_9/sky130_fd_sc_hs__nor2b_1_1/a_27_112# prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_27/a_138_385#
+ prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_23/a_230_79# prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_67/a_138_385#
+ prbs_generator_syn_9/sky130_fd_sc_hs__nand2_1_41/B prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_9/a_222_392#
+ prbs_generator_syn_9/sky130_fd_sc_hs__nand2_1_27/a_117_74# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_32/a_206_368#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_23/a_651_503# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_41/a_437_503#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_73/a_27_74# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_61/a_651_503#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_63/a_544_485# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_49/a_735_102#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_73/a_696_458# prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_37/a_112_119#
+ prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_51/a_222_392# prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_43/X
+ prbs_generator_syn_9/sky130_fd_sc_hs__nand2_2_1/B prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_9/a_651_503#
+ prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_53/a_52_123# prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_49/X
+ prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_25/a_376_368# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_1/a_544_485#
+ prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_65/a_376_368# prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_57/a_138_385#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_27/a_27_74# prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_39/a_132_392#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_7/a_1034_424# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_13/a_651_503#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_32/a_437_503# prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_27/a_230_79#
+ prbs_generator_syn_9/m3_13600_12265# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_51/a_651_503#
+ prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_59/B prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_47/A
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_61/a_1034_424# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_41/a_1141_508#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_59/a_1141_508# prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_41/a_222_392#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_53/a_1226_296# prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_3/A
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_71/a_1178_124# prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_9/a_112_119#
+ prbs_generator_syn_9/sky130_fd_sc_hs__nand2_1_3/a_117_74# prbs_generator_syn_9/m3_13600_8483#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_39/a_1178_124# prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_57/a_52_123#
+ prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_46/a_138_385# prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_23/a_52_123#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_67/a_27_74# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_53/a_696_458#
+ prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_17/a_112_119# prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_11/A
+ prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_55/a_112_119# prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_1/A
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_51/a_1226_296# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_29/a_1034_424#
+ prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_59/A prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_23/A
+ prbs_generator_syn_9/sky130_fd_sc_hs__nand2_1_39/B prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_5/a_27_74#
+ prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_57/a_293_74# prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_37/a_138_385#
+ prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_59/a_132_392# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_33/a_651_503#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_71/a_651_503# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_43/a_696_458#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_73/a_544_485# prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_27/a_52_123#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_57/a_1141_508# prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_21/a_222_392#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_35/a_27_74# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_69/a_1226_296#
+ prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_37/B prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_19/a_1226_296#
+ prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_35/a_376_368# prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_47/a_230_79#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_37/a_1178_124# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_5/a_1034_424#
+ prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_49/a_132_392# prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_7/a_222_392#
+ prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_27/a_293_74# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_21/a_651_503#
+ prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_9/a_138_385# prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_11/a_222_392#
+ prbs_generator_syn_9/m3_13600_14095# prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_50/A
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_27/a_1034_424# prbs_generator_syn_9/sky130_fd_sc_hs__nand2_1_13/B
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_8/a_651_503# prbs_generator_syn_9/m3_13600_9703#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_35/a_1178_124# prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_17/a_138_385#
+ prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_55/a_138_385# prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_7/a_230_79#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_4/a_1034_424# prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_7/a_376_368#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_69/a_206_368# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_23/a_696_458#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_53/a_544_485# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_39/a_735_102#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_61/a_696_458# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_55/a_1141_508#
+ prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_25/a_112_119# prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_65/a_112_119#
+ prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_43/a_293_74# prbs_generator_syn_9/sky130_fd_sc_hs__nand2_1_57/B
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_25/a_1034_424# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_7/a_206_368#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_17/a_1226_296# prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_15/a_376_368#
+ prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_53/a_376_368# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_9/a_696_458#
+ prbs_generator_syn_9/m3_13600_431# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_45/a_27_74#
+ prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_47/a_52_123# prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_29/a_132_392#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_59/a_206_368# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_69/a_437_503#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_41/a_651_503# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_43/a_544_485#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_13/a_696_458# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_29/a_735_102#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_51/a_696_458# prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_61/Y
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_67/a_1226_296# prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_5/a_132_392#
+ prbs_generator_syn_9/sky130_fd_sc_hs__and2b_2_1/a_198_48# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_7/a_437_503#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_15/a_1226_296# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_69/a_27_74#
+ prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_46/a_293_74# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_1/a_1034_424#
+ prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_19/a_132_392# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_49/a_206_368#
+ prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_7/a_52_123# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_59/a_437_503#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_32/a_651_503# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_7/a_27_74#
+ prbs_generator_syn_9/sky130_fd_sc_hs__nand2_2_1/a_27_74# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_19/a_735_102#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_57/a_735_102# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_65/a_1226_296#
+ prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_37/A prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_33/a_376_368#
+ prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_37/a_230_79# prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_25/a_138_385#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_39/a_27_74# prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_65/a_138_385#
+ prbs_generator_syn_9/sky130_fd_sc_hs__nor2b_1_9/a_278_368# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_49/a_437_503#
+ prbs_generator_syn_9/sky130_fd_sc_hs__and2b_2_1/a_505_74# prbs_generator_syn_9/sky130_fd_sc_hs__nand2_1_51/a_117_74#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_23/a_544_485# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_33/a_696_458#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_61/a_544_485# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_9/a_1226_296#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_53/a_1141_508# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_71/a_696_458#
+ prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_35/a_112_119# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_23/a_1034_424#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_9/a_544_485# prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_63/a_376_368#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_33/a_1178_124# prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_5/a_376_368#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_13/a_544_485# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_73/a_1034_424#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_21/a_696_458# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_51/a_544_485#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_8/a_1226_296# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_51/a_1141_508#
+ prbs_generator_syn_9/sky130_fd_sc_hs__nand2_1_55/a_117_74# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_21/a_1034_424#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_63/a_1226_296# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_23/a_27_74#
+ prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_7/a_112_119# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_13/a_1226_296#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_8/a_696_458# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_32/a_1178_124#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_49/a_1178_124# prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_37/a_52_123#
+ prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_27/a_132_392# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_71/Q
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_67/a_735_102# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_69/a_1141_508#
+ prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_15/a_112_119# prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_53/a_112_119#
+ prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_39/a_222_392# prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_55/a_230_79#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_19/a_1141_508# prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_37/a_293_74#
+ prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_43/a_376_368# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_5/a_735_102#
+ prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_35/a_138_385# prbs_generator_syn_9/sky130_fd_sc_hs__sdlclkp_2_1/a_114_424#
+ prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_57/a_132_392# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_71/a_1034_424#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_7/a_1226_296# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_33/a_544_485#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_41/a_696_458# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_71/a_544_485#
+ prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_21/B prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_61/a_1226_296#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_39/a_1034_424# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_17/a_27_74#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_9/a_27_74# prbs_generator_syn_9/sky130_fd_sc_hs__nor2b_1_5/a_27_112#
+ prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_47/a_132_392# prbs_generator_syn_9/sky130_fd_sc_hs__nor2b_1_8/a_278_368#
+ prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_9/B prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_39/a_206_368#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_33/a_27_74# prbs_generator_syn_9/sky130_fd_sc_hs__nand2_1_41/a_117_74#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_69/a_651_503# prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_51/a_293_74#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_21/a_544_485# prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_7/a_138_385#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_32/a_696_458# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_47/a_735_102#
+ prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_33/a_112_119# prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_59/a_222_392#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_17/a_1141_508# prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_55/a_52_123#
+ prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_3/a_293_74# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_7/a_651_503#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_29/a_1226_296# prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_23/a_376_368#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_8/a_544_485# prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_47/B
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_47/a_1178_124# prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_15/a_138_385#
+ prbs_generator_syn_9/sky130_fd_sc_hs__sdlclkp_2_1/a_1195_374# prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_53/a_138_385#
+ prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_37/a_132_392# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_29/a_206_368#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_39/a_437_503# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_59/a_651_503#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_37/a_735_102# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_67/a_1141_508#
+ prbs_generator_syn_9/sky130_fd_sc_hs__and2b_2_1/a_27_74# prbs_generator_syn_9/sky130_fd_sc_hs__conb_1_1/a_165_290#
+ prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_55/a_293_74# prbs_generator_syn_9/sky130_fd_sc_hs__nand2_1_45/a_117_74#
+ prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_63/a_112_119# prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_49/a_222_392#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_37/a_1034_424# prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_23/a_293_74#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_15/a_1141_508# prbs_generator_syn_9/sky130_fd_sc_hs__nand2_1_5/a_117_74#
+ prbs_generator_syn_9/m3_13600_13485# prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_5/a_112_119#
+ prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_13/a_376_368# prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_51/a_376_368#
+ prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_7/a_293_74# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_19/a_206_368#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_57/a_206_368# prbs_generator_syn_9/sky130_fd_sc_hs__sdlclkp_2_1/a_318_74#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_29/a_437_503# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_49/a_651_503#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_25/a_27_74# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_5/a_1226_296#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_41/a_544_485# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_27/a_735_102#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_65/a_1141_508# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_65/a_735_102#
+ prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_3/a_230_79# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_35/a_1034_424#
+ prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_13/a_230_79# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_41/a_27_74#
+ prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_3/a_132_392# prbs_generator_syn_9/sky130_fd_sc_hs__nand2_1_49/a_117_74#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_27/a_1226_296# prbs_generator_syn_9/sky130_fd_sc_hs__nand2_1_15/a_117_74#
+ prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_41/a_376_368# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_45/a_1178_124#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_4/a_735_102# prbs_generator_syn_9/sky130_fd_sc_hs__nand2_1_9/a_117_74#
+ prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_33/a_138_385# prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_17/a_132_392#
+ prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_55/a_132_392# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_9/a_1141_508#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_19/a_437_503# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_57/a_437_503#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_4/a_1226_296# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_32/a_544_485#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_17/a_735_102# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_55/a_735_102#
+ prbs_generator_syn_9/m3_13600_2261# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_65/a_27_74#
+ prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_29/a_222_392# prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_43/a_112_119#
+ prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_19/X prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_25/a_1226_296#
+ prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_31/a_376_368# prbs_generator_syn_9/sky130_fd_sc_hs__or2_1_1/a_63_368#
+ prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_17/a_230_79# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_4/a_27_74#
+ prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_61/a_230_79# prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_63/a_138_385#
+ prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_5/a_222_392# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_8/a_1141_508#
+ prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_41/a_293_74# prbs_generator_syn_9/sky130_fd_sc_hs__nand2_1_31/a_117_74#
+ prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_5/a_138_385# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_63/a_1141_508#
+ prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_19/a_222_392# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_13/a_1141_508#
+ prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_3/a_52_123# prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_13/a_52_123#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_43/a_1178_124# prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_61/a_376_368#
+ prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_35/a_132_392# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_67/a_206_368#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_1/a_1226_296# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_69/a_696_458#
+ prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_31/a_230_79# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_35/a_735_102#
+ prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_23/a_112_119# prbs_generator_syn_9/sky130_fd_sc_hs__nand2_1_35/a_117_74#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_59/a_27_74# prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_13/a_293_74#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_5/a_206_368# prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_50/a_376_368#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_7/a_696_458# prbs_generator_syn_9/sky130_fd_sc_hs__nor2b_1_7/a_278_368#
+ prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_17/a_52_123# prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_43/a_138_385#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_7/a_1141_508# prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_61/a_52_123#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_67/a_437_503# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_61/a_1141_508#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_25/a_735_102# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_59/a_696_458#
+ prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_13/a_112_119# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_33/a_1034_424#
+ prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_51/a_112_119# prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_35/a_230_79#
+ prbs_generator_syn_9/m3_13600_4091# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_23/a_1226_296#
+ prbs_generator_syn_9/sky130_fd_sc_hs__nand2_1_39/a_117_74# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_29/a_27_74#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_5/a_437_503# prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_17/a_293_74#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_41/a_1178_124# prbs_generator_syn_9/sky130_fd_sc_hs__or2_1_1/a_152_368#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_59/a_1178_124# prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_61/a_293_74#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_47/a_206_368# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_39/a_651_503#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_49/a_696_458# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_15/a_735_102#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_32/a_1034_424# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_73/a_1226_296#
+ prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_27/a_222_392# prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_41/a_112_119#
+ prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_31/a_52_123# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_49/a_1034_424#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_29/a_1141_508# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_21/a_1226_296#
+ prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_39/a_230_79# prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_23/a_138_385#
+ prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_51/a_230_79# prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_45/a_132_392#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_37/a_206_368# prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_65/a_293_74#
+ prbs_generator_syn_9/sky130_fd_sc_hs__nand2_1_53/a_117_74# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_47/a_437_503#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_29/a_651_503# prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_31/a_293_74#
+ prbs_generator_syn_9/sky130_fd_sc_hs__nand2_1_21/a_117_74# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_69/a_544_485#
+ prbs_generator_syn_9/sky130_fd_sc_hs__clkbuf_16_1/a_114_74# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_45/a_735_102#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_13/a_27_74# prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_31/a_112_119#
+ prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_57/a_222_392# prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_35/a_52_123#
+ prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_21/a_376_368# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_7/a_544_485#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_57/a_1178_124# prbs_generator_syn_9/m3_13600_6043#
+ prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_13/a_138_385# prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_51/a_138_385#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_5/a_1141_508# prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_3/a_376_368#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_27/a_206_368# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_65/a_206_368#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_37/a_437_503# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_19/a_651_503#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_57/a_651_503# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_59/a_544_485#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_71/a_1226_296# prbs_generator_syn_9/sky130_fd_sc_hs__nand2_1_25/a_117_74#
+ prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_61/a_112_119# prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_47/a_222_392#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_27/a_1141_508# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_53/a_27_74#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_4/a_206_368# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_39/a_1226_296#
+ prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_11/a_376_368# prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_39/a_52_123#
+ prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_41/a_138_385# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_4/a_1141_508#
+ prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_25/a_132_392# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_17/a_206_368#
+ prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_41/A prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_55/a_206_368#
+ prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_51/a_52_123# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_27/a_437_503#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_65/a_437_503# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_49/a_544_485#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_63/a_735_102# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_47/a_1034_424#
+ prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_50/a_112_119# prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_37/a_222_392#
+ prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_59/a_230_79# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_25/a_1141_508#
+ prbs_generator_syn_9/sky130_fd_sc_hs__nor2b_1_4/a_27_112# prbs_generator_syn_9/sky130_fd_sc_hs__sdlclkp_2_1/a_685_81#
+ prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_1/a_132_392# prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_39/a_293_74#
+ prbs_generator_syn_9/sky130_fd_sc_hs__nand2_1_29/a_117_74# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_4/a_437_503#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_55/a_1178_124# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_21/a_27_74#
+ prbs_generator_syn_9/m3_13600_12875# prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_50/a_293_74#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_1/a_735_102# prbs_generator_syn_9/sky130_fd_sc_hs__xnor2_1_31/a_138_385#
+ prbs_generator_syn_9/sky130_fd_sc_hs__a22o_1_15/a_132_392# prbs_generator_syn_9/sky130_fd_sc_hs__nand2_1_1/a_117_74#
+ prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_17/a_437_503# prbs_generator_syn_9/sky130_fd_sc_hs__dfxtp_4_55/a_437_503#
+ prbs_generator_syn
Xsky130_fd_sc_hs__clkbuf_4_101 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__clkbuf_4_109/X
+ fine_freq_track_1/fftl_en sky130_fd_sc_hs__clkbuf_4_101/a_83_270# sky130_fd_sc_hs__clkbuf_4
Xsky130_fd_sc_hs__clkbuf_4_112 DVSS: DVDD: DVDD: DVSS: CTL_BUF_P[4] sky130_fd_sc_hs__clkbuf_4_113/X
+ sky130_fd_sc_hs__clkbuf_4_113/a_83_270# sky130_fd_sc_hs__clkbuf_4
Xsky130_fd_sc_hs__clkbuf_4_123 DVSS: DVDD: DVDD: DVSS: CTL_BUF_N[5] sky130_fd_sc_hs__clkbuf_4_123/X
+ sky130_fd_sc_hs__clkbuf_4_123/a_83_270# sky130_fd_sc_hs__clkbuf_4
Xsky130_fd_sc_hs__clkbuf_4_134 DVSS: DVDD: DVDD: DVSS: rst_prbs sky130_fd_sc_hs__clkbuf_8_93/A
+ sky130_fd_sc_hs__clkbuf_4_135/a_83_270# sky130_fd_sc_hs__clkbuf_4
Xsky130_fd_sc_hs__o21ai_2_3 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__inv_4_13/Y sky130_fd_sc_hs__o21ai_2_3/A2
+ sky130_fd_sc_hs__nand2_2_9/B sky130_fd_sc_hs__buf_2_41/A sky130_fd_sc_hs__o21ai_2_3/a_116_368#
+ sky130_fd_sc_hs__o21ai_2_3/a_27_74# sky130_fd_sc_hs__o21ai_2
Xsky130_fd_sc_hs__clkbuf_4_30 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__buf_2_11/X
+ sky130_fd_sc_hs__clkbuf_8_27/A sky130_fd_sc_hs__clkbuf_4_31/a_83_270# sky130_fd_sc_hs__clkbuf_4
Xsky130_fd_sc_hs__clkbuf_4_41 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__clkbuf_4_47/X
+ sky130_fd_sc_hs__clkbuf_4_41/X sky130_fd_sc_hs__clkbuf_4_41/a_83_270# sky130_fd_sc_hs__clkbuf_4
Xsky130_fd_sc_hs__clkbuf_4_52 DVSS: DVDD: DVDD: DVSS: fine_con_step_size[3] sky130_fd_sc_hs__clkbuf_4_53/X
+ sky130_fd_sc_hs__clkbuf_4_53/a_83_270# sky130_fd_sc_hs__clkbuf_4
Xsky130_fd_sc_hs__clkbuf_4_63 DVSS: DVDD: DVDD: DVSS: fine_control_avg_window_select[2]
+ sky130_fd_sc_hs__clkbuf_4_63/X sky130_fd_sc_hs__clkbuf_4_63/a_83_270# sky130_fd_sc_hs__clkbuf_4
Xsky130_fd_sc_hs__clkbuf_4_74 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__or2b_4_5/A
+ sky130_fd_sc_hs__o21ai_2_9/A2 sky130_fd_sc_hs__clkbuf_4_75/a_83_270# sky130_fd_sc_hs__clkbuf_4
Xsky130_fd_sc_hs__clkbuf_4_85 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__buf_2_131/X
+ sky130_fd_sc_hs__inv_4_23/A sky130_fd_sc_hs__clkbuf_4_85/a_83_270# sky130_fd_sc_hs__clkbuf_4
Xsky130_fd_sc_hs__clkbuf_4_96 DVSS: DVDD: DVDD: DVSS: div_ratio_half[1] sky130_fd_sc_hs__clkbuf_4_97/X
+ sky130_fd_sc_hs__clkbuf_4_97/a_83_270# sky130_fd_sc_hs__clkbuf_4
Xsky130_fd_sc_hs__clkinv_8_11 DVSS: DVDD: DVDD: DVSS: prbs_generator_syn_5/out hr_16t4_mux_top_3/din[7]
+ sky130_fd_sc_hs__clkinv_8
Xsky130_fd_sc_hs__einvn_4_0 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__clkinv_8_15/Y
+ osc_core_1/p3 qr_4t1_mux_top_3/clk_IB sky130_fd_sc_hs__einvn_4_1/a_114_74# sky130_fd_sc_hs__einvn_4_1/a_241_368#
+ sky130_fd_sc_hs__einvn_4_1/a_281_74# sky130_fd_sc_hs__einvn_4
Xsky130_fd_sc_hs__conb_1_120 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__conb_1_121/LO
+ sky130_fd_sc_hs__conb_1_121/HI sky130_fd_sc_hs__conb_1_121/a_165_290# sky130_fd_sc_hs__conb_1_121/a_21_290#
+ sky130_fd_sc_hs__conb_1
Xsky130_fd_sc_hs__conb_1_131 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__conb_1_131/LO
+ sky130_fd_sc_hs__conb_1_131/HI sky130_fd_sc_hs__conb_1_131/a_165_290# sky130_fd_sc_hs__conb_1_131/a_21_290#
+ sky130_fd_sc_hs__conb_1
Xsky130_fd_sc_hs__conb_1_142 DVSS: DVDD: DVDD: DVSS: prbs_generator_syn_15/eqn[31]
+ prbs_generator_syn_15/cke sky130_fd_sc_hs__conb_1_143/a_165_290# sky130_fd_sc_hs__conb_1_143/a_21_290#
+ sky130_fd_sc_hs__conb_1
Xsky130_fd_sc_hs__conb_1_153 DVSS: DVDD: DVDD: DVSS: prbs_generator_syn_17/eqn[9]
+ sky130_fd_sc_hs__conb_1_153/HI sky130_fd_sc_hs__conb_1_153/a_165_290# sky130_fd_sc_hs__conb_1_153/a_21_290#
+ sky130_fd_sc_hs__conb_1
Xsky130_fd_sc_hs__conb_1_164 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__conb_1_165/LO
+ sky130_fd_sc_hs__conb_1_165/HI sky130_fd_sc_hs__conb_1_165/a_165_290# sky130_fd_sc_hs__conb_1_165/a_21_290#
+ sky130_fd_sc_hs__conb_1
Xsky130_fd_sc_hs__conb_1_175 DVSS: DVDD: DVDD: DVSS: prbs_generator_syn_23/eqn[9]
+ sky130_fd_sc_hs__conb_1_175/HI sky130_fd_sc_hs__conb_1_175/a_165_290# sky130_fd_sc_hs__conb_1_175/a_21_290#
+ sky130_fd_sc_hs__conb_1
Xsky130_fd_sc_hs__conb_1_186 DVSS: DVDD: DVDD: DVSS: prbs_generator_syn_23/eqn[0]
+ sky130_fd_sc_hs__conb_1_187/HI sky130_fd_sc_hs__conb_1_187/a_165_290# sky130_fd_sc_hs__conb_1_187/a_21_290#
+ sky130_fd_sc_hs__conb_1
Xsky130_fd_sc_hs__conb_1_197 DVSS: DVDD: DVDD: DVSS: prbs_generator_syn_19/eqn[22]
+ prbs_generator_syn_19/eqn[20] sky130_fd_sc_hs__conb_1_197/a_165_290# sky130_fd_sc_hs__conb_1_197/a_21_290#
+ sky130_fd_sc_hs__conb_1
Xsky130_fd_sc_hs__einvp_2_120 DVSS: DVDD: DVDD: DVSS: dout_n sky130_fd_sc_hs__buf_8_1/X
+ sky130_fd_sc_hs__buf_2_119/X sky130_fd_sc_hs__einvp_2_121/a_263_323# sky130_fd_sc_hs__einvp_2_121/a_36_74#
+ sky130_fd_sc_hs__einvp_2_121/a_27_368# sky130_fd_sc_hs__einvp_2
Xsky130_fd_sc_hs__einvp_2_131 DVSS: DVDD: DVDD: DVSS: dout_n sky130_fd_sc_hs__buf_8_1/X
+ sky130_fd_sc_hs__dlrtp_1_127/Q sky130_fd_sc_hs__einvp_2_131/a_263_323# sky130_fd_sc_hs__einvp_2_131/a_36_74#
+ sky130_fd_sc_hs__einvp_2_131/a_27_368# sky130_fd_sc_hs__einvp_2
Xsky130_fd_sc_hs__einvp_2_142 DVSS: DVDD: DVDD: DVSS: dout_p sky130_fd_sc_hs__einvp_2_99/A
+ sky130_fd_sc_hs__dlrtp_1_139/Q sky130_fd_sc_hs__einvp_2_143/a_263_323# sky130_fd_sc_hs__einvp_2_143/a_36_74#
+ sky130_fd_sc_hs__einvp_2_143/a_27_368# sky130_fd_sc_hs__einvp_2
Xsky130_fd_sc_hs__einvp_2_153 DVSS: DVDD: DVDD: DVSS: dout_p sky130_fd_sc_hs__einvp_2_99/A
+ sky130_fd_sc_hs__dlrtp_1_157/Q sky130_fd_sc_hs__einvp_2_153/a_263_323# sky130_fd_sc_hs__einvp_2_153/a_36_74#
+ sky130_fd_sc_hs__einvp_2_153/a_27_368# sky130_fd_sc_hs__einvp_2
Xsky130_fd_sc_hs__clkbuf_16_14 DVSS: DVDD: DVDD: DVSS: prbs_generator_syn_9/clk sky130_fd_sc_hs__clkbuf_16_75/X
+ sky130_fd_sc_hs__clkbuf_16_15/a_114_74# sky130_fd_sc_hs__clkbuf_16
Xsky130_fd_sc_hs__clkbuf_16_25 DVSS: DVDD: DVDD: DVSS: osc_core_1/pi3_l[3] sky130_fd_sc_hs__clkbuf_8_11/X
+ sky130_fd_sc_hs__clkbuf_16_25/a_114_74# sky130_fd_sc_hs__clkbuf_16
Xsky130_fd_sc_hs__clkbuf_16_36 DVSS: DVDD: DVDD: DVSS: osc_core_1/pi2_l[2] sky130_fd_sc_hs__clkbuf_8_3/X
+ sky130_fd_sc_hs__clkbuf_16_37/a_114_74# sky130_fd_sc_hs__clkbuf_16
Xsky130_fd_sc_hs__clkbuf_16_47 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__buf_8_1/A
+ sky130_fd_sc_hs__nand2_2_1/Y sky130_fd_sc_hs__clkbuf_16_47/a_114_74# sky130_fd_sc_hs__clkbuf_16
Xsky130_fd_sc_hs__clkbuf_16_58 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__o21ai_4_1/A1
+ sky130_fd_sc_hs__clkbuf_16_93/X sky130_fd_sc_hs__clkbuf_16_59/a_114_74# sky130_fd_sc_hs__clkbuf_16
Xsky130_fd_sc_hs__clkbuf_16_69 DVSS: DVDD: DVDD: DVSS: qr_4t1_mux_top_1/rst qr_4t1_mux_top_3/rst
+ sky130_fd_sc_hs__clkbuf_16_69/a_114_74# sky130_fd_sc_hs__clkbuf_16
Xsky130_fd_sc_hs__clkbuf_16_102 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__clkbuf_8_67/A
+ sky130_fd_sc_hs__clkbuf_4_127/X sky130_fd_sc_hs__clkbuf_16_103/a_114_74# sky130_fd_sc_hs__clkbuf_16
Xsky130_fd_sc_hs__clkbuf_16_113 DVSS: DVDD: DVDD: DVSS: prbs_generator_syn_31/inj_err
+ prbs_generator_syn_27/inj_err sky130_fd_sc_hs__clkbuf_16_113/a_114_74# sky130_fd_sc_hs__clkbuf_16
Xsky130_fd_sc_hs__clkbuf_16_124 DVSS: DVDD: DVDD: DVSS: osc_core_1/pi5_l[2] sky130_fd_sc_hs__clkbuf_4_131/X
+ sky130_fd_sc_hs__clkbuf_16_125/a_114_74# sky130_fd_sc_hs__clkbuf_16
Xsky130_fd_sc_hs__clkbuf_4_102 DVSS: DVDD: DVDD: DVSS: con_perb[1] osc_core_1/con_perb_5[1]
+ sky130_fd_sc_hs__clkbuf_4_103/a_83_270# sky130_fd_sc_hs__clkbuf_4
Xsky130_fd_sc_hs__clkbuf_4_113 DVSS: DVDD: DVDD: DVSS: CTL_BUF_P[4] sky130_fd_sc_hs__clkbuf_4_113/X
+ sky130_fd_sc_hs__clkbuf_4_113/a_83_270# sky130_fd_sc_hs__clkbuf_4
Xsky130_fd_sc_hs__clkbuf_4_124 DVSS: DVDD: DVDD: DVSS: pi5_con[1] sky130_fd_sc_hs__clkbuf_4_125/X
+ sky130_fd_sc_hs__clkbuf_4_125/a_83_270# sky130_fd_sc_hs__clkbuf_4
Xsky130_fd_sc_hs__clkbuf_4_135 DVSS: DVDD: DVDD: DVSS: rst_prbs sky130_fd_sc_hs__clkbuf_8_93/A
+ sky130_fd_sc_hs__clkbuf_4_135/a_83_270# sky130_fd_sc_hs__clkbuf_4
Xsky130_fd_sc_hs__o21ai_2_4 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__inv_4_13/Y sky130_fd_sc_hs__o21ai_2_9/A2
+ sky130_fd_sc_hs__nand2_2_9/B sky130_fd_sc_hs__o21ai_2_5/Y sky130_fd_sc_hs__o21ai_2_5/a_116_368#
+ sky130_fd_sc_hs__o21ai_2_5/a_27_74# sky130_fd_sc_hs__o21ai_2
Xsky130_fd_sc_hs__clkbuf_4_20 DVSS: DVDD: DVDD: DVSS: pi1_con[2] sky130_fd_sc_hs__clkbuf_4_21/X
+ sky130_fd_sc_hs__clkbuf_4_21/a_83_270# sky130_fd_sc_hs__clkbuf_4
Xsky130_fd_sc_hs__clkbuf_4_31 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__buf_2_11/X
+ sky130_fd_sc_hs__clkbuf_8_27/A sky130_fd_sc_hs__clkbuf_4_31/a_83_270# sky130_fd_sc_hs__clkbuf_4
Xsky130_fd_sc_hs__clkbuf_4_42 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__einvn_8_1/Z
+ qr_4t1_mux_top_1/clk_Q sky130_fd_sc_hs__clkbuf_4_43/a_83_270# sky130_fd_sc_hs__clkbuf_4
Xsky130_fd_sc_hs__clkbuf_4_53 DVSS: DVDD: DVDD: DVSS: fine_con_step_size[3] sky130_fd_sc_hs__clkbuf_4_53/X
+ sky130_fd_sc_hs__clkbuf_4_53/a_83_270# sky130_fd_sc_hs__clkbuf_4
Xsky130_fd_sc_hs__clkbuf_4_64 DVSS: DVDD: DVDD: DVSS: fine_control_avg_window_select[4]
+ sky130_fd_sc_hs__clkbuf_4_65/X sky130_fd_sc_hs__clkbuf_4_65/a_83_270# sky130_fd_sc_hs__clkbuf_4
Xsky130_fd_sc_hs__clkbuf_4_75 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__or2b_4_5/A
+ sky130_fd_sc_hs__o21ai_2_9/A2 sky130_fd_sc_hs__clkbuf_4_75/a_83_270# sky130_fd_sc_hs__clkbuf_4
Xsky130_fd_sc_hs__clkbuf_4_86 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__or2b_2_3/A
+ sky130_fd_sc_hs__o21ai_2_51/A1 sky130_fd_sc_hs__clkbuf_4_87/a_83_270# sky130_fd_sc_hs__clkbuf_4
Xsky130_fd_sc_hs__clkbuf_4_97 DVSS: DVDD: DVDD: DVSS: div_ratio_half[1] sky130_fd_sc_hs__clkbuf_4_97/X
+ sky130_fd_sc_hs__clkbuf_4_97/a_83_270# sky130_fd_sc_hs__clkbuf_4
Xsky130_fd_sc_hs__clkinv_8_12 DVSS: DVDD: DVDD: DVSS: prbs_generator_syn_9/out hr_16t4_mux_top_3/din[3]
+ sky130_fd_sc_hs__clkinv_8
Xsky130_fd_sc_hs__einvn_4_1 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__clkinv_8_15/Y
+ osc_core_1/p3 qr_4t1_mux_top_3/clk_IB sky130_fd_sc_hs__einvn_4_1/a_114_74# sky130_fd_sc_hs__einvn_4_1/a_241_368#
+ sky130_fd_sc_hs__einvn_4_1/a_281_74# sky130_fd_sc_hs__einvn_4
Xsky130_fd_sc_hs__conb_1_110 DVSS: DVDD: DVDD: DVSS: prbs_generator_syn_15/eqn[13]
+ sky130_fd_sc_hs__conb_1_111/HI sky130_fd_sc_hs__conb_1_111/a_165_290# sky130_fd_sc_hs__conb_1_111/a_21_290#
+ sky130_fd_sc_hs__conb_1
Xsky130_fd_sc_hs__conb_1_121 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__conb_1_121/LO
+ sky130_fd_sc_hs__conb_1_121/HI sky130_fd_sc_hs__conb_1_121/a_165_290# sky130_fd_sc_hs__conb_1_121/a_21_290#
+ sky130_fd_sc_hs__conb_1
Xsky130_fd_sc_hs__conb_1_132 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__conb_1_133/LO
+ sky130_fd_sc_hs__conb_1_133/HI sky130_fd_sc_hs__conb_1_133/a_165_290# sky130_fd_sc_hs__conb_1_133/a_21_290#
+ sky130_fd_sc_hs__conb_1
Xsky130_fd_sc_hs__conb_1_143 DVSS: DVDD: DVDD: DVSS: prbs_generator_syn_15/eqn[31]
+ prbs_generator_syn_15/cke sky130_fd_sc_hs__conb_1_143/a_165_290# sky130_fd_sc_hs__conb_1_143/a_21_290#
+ sky130_fd_sc_hs__conb_1
Xsky130_fd_sc_hs__conb_1_154 DVSS: DVDD: DVDD: DVSS: prbs_generator_syn_17/eqn[22]
+ prbs_generator_syn_17/eqn[20] sky130_fd_sc_hs__conb_1_155/a_165_290# sky130_fd_sc_hs__conb_1_155/a_21_290#
+ sky130_fd_sc_hs__conb_1
Xsky130_fd_sc_hs__conb_1_165 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__conb_1_165/LO
+ sky130_fd_sc_hs__conb_1_165/HI sky130_fd_sc_hs__conb_1_165/a_165_290# sky130_fd_sc_hs__conb_1_165/a_21_290#
+ sky130_fd_sc_hs__conb_1
Xsky130_fd_sc_hs__conb_1_176 DVSS: DVDD: DVDD: DVSS: prbs_generator_syn_21/eqn[0]
+ sky130_fd_sc_hs__conb_1_177/HI sky130_fd_sc_hs__conb_1_177/a_165_290# sky130_fd_sc_hs__conb_1_177/a_21_290#
+ sky130_fd_sc_hs__conb_1
Xsky130_fd_sc_hs__conb_1_187 DVSS: DVDD: DVDD: DVSS: prbs_generator_syn_23/eqn[0]
+ sky130_fd_sc_hs__conb_1_187/HI sky130_fd_sc_hs__conb_1_187/a_165_290# sky130_fd_sc_hs__conb_1_187/a_21_290#
+ sky130_fd_sc_hs__conb_1
Xsky130_fd_sc_hs__conb_1_198 DVSS: DVDD: DVDD: DVSS: prbs_generator_syn_19/eqn[2]
+ prbs_generator_syn_19/eqn[1] sky130_fd_sc_hs__conb_1_199/a_165_290# sky130_fd_sc_hs__conb_1_199/a_21_290#
+ sky130_fd_sc_hs__conb_1
Xsky130_fd_sc_hs__einvp_2_110 DVSS: DVDD: DVDD: DVSS: dout_n sky130_fd_sc_hs__einvp_2_9/A
+ sky130_fd_sc_hs__dlrtp_1_97/Q sky130_fd_sc_hs__einvp_2_111/a_263_323# sky130_fd_sc_hs__einvp_2_111/a_36_74#
+ sky130_fd_sc_hs__einvp_2_111/a_27_368# sky130_fd_sc_hs__einvp_2
Xsky130_fd_sc_hs__einvp_2_121 DVSS: DVDD: DVDD: DVSS: dout_n sky130_fd_sc_hs__buf_8_1/X
+ sky130_fd_sc_hs__buf_2_119/X sky130_fd_sc_hs__einvp_2_121/a_263_323# sky130_fd_sc_hs__einvp_2_121/a_36_74#
+ sky130_fd_sc_hs__einvp_2_121/a_27_368# sky130_fd_sc_hs__einvp_2
Xsky130_fd_sc_hs__einvp_2_132 DVSS: DVDD: DVDD: DVSS: dout_p sky130_fd_sc_hs__einvp_2_99/A
+ sky130_fd_sc_hs__dlrtp_1_131/Q sky130_fd_sc_hs__einvp_2_133/a_263_323# sky130_fd_sc_hs__einvp_2_133/a_36_74#
+ sky130_fd_sc_hs__einvp_2_133/a_27_368# sky130_fd_sc_hs__einvp_2
Xsky130_fd_sc_hs__einvp_2_143 DVSS: DVDD: DVDD: DVSS: dout_p sky130_fd_sc_hs__einvp_2_99/A
+ sky130_fd_sc_hs__dlrtp_1_139/Q sky130_fd_sc_hs__einvp_2_143/a_263_323# sky130_fd_sc_hs__einvp_2_143/a_36_74#
+ sky130_fd_sc_hs__einvp_2_143/a_27_368# sky130_fd_sc_hs__einvp_2
Xsky130_fd_sc_hs__einvp_2_154 DVSS: DVDD: DVDD: DVSS: dout_p sky130_fd_sc_hs__einvp_2_99/A
+ sky130_fd_sc_hs__buf_2_161/X sky130_fd_sc_hs__einvp_2_155/a_263_323# sky130_fd_sc_hs__einvp_2_155/a_36_74#
+ sky130_fd_sc_hs__einvp_2_155/a_27_368# sky130_fd_sc_hs__einvp_2
Xsky130_fd_sc_hs__clkbuf_16_15 DVSS: DVDD: DVDD: DVSS: prbs_generator_syn_9/clk sky130_fd_sc_hs__clkbuf_16_75/X
+ sky130_fd_sc_hs__clkbuf_16_15/a_114_74# sky130_fd_sc_hs__clkbuf_16
Xsky130_fd_sc_hs__clkbuf_16_26 DVSS: DVDD: DVDD: DVSS: osc_core_1/pi3_l[2] sky130_fd_sc_hs__clkbuf_8_7/X
+ sky130_fd_sc_hs__clkbuf_16_27/a_114_74# sky130_fd_sc_hs__clkbuf_16
Xsky130_fd_sc_hs__clkbuf_16_37 DVSS: DVDD: DVDD: DVSS: osc_core_1/pi2_l[2] sky130_fd_sc_hs__clkbuf_8_3/X
+ sky130_fd_sc_hs__clkbuf_16_37/a_114_74# sky130_fd_sc_hs__clkbuf_16
Xsky130_fd_sc_hs__clkbuf_16_48 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__einvp_2_97/A
+ sky130_fd_sc_hs__inv_4_9/Y sky130_fd_sc_hs__clkbuf_16_49/a_114_74# sky130_fd_sc_hs__clkbuf_16
Xsky130_fd_sc_hs__clkbuf_16_59 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__o21ai_4_1/A1
+ sky130_fd_sc_hs__clkbuf_16_93/X sky130_fd_sc_hs__clkbuf_16_59/a_114_74# sky130_fd_sc_hs__clkbuf_16
Xsky130_fd_sc_hs__clkbuf_16_103 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__clkbuf_8_67/A
+ sky130_fd_sc_hs__clkbuf_4_127/X sky130_fd_sc_hs__clkbuf_16_103/a_114_74# sky130_fd_sc_hs__clkbuf_16
Xsky130_fd_sc_hs__clkbuf_16_114 DVSS: DVDD: DVDD: DVSS: osc_core_1/pi4_l[1] pi4_con[1]
+ sky130_fd_sc_hs__clkbuf_16_115/a_114_74# sky130_fd_sc_hs__clkbuf_16
Xsky130_fd_sc_hs__clkbuf_16_125 DVSS: DVDD: DVDD: DVSS: osc_core_1/pi5_l[2] sky130_fd_sc_hs__clkbuf_4_131/X
+ sky130_fd_sc_hs__clkbuf_16_125/a_114_74# sky130_fd_sc_hs__clkbuf_16
Xsky130_fd_sc_hs__clkbuf_4_103 DVSS: DVDD: DVDD: DVSS: con_perb[1] osc_core_1/con_perb_5[1]
+ sky130_fd_sc_hs__clkbuf_4_103/a_83_270# sky130_fd_sc_hs__clkbuf_4
Xsky130_fd_sc_hs__clkbuf_4_114 DVSS: DVDD: DVDD: DVSS: CTL_BUF_P[5] sky130_fd_sc_hs__clkbuf_4_115/X
+ sky130_fd_sc_hs__clkbuf_4_115/a_83_270# sky130_fd_sc_hs__clkbuf_4
Xsky130_fd_sc_hs__clkbuf_4_125 DVSS: DVDD: DVDD: DVSS: pi5_con[1] sky130_fd_sc_hs__clkbuf_4_125/X
+ sky130_fd_sc_hs__clkbuf_4_125/a_83_270# sky130_fd_sc_hs__clkbuf_4
Xsky130_fd_sc_hs__clkbuf_4_136 DVSS: DVDD: DVDD: DVSS: pi5_con[3] sky130_fd_sc_hs__clkbuf_4_137/X
+ sky130_fd_sc_hs__clkbuf_4_137/a_83_270# sky130_fd_sc_hs__clkbuf_4
Xsky130_fd_sc_hs__o21ai_2_5 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__inv_4_13/Y sky130_fd_sc_hs__o21ai_2_9/A2
+ sky130_fd_sc_hs__nand2_2_9/B sky130_fd_sc_hs__o21ai_2_5/Y sky130_fd_sc_hs__o21ai_2_5/a_116_368#
+ sky130_fd_sc_hs__o21ai_2_5/a_27_74# sky130_fd_sc_hs__o21ai_2
Xsky130_fd_sc_hs__clkbuf_4_10 DVSS: DVDD: DVDD: DVSS: manual_control_osc[12] sky130_fd_sc_hs__clkbuf_8_15/A
+ sky130_fd_sc_hs__clkbuf_4_11/a_83_270# sky130_fd_sc_hs__clkbuf_4
Xsky130_fd_sc_hs__clkbuf_4_21 DVSS: DVDD: DVDD: DVSS: pi1_con[2] sky130_fd_sc_hs__clkbuf_4_21/X
+ sky130_fd_sc_hs__clkbuf_4_21/a_83_270# sky130_fd_sc_hs__clkbuf_4
Xsky130_fd_sc_hs__clkbuf_4_32 DVSS: DVDD: DVDD: DVSS: manual_control_osc[5] sky130_fd_sc_hs__clkbuf_8_23/A
+ sky130_fd_sc_hs__clkbuf_4_33/a_83_270# sky130_fd_sc_hs__clkbuf_4
Xsky130_fd_sc_hs__clkbuf_4_43 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__einvn_8_1/Z
+ qr_4t1_mux_top_1/clk_Q sky130_fd_sc_hs__clkbuf_4_43/a_83_270# sky130_fd_sc_hs__clkbuf_4
Xsky130_fd_sc_hs__clkbuf_4_54 DVSS: DVDD: DVDD: DVSS: fine_con_step_size[0] sky130_fd_sc_hs__clkbuf_4_55/X
+ sky130_fd_sc_hs__clkbuf_4_55/a_83_270# sky130_fd_sc_hs__clkbuf_4
Xsky130_fd_sc_hs__clkbuf_4_65 DVSS: DVDD: DVDD: DVSS: fine_control_avg_window_select[4]
+ sky130_fd_sc_hs__clkbuf_4_65/X sky130_fd_sc_hs__clkbuf_4_65/a_83_270# sky130_fd_sc_hs__clkbuf_4
Xsky130_fd_sc_hs__clkbuf_4_76 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__buf_2_89/X
+ sky130_fd_sc_hs__dlrtp_1_21/D sky130_fd_sc_hs__clkbuf_4_77/a_83_270# sky130_fd_sc_hs__clkbuf_4
Xsky130_fd_sc_hs__clkbuf_4_87 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__or2b_2_3/A
+ sky130_fd_sc_hs__o21ai_2_51/A1 sky130_fd_sc_hs__clkbuf_4_87/a_83_270# sky130_fd_sc_hs__clkbuf_4
Xsky130_fd_sc_hs__clkbuf_4_98 DVSS: DVDD: DVDD: DVSS: div_ratio_half[0] sky130_fd_sc_hs__clkbuf_4_99/X
+ sky130_fd_sc_hs__clkbuf_4_99/a_83_270# sky130_fd_sc_hs__clkbuf_4
Xsky130_fd_sc_hs__clkinv_8_13 DVSS: DVDD: DVDD: DVSS: prbs_generator_syn_9/out hr_16t4_mux_top_3/din[3]
+ sky130_fd_sc_hs__clkinv_8
Xsky130_fd_sc_hs__conb_1_100 DVSS: DVDD: DVDD: DVSS: prbs_generator_syn_13/eqn[22]
+ prbs_generator_syn_13/eqn[20] sky130_fd_sc_hs__conb_1_101/a_165_290# sky130_fd_sc_hs__conb_1_101/a_21_290#
+ sky130_fd_sc_hs__conb_1
Xsky130_fd_sc_hs__conb_1_111 DVSS: DVDD: DVDD: DVSS: prbs_generator_syn_15/eqn[13]
+ sky130_fd_sc_hs__conb_1_111/HI sky130_fd_sc_hs__conb_1_111/a_165_290# sky130_fd_sc_hs__conb_1_111/a_21_290#
+ sky130_fd_sc_hs__conb_1
Xsky130_fd_sc_hs__conb_1_122 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__conb_1_123/LO
+ sky130_fd_sc_hs__conb_1_123/HI sky130_fd_sc_hs__conb_1_123/a_165_290# sky130_fd_sc_hs__conb_1_123/a_21_290#
+ sky130_fd_sc_hs__conb_1
Xsky130_fd_sc_hs__conb_1_133 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__conb_1_133/LO
+ sky130_fd_sc_hs__conb_1_133/HI sky130_fd_sc_hs__conb_1_133/a_165_290# sky130_fd_sc_hs__conb_1_133/a_21_290#
+ sky130_fd_sc_hs__conb_1
Xsky130_fd_sc_hs__conb_1_144 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__conb_1_145/LO
+ sky130_fd_sc_hs__conb_1_145/HI sky130_fd_sc_hs__conb_1_145/a_165_290# sky130_fd_sc_hs__conb_1_145/a_21_290#
+ sky130_fd_sc_hs__conb_1
Xsky130_fd_sc_hs__conb_1_155 DVSS: DVDD: DVDD: DVSS: prbs_generator_syn_17/eqn[22]
+ prbs_generator_syn_17/eqn[20] sky130_fd_sc_hs__conb_1_155/a_165_290# sky130_fd_sc_hs__conb_1_155/a_21_290#
+ sky130_fd_sc_hs__conb_1
Xsky130_fd_sc_hs__conb_1_166 DVSS: DVDD: DVDD: DVSS: prbs_generator_syn_21/eqn[9]
+ sky130_fd_sc_hs__conb_1_167/HI sky130_fd_sc_hs__conb_1_167/a_165_290# sky130_fd_sc_hs__conb_1_167/a_21_290#
+ sky130_fd_sc_hs__conb_1
Xsky130_fd_sc_hs__conb_1_177 DVSS: DVDD: DVDD: DVSS: prbs_generator_syn_21/eqn[0]
+ sky130_fd_sc_hs__conb_1_177/HI sky130_fd_sc_hs__conb_1_177/a_165_290# sky130_fd_sc_hs__conb_1_177/a_21_290#
+ sky130_fd_sc_hs__conb_1
Xsky130_fd_sc_hs__conb_1_188 DVSS: DVDD: DVDD: DVSS: prbs_generator_syn_29/eqn[22]
+ prbs_generator_syn_29/eqn[20] sky130_fd_sc_hs__conb_1_189/a_165_290# sky130_fd_sc_hs__conb_1_189/a_21_290#
+ sky130_fd_sc_hs__conb_1
Xsky130_fd_sc_hs__conb_1_199 DVSS: DVDD: DVDD: DVSS: prbs_generator_syn_19/eqn[2]
+ prbs_generator_syn_19/eqn[1] sky130_fd_sc_hs__conb_1_199/a_165_290# sky130_fd_sc_hs__conb_1_199/a_21_290#
+ sky130_fd_sc_hs__conb_1
Xsky130_fd_sc_hs__nand2_8_0 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__nor4_2_1/C sky130_fd_sc_hs__nor4_2_1/A
+ sky130_fd_sc_hs__nand2_8_1/Y sky130_fd_sc_hs__nand2_8_1/a_27_74# sky130_fd_sc_hs__nand2_8
Xsky130_fd_sc_hs__einvp_2_100 DVSS: DVDD: DVDD: DVSS: dout_p sky130_fd_sc_hs__einvp_2_97/A
+ sky130_fd_sc_hs__dlrtp_1_75/Q sky130_fd_sc_hs__einvp_2_101/a_263_323# sky130_fd_sc_hs__einvp_2_101/a_36_74#
+ sky130_fd_sc_hs__einvp_2_101/a_27_368# sky130_fd_sc_hs__einvp_2
Xsky130_fd_sc_hs__einvp_2_111 DVSS: DVDD: DVDD: DVSS: dout_n sky130_fd_sc_hs__einvp_2_9/A
+ sky130_fd_sc_hs__dlrtp_1_97/Q sky130_fd_sc_hs__einvp_2_111/a_263_323# sky130_fd_sc_hs__einvp_2_111/a_36_74#
+ sky130_fd_sc_hs__einvp_2_111/a_27_368# sky130_fd_sc_hs__einvp_2
Xsky130_fd_sc_hs__einvp_2_122 DVSS: DVDD: DVDD: DVSS: dout_n sky130_fd_sc_hs__buf_8_1/X
+ sky130_fd_sc_hs__dlrtp_1_119/Q sky130_fd_sc_hs__einvp_2_123/a_263_323# sky130_fd_sc_hs__einvp_2_123/a_36_74#
+ sky130_fd_sc_hs__einvp_2_123/a_27_368# sky130_fd_sc_hs__einvp_2
Xsky130_fd_sc_hs__einvp_2_133 DVSS: DVDD: DVDD: DVSS: dout_p sky130_fd_sc_hs__einvp_2_99/A
+ sky130_fd_sc_hs__dlrtp_1_131/Q sky130_fd_sc_hs__einvp_2_133/a_263_323# sky130_fd_sc_hs__einvp_2_133/a_36_74#
+ sky130_fd_sc_hs__einvp_2_133/a_27_368# sky130_fd_sc_hs__einvp_2
Xsky130_fd_sc_hs__einvp_2_144 DVSS: DVDD: DVDD: DVSS: dout_p sky130_fd_sc_hs__einvp_2_99/A
+ sky130_fd_sc_hs__dlrtp_1_147/Q sky130_fd_sc_hs__einvp_2_145/a_263_323# sky130_fd_sc_hs__einvp_2_145/a_36_74#
+ sky130_fd_sc_hs__einvp_2_145/a_27_368# sky130_fd_sc_hs__einvp_2
Xsky130_fd_sc_hs__einvp_2_155 DVSS: DVDD: DVDD: DVSS: dout_p sky130_fd_sc_hs__einvp_2_99/A
+ sky130_fd_sc_hs__buf_2_161/X sky130_fd_sc_hs__einvp_2_155/a_263_323# sky130_fd_sc_hs__einvp_2_155/a_36_74#
+ sky130_fd_sc_hs__einvp_2_155/a_27_368# sky130_fd_sc_hs__einvp_2
Xsky130_fd_sc_hs__clkbuf_16_16 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__clkbuf_16_17/X
+ sky130_fd_sc_hs__clkbuf_4_27/X sky130_fd_sc_hs__clkbuf_16_17/a_114_74# sky130_fd_sc_hs__clkbuf_16
Xsky130_fd_sc_hs__clkbuf_16_27 DVSS: DVDD: DVDD: DVSS: osc_core_1/pi3_l[2] sky130_fd_sc_hs__clkbuf_8_7/X
+ sky130_fd_sc_hs__clkbuf_16_27/a_114_74# sky130_fd_sc_hs__clkbuf_16
Xsky130_fd_sc_hs__clkbuf_16_38 DVSS: DVDD: DVDD: DVSS: osc_core_1/pi2_l[1] sky130_fd_sc_hs__clkbuf_16_3/X
+ sky130_fd_sc_hs__clkbuf_16_39/a_114_74# sky130_fd_sc_hs__clkbuf_16
Xsky130_fd_sc_hs__clkbuf_16_49 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__einvp_2_97/A
+ sky130_fd_sc_hs__inv_4_9/Y sky130_fd_sc_hs__clkbuf_16_49/a_114_74# sky130_fd_sc_hs__clkbuf_16
Xsky130_fd_sc_hs__clkbuf_16_0 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__clkbuf_16_1/X
+ pi3_con[0] sky130_fd_sc_hs__clkbuf_16_1/a_114_74# sky130_fd_sc_hs__clkbuf_16
Xsky130_fd_sc_hs__clkbuf_16_104 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__clkbuf_16_63/A
+ sky130_fd_sc_hs__clkbuf_4_119/X sky130_fd_sc_hs__clkbuf_16_105/a_114_74# sky130_fd_sc_hs__clkbuf_16
Xsky130_fd_sc_hs__clkbuf_16_115 DVSS: DVDD: DVDD: DVSS: osc_core_1/pi4_l[1] pi4_con[1]
+ sky130_fd_sc_hs__clkbuf_16_115/a_114_74# sky130_fd_sc_hs__clkbuf_16
Xsky130_fd_sc_hs__clkbuf_16_126 DVSS: DVDD: DVDD: DVSS: osc_core_1/pi5_l[1] sky130_fd_sc_hs__clkbuf_4_125/X
+ sky130_fd_sc_hs__clkbuf_16_127/a_114_74# sky130_fd_sc_hs__clkbuf_16
Xsky130_fd_sc_hs__clkbuf_4_104 DVSS: DVDD: DVDD: DVSS: con_perb[0] osc_core_1/con_perb_5[0]
+ sky130_fd_sc_hs__clkbuf_4_105/a_83_270# sky130_fd_sc_hs__clkbuf_4
Xsky130_fd_sc_hs__clkbuf_4_115 DVSS: DVDD: DVDD: DVSS: CTL_BUF_P[5] sky130_fd_sc_hs__clkbuf_4_115/X
+ sky130_fd_sc_hs__clkbuf_4_115/a_83_270# sky130_fd_sc_hs__clkbuf_4
Xsky130_fd_sc_hs__clkbuf_4_126 DVSS: DVDD: DVDD: DVSS: CTL_BUF_N[2] sky130_fd_sc_hs__clkbuf_4_127/X
+ sky130_fd_sc_hs__clkbuf_4_127/a_83_270# sky130_fd_sc_hs__clkbuf_4
Xsky130_fd_sc_hs__clkbuf_4_137 DVSS: DVDD: DVDD: DVSS: pi5_con[3] sky130_fd_sc_hs__clkbuf_4_137/X
+ sky130_fd_sc_hs__clkbuf_4_137/a_83_270# sky130_fd_sc_hs__clkbuf_4
Xsky130_fd_sc_hs__o21ai_2_6 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__inv_4_11/Y sky130_fd_sc_hs__nand2_2_3/B
+ sky130_fd_sc_hs__o21ai_2_9/A2 sky130_fd_sc_hs__buf_2_45/A sky130_fd_sc_hs__o21ai_2_7/a_116_368#
+ sky130_fd_sc_hs__o21ai_2_7/a_27_74# sky130_fd_sc_hs__o21ai_2
Xsky130_fd_sc_hs__clkbuf_4_11 DVSS: DVDD: DVDD: DVSS: manual_control_osc[12] sky130_fd_sc_hs__clkbuf_8_15/A
+ sky130_fd_sc_hs__clkbuf_4_11/a_83_270# sky130_fd_sc_hs__clkbuf_4
Xsky130_fd_sc_hs__clkbuf_4_22 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__buf_2_5/X sky130_fd_sc_hs__clkbuf_8_21/A
+ sky130_fd_sc_hs__clkbuf_4_23/a_83_270# sky130_fd_sc_hs__clkbuf_4
Xsky130_fd_sc_hs__clkbuf_4_33 DVSS: DVDD: DVDD: DVSS: manual_control_osc[5] sky130_fd_sc_hs__clkbuf_8_23/A
+ sky130_fd_sc_hs__clkbuf_4_33/a_83_270# sky130_fd_sc_hs__clkbuf_4
Xsky130_fd_sc_hs__clkbuf_4_44 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__buf_2_13/X
+ sky130_fd_sc_hs__clkbuf_8_31/A sky130_fd_sc_hs__clkbuf_4_45/a_83_270# sky130_fd_sc_hs__clkbuf_4
Xsky130_fd_sc_hs__clkbuf_4_55 DVSS: DVDD: DVDD: DVSS: fine_con_step_size[0] sky130_fd_sc_hs__clkbuf_4_55/X
+ sky130_fd_sc_hs__clkbuf_4_55/a_83_270# sky130_fd_sc_hs__clkbuf_4
Xsky130_fd_sc_hs__clkbuf_4_66 DVSS: DVDD: DVDD: DVSS: fine_control_avg_window_select[0]
+ sky130_fd_sc_hs__clkbuf_4_67/X sky130_fd_sc_hs__clkbuf_4_67/a_83_270# sky130_fd_sc_hs__clkbuf_4
Xsky130_fd_sc_hs__clkbuf_4_77 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__buf_2_89/X
+ sky130_fd_sc_hs__dlrtp_1_21/D sky130_fd_sc_hs__clkbuf_4_77/a_83_270# sky130_fd_sc_hs__clkbuf_4
Xsky130_fd_sc_hs__clkbuf_4_88 DVSS: DVDD: DVDD: DVSS: div_ratio_half[5] sky130_fd_sc_hs__clkbuf_4_89/X
+ sky130_fd_sc_hs__clkbuf_4_89/a_83_270# sky130_fd_sc_hs__clkbuf_4
Xsky130_fd_sc_hs__clkbuf_4_99 DVSS: DVDD: DVDD: DVSS: div_ratio_half[0] sky130_fd_sc_hs__clkbuf_4_99/X
+ sky130_fd_sc_hs__clkbuf_4_99/a_83_270# sky130_fd_sc_hs__clkbuf_4
Xsky130_fd_sc_hs__clkinv_8_14 DVSS: DVDD: DVDD: DVSS: osc_core_1/glob_en sky130_fd_sc_hs__clkinv_8_15/Y
+ sky130_fd_sc_hs__clkinv_8
Xsky130_fd_sc_hs__buf_8_0 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__buf_8_1/X sky130_fd_sc_hs__buf_8_1/A
+ sky130_fd_sc_hs__buf_8_1/a_27_74# sky130_fd_sc_hs__buf_8
Xsky130_fd_sc_hs__inv_8_0 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__or4_2_1/A sky130_fd_sc_hs__inv_8_1/Y
+ sky130_fd_sc_hs__inv_8
Xsky130_fd_sc_hs__conb_1_101 DVSS: DVDD: DVDD: DVSS: prbs_generator_syn_13/eqn[22]
+ prbs_generator_syn_13/eqn[20] sky130_fd_sc_hs__conb_1_101/a_165_290# sky130_fd_sc_hs__conb_1_101/a_21_290#
+ sky130_fd_sc_hs__conb_1
Xsky130_fd_sc_hs__conb_1_112 DVSS: DVDD: DVDD: DVSS: prbs_generator_syn_15/eqn[9]
+ sky130_fd_sc_hs__conb_1_113/HI sky130_fd_sc_hs__conb_1_113/a_165_290# sky130_fd_sc_hs__conb_1_113/a_21_290#
+ sky130_fd_sc_hs__conb_1
Xsky130_fd_sc_hs__conb_1_123 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__conb_1_123/LO
+ sky130_fd_sc_hs__conb_1_123/HI sky130_fd_sc_hs__conb_1_123/a_165_290# sky130_fd_sc_hs__conb_1_123/a_21_290#
+ sky130_fd_sc_hs__conb_1
Xsky130_fd_sc_hs__conb_1_134 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__conb_1_135/LO
+ sky130_fd_sc_hs__conb_1_135/HI sky130_fd_sc_hs__conb_1_135/a_165_290# sky130_fd_sc_hs__conb_1_135/a_21_290#
+ sky130_fd_sc_hs__conb_1
Xsky130_fd_sc_hs__conb_1_145 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__conb_1_145/LO
+ sky130_fd_sc_hs__conb_1_145/HI sky130_fd_sc_hs__conb_1_145/a_165_290# sky130_fd_sc_hs__conb_1_145/a_21_290#
+ sky130_fd_sc_hs__conb_1
Xsky130_fd_sc_hs__conb_1_156 DVSS: DVDD: DVDD: DVSS: prbs_generator_syn_17/eqn[30]
+ sky130_fd_sc_hs__conb_1_157/HI sky130_fd_sc_hs__conb_1_157/a_165_290# sky130_fd_sc_hs__conb_1_157/a_21_290#
+ sky130_fd_sc_hs__conb_1
Xsky130_fd_sc_hs__conb_1_167 DVSS: DVDD: DVDD: DVSS: prbs_generator_syn_21/eqn[9]
+ sky130_fd_sc_hs__conb_1_167/HI sky130_fd_sc_hs__conb_1_167/a_165_290# sky130_fd_sc_hs__conb_1_167/a_21_290#
+ sky130_fd_sc_hs__conb_1
Xsky130_fd_sc_hs__conb_1_178 DVSS: DVDD: DVDD: DVSS: prbs_generator_syn_23/eqn[22]
+ prbs_generator_syn_23/eqn[20] sky130_fd_sc_hs__conb_1_179/a_165_290# sky130_fd_sc_hs__conb_1_179/a_21_290#
+ sky130_fd_sc_hs__conb_1
Xsky130_fd_sc_hs__conb_1_189 DVSS: DVDD: DVDD: DVSS: prbs_generator_syn_29/eqn[22]
+ prbs_generator_syn_29/eqn[20] sky130_fd_sc_hs__conb_1_189/a_165_290# sky130_fd_sc_hs__conb_1_189/a_21_290#
+ sky130_fd_sc_hs__conb_1
Xsky130_fd_sc_hs__nand2_8_1 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__nor4_2_1/C sky130_fd_sc_hs__nor4_2_1/A
+ sky130_fd_sc_hs__nand2_8_1/Y sky130_fd_sc_hs__nand2_8_1/a_27_74# sky130_fd_sc_hs__nand2_8
Xsky130_fd_sc_hs__einvn_2_0 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__clkinv_8_15/Y
+ osc_core_1/p1 sky130_fd_sc_hs__einvn_2_1/Z sky130_fd_sc_hs__einvn_2_1/a_227_368#
+ sky130_fd_sc_hs__einvn_2_1/a_231_74# sky130_fd_sc_hs__einvn_2_1/a_115_464# sky130_fd_sc_hs__einvn_2
Xsky130_fd_sc_hs__einvp_2_101 DVSS: DVDD: DVDD: DVSS: dout_p sky130_fd_sc_hs__einvp_2_97/A
+ sky130_fd_sc_hs__dlrtp_1_75/Q sky130_fd_sc_hs__einvp_2_101/a_263_323# sky130_fd_sc_hs__einvp_2_101/a_36_74#
+ sky130_fd_sc_hs__einvp_2_101/a_27_368# sky130_fd_sc_hs__einvp_2
Xsky130_fd_sc_hs__einvp_2_112 DVSS: DVDD: DVDD: DVSS: dout_n sky130_fd_sc_hs__einvp_2_9/A
+ sky130_fd_sc_hs__dlrtp_1_103/Q sky130_fd_sc_hs__einvp_2_113/a_263_323# sky130_fd_sc_hs__einvp_2_113/a_36_74#
+ sky130_fd_sc_hs__einvp_2_113/a_27_368# sky130_fd_sc_hs__einvp_2
Xsky130_fd_sc_hs__einvp_2_123 DVSS: DVDD: DVDD: DVSS: dout_n sky130_fd_sc_hs__buf_8_1/X
+ sky130_fd_sc_hs__dlrtp_1_119/Q sky130_fd_sc_hs__einvp_2_123/a_263_323# sky130_fd_sc_hs__einvp_2_123/a_36_74#
+ sky130_fd_sc_hs__einvp_2_123/a_27_368# sky130_fd_sc_hs__einvp_2
Xsky130_fd_sc_hs__einvp_2_134 DVSS: DVDD: DVDD: DVSS: dout_p sky130_fd_sc_hs__einvp_2_99/A
+ sky130_fd_sc_hs__dlrtp_1_135/Q sky130_fd_sc_hs__einvp_2_135/a_263_323# sky130_fd_sc_hs__einvp_2_135/a_36_74#
+ sky130_fd_sc_hs__einvp_2_135/a_27_368# sky130_fd_sc_hs__einvp_2
Xsky130_fd_sc_hs__einvp_2_145 DVSS: DVDD: DVDD: DVSS: dout_p sky130_fd_sc_hs__einvp_2_99/A
+ sky130_fd_sc_hs__dlrtp_1_147/Q sky130_fd_sc_hs__einvp_2_145/a_263_323# sky130_fd_sc_hs__einvp_2_145/a_36_74#
+ sky130_fd_sc_hs__einvp_2_145/a_27_368# sky130_fd_sc_hs__einvp_2
Xsky130_fd_sc_hs__einvp_2_156 DVSS: DVDD: DVDD: DVSS: dout_p sky130_fd_sc_hs__einvp_2_97/A
+ sky130_fd_sc_hs__dlrtp_1_153/Q sky130_fd_sc_hs__einvp_2_157/a_263_323# sky130_fd_sc_hs__einvp_2_157/a_36_74#
+ sky130_fd_sc_hs__einvp_2_157/a_27_368# sky130_fd_sc_hs__einvp_2
Xsky130_fd_sc_hs__clkbuf_16_17 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__clkbuf_16_17/X
+ sky130_fd_sc_hs__clkbuf_4_27/X sky130_fd_sc_hs__clkbuf_16_17/a_114_74# sky130_fd_sc_hs__clkbuf_16
Xsky130_fd_sc_hs__clkbuf_16_28 DVSS: DVDD: DVDD: DVSS: osc_core_1/ref_clk ref_clk_ext_p
+ sky130_fd_sc_hs__clkbuf_16_29/a_114_74# sky130_fd_sc_hs__clkbuf_16
Xsky130_fd_sc_hs__clkbuf_16_39 DVSS: DVDD: DVDD: DVSS: osc_core_1/pi2_l[1] sky130_fd_sc_hs__clkbuf_16_3/X
+ sky130_fd_sc_hs__clkbuf_16_39/a_114_74# sky130_fd_sc_hs__clkbuf_16
Xsky130_fd_sc_hs__clkbuf_16_1 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__clkbuf_16_1/X
+ pi3_con[0] sky130_fd_sc_hs__clkbuf_16_1/a_114_74# sky130_fd_sc_hs__clkbuf_16
Xsky130_fd_sc_hs__clkbuf_16_105 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__clkbuf_16_63/A
+ sky130_fd_sc_hs__clkbuf_4_119/X sky130_fd_sc_hs__clkbuf_16_105/a_114_74# sky130_fd_sc_hs__clkbuf_16
Xsky130_fd_sc_hs__clkbuf_16_116 DVSS: DVDD: DVDD: DVSS: osc_core_1/pi4_l[2] pi4_con[2]
+ sky130_fd_sc_hs__clkbuf_16_117/a_114_74# sky130_fd_sc_hs__clkbuf_16
Xsky130_fd_sc_hs__clkbuf_16_127 DVSS: DVDD: DVDD: DVSS: osc_core_1/pi5_l[1] sky130_fd_sc_hs__clkbuf_4_125/X
+ sky130_fd_sc_hs__clkbuf_16_127/a_114_74# sky130_fd_sc_hs__clkbuf_16
Xsky130_fd_sc_hs__clkbuf_4_105 DVSS: DVDD: DVDD: DVSS: con_perb[0] osc_core_1/con_perb_5[0]
+ sky130_fd_sc_hs__clkbuf_4_105/a_83_270# sky130_fd_sc_hs__clkbuf_4
Xsky130_fd_sc_hs__clkbuf_4_116 DVSS: DVDD: DVDD: DVSS: CTL_BUF_P[3] sky130_fd_sc_hs__clkbuf_8_75/A
+ sky130_fd_sc_hs__clkbuf_4_117/a_83_270# sky130_fd_sc_hs__clkbuf_4
Xsky130_fd_sc_hs__clkbuf_4_127 DVSS: DVDD: DVDD: DVSS: CTL_BUF_N[2] sky130_fd_sc_hs__clkbuf_4_127/X
+ sky130_fd_sc_hs__clkbuf_4_127/a_83_270# sky130_fd_sc_hs__clkbuf_4
Xsky130_fd_sc_hs__o21ai_2_7 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__inv_4_11/Y sky130_fd_sc_hs__nand2_2_3/B
+ sky130_fd_sc_hs__o21ai_2_9/A2 sky130_fd_sc_hs__buf_2_45/A sky130_fd_sc_hs__o21ai_2_7/a_116_368#
+ sky130_fd_sc_hs__o21ai_2_7/a_27_74# sky130_fd_sc_hs__o21ai_2
Xsky130_fd_sc_hs__clkbuf_4_12 DVSS: DVDD: DVDD: DVSS: pi1_con[3] sky130_fd_sc_hs__clkbuf_4_13/X
+ sky130_fd_sc_hs__clkbuf_4_13/a_83_270# sky130_fd_sc_hs__clkbuf_4
Xsky130_fd_sc_hs__clkbuf_4_23 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__buf_2_5/X sky130_fd_sc_hs__clkbuf_8_21/A
+ sky130_fd_sc_hs__clkbuf_4_23/a_83_270# sky130_fd_sc_hs__clkbuf_4
Xsky130_fd_sc_hs__clkbuf_4_34 DVSS: DVDD: DVDD: DVSS: manual_control_osc[4] sky130_fd_sc_hs__clkbuf_8_25/A
+ sky130_fd_sc_hs__clkbuf_4_35/a_83_270# sky130_fd_sc_hs__clkbuf_4
Xsky130_fd_sc_hs__clkbuf_4_45 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__buf_2_13/X
+ sky130_fd_sc_hs__clkbuf_8_31/A sky130_fd_sc_hs__clkbuf_4_45/a_83_270# sky130_fd_sc_hs__clkbuf_4
Xsky130_fd_sc_hs__clkbuf_4_56 DVSS: DVDD: DVDD: DVSS: fine_con_step_size[2] sky130_fd_sc_hs__clkbuf_4_57/X
+ sky130_fd_sc_hs__clkbuf_4_57/a_83_270# sky130_fd_sc_hs__clkbuf_4
Xsky130_fd_sc_hs__clkbuf_4_67 DVSS: DVDD: DVDD: DVSS: fine_control_avg_window_select[0]
+ sky130_fd_sc_hs__clkbuf_4_67/X sky130_fd_sc_hs__clkbuf_4_67/a_83_270# sky130_fd_sc_hs__clkbuf_4
Xsky130_fd_sc_hs__clkbuf_4_78 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__nand2_2_17/Y
+ sky130_fd_sc_hs__inv_4_21/A sky130_fd_sc_hs__clkbuf_4_79/a_83_270# sky130_fd_sc_hs__clkbuf_4
Xsky130_fd_sc_hs__clkbuf_4_89 DVSS: DVDD: DVDD: DVSS: div_ratio_half[5] sky130_fd_sc_hs__clkbuf_4_89/X
+ sky130_fd_sc_hs__clkbuf_4_89/a_83_270# sky130_fd_sc_hs__clkbuf_4
Xsky130_fd_sc_hs__clkinv_8_15 DVSS: DVDD: DVDD: DVSS: osc_core_1/glob_en sky130_fd_sc_hs__clkinv_8_15/Y
+ sky130_fd_sc_hs__clkinv_8
Xsky130_fd_sc_hs__buf_8_1 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__buf_8_1/X sky130_fd_sc_hs__buf_8_1/A
+ sky130_fd_sc_hs__buf_8_1/a_27_74# sky130_fd_sc_hs__buf_8
Xsky130_fd_sc_hs__inv_8_1 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__or4_2_1/A sky130_fd_sc_hs__inv_8_1/Y
+ sky130_fd_sc_hs__inv_8
Xsky130_fd_sc_hs__conb_1_102 DVSS: DVDD: DVDD: DVSS: prbs_generator_syn_13/eqn[2]
+ prbs_generator_syn_13/eqn[1] sky130_fd_sc_hs__conb_1_103/a_165_290# sky130_fd_sc_hs__conb_1_103/a_21_290#
+ sky130_fd_sc_hs__conb_1
Xsky130_fd_sc_hs__conb_1_113 DVSS: DVDD: DVDD: DVSS: prbs_generator_syn_15/eqn[9]
+ sky130_fd_sc_hs__conb_1_113/HI sky130_fd_sc_hs__conb_1_113/a_165_290# sky130_fd_sc_hs__conb_1_113/a_21_290#
+ sky130_fd_sc_hs__conb_1
Xsky130_fd_sc_hs__conb_1_124 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__conb_1_125/LO
+ sky130_fd_sc_hs__conb_1_125/HI sky130_fd_sc_hs__conb_1_125/a_165_290# sky130_fd_sc_hs__conb_1_125/a_21_290#
+ sky130_fd_sc_hs__conb_1
Xsky130_fd_sc_hs__conb_1_135 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__conb_1_135/LO
+ sky130_fd_sc_hs__conb_1_135/HI sky130_fd_sc_hs__conb_1_135/a_165_290# sky130_fd_sc_hs__conb_1_135/a_21_290#
+ sky130_fd_sc_hs__conb_1
Xsky130_fd_sc_hs__conb_1_146 DVSS: DVDD: DVDD: DVSS: prbs_generator_syn_17/eqn[13]
+ sky130_fd_sc_hs__conb_1_147/HI sky130_fd_sc_hs__conb_1_147/a_165_290# sky130_fd_sc_hs__conb_1_147/a_21_290#
+ sky130_fd_sc_hs__conb_1
Xsky130_fd_sc_hs__conb_1_157 DVSS: DVDD: DVDD: DVSS: prbs_generator_syn_17/eqn[30]
+ sky130_fd_sc_hs__conb_1_157/HI sky130_fd_sc_hs__conb_1_157/a_165_290# sky130_fd_sc_hs__conb_1_157/a_21_290#
+ sky130_fd_sc_hs__conb_1
Xsky130_fd_sc_hs__conb_1_168 DVSS: DVDD: DVDD: DVSS: prbs_generator_syn_21/eqn[22]
+ prbs_generator_syn_21/eqn[20] sky130_fd_sc_hs__conb_1_169/a_165_290# sky130_fd_sc_hs__conb_1_169/a_21_290#
+ sky130_fd_sc_hs__conb_1
Xsky130_fd_sc_hs__conb_1_179 DVSS: DVDD: DVDD: DVSS: prbs_generator_syn_23/eqn[22]
+ prbs_generator_syn_23/eqn[20] sky130_fd_sc_hs__conb_1_179/a_165_290# sky130_fd_sc_hs__conb_1_179/a_21_290#
+ sky130_fd_sc_hs__conb_1
Xsky130_fd_sc_hs__nand2_8_2 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__or4_2_1/C sky130_fd_sc_hs__or4_2_1/B
+ sky130_fd_sc_hs__or2b_4_5/A sky130_fd_sc_hs__nand2_8_3/a_27_74# sky130_fd_sc_hs__nand2_8
Xsky130_fd_sc_hs__einvn_2_1 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__clkinv_8_15/Y
+ osc_core_1/p1 sky130_fd_sc_hs__einvn_2_1/Z sky130_fd_sc_hs__einvn_2_1/a_227_368#
+ sky130_fd_sc_hs__einvn_2_1/a_231_74# sky130_fd_sc_hs__einvn_2_1/a_115_464# sky130_fd_sc_hs__einvn_2
Xsky130_fd_sc_hs__einvp_2_102 DVSS: DVDD: DVDD: DVSS: dout_p sky130_fd_sc_hs__einvp_2_97/A
+ sky130_fd_sc_hs__dlrtp_1_74/Q sky130_fd_sc_hs__einvp_2_103/a_263_323# sky130_fd_sc_hs__einvp_2_103/a_36_74#
+ sky130_fd_sc_hs__einvp_2_103/a_27_368# sky130_fd_sc_hs__einvp_2
Xsky130_fd_sc_hs__einvp_2_113 DVSS: DVDD: DVDD: DVSS: dout_n sky130_fd_sc_hs__einvp_2_9/A
+ sky130_fd_sc_hs__dlrtp_1_103/Q sky130_fd_sc_hs__einvp_2_113/a_263_323# sky130_fd_sc_hs__einvp_2_113/a_36_74#
+ sky130_fd_sc_hs__einvp_2_113/a_27_368# sky130_fd_sc_hs__einvp_2
Xsky130_fd_sc_hs__einvp_2_124 DVSS: DVDD: DVDD: DVSS: dout_n sky130_fd_sc_hs__buf_8_1/X
+ sky130_fd_sc_hs__dlrtp_1_121/Q sky130_fd_sc_hs__einvp_2_125/a_263_323# sky130_fd_sc_hs__einvp_2_125/a_36_74#
+ sky130_fd_sc_hs__einvp_2_125/a_27_368# sky130_fd_sc_hs__einvp_2
Xsky130_fd_sc_hs__einvp_2_135 DVSS: DVDD: DVDD: DVSS: dout_p sky130_fd_sc_hs__einvp_2_99/A
+ sky130_fd_sc_hs__dlrtp_1_135/Q sky130_fd_sc_hs__einvp_2_135/a_263_323# sky130_fd_sc_hs__einvp_2_135/a_36_74#
+ sky130_fd_sc_hs__einvp_2_135/a_27_368# sky130_fd_sc_hs__einvp_2
Xsky130_fd_sc_hs__einvp_2_146 DVSS: DVDD: DVDD: DVSS: dout_p sky130_fd_sc_hs__einvp_2_99/A
+ sky130_fd_sc_hs__dlrtp_1_149/Q sky130_fd_sc_hs__einvp_2_147/a_263_323# sky130_fd_sc_hs__einvp_2_147/a_36_74#
+ sky130_fd_sc_hs__einvp_2_147/a_27_368# sky130_fd_sc_hs__einvp_2
Xsky130_fd_sc_hs__einvp_2_157 DVSS: DVDD: DVDD: DVSS: dout_p sky130_fd_sc_hs__einvp_2_97/A
+ sky130_fd_sc_hs__dlrtp_1_153/Q sky130_fd_sc_hs__einvp_2_157/a_263_323# sky130_fd_sc_hs__einvp_2_157/a_36_74#
+ sky130_fd_sc_hs__einvp_2_157/a_27_368# sky130_fd_sc_hs__einvp_2
Xsky130_fd_sc_hs__clkbuf_16_18 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__clkbuf_16_19/X
+ sky130_fd_sc_hs__clkbuf_4_25/X sky130_fd_sc_hs__clkbuf_16_19/a_114_74# sky130_fd_sc_hs__clkbuf_16
Xsky130_fd_sc_hs__clkbuf_16_29 DVSS: DVDD: DVDD: DVSS: osc_core_1/ref_clk ref_clk_ext_p
+ sky130_fd_sc_hs__clkbuf_16_29/a_114_74# sky130_fd_sc_hs__clkbuf_16
Xsky130_fd_sc_hs__clkbuf_16_2 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__clkbuf_16_3/X
+ pi2_con[1] sky130_fd_sc_hs__clkbuf_16_3/a_114_74# sky130_fd_sc_hs__clkbuf_16
Xsky130_fd_sc_hs__clkbuf_16_106 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__einvp_8_3/TE
+ test_mux_clk_Q_select[0] sky130_fd_sc_hs__clkbuf_16_107/a_114_74# sky130_fd_sc_hs__clkbuf_16
Xsky130_fd_sc_hs__clkbuf_16_117 DVSS: DVDD: DVDD: DVSS: osc_core_1/pi4_l[2] pi4_con[2]
+ sky130_fd_sc_hs__clkbuf_16_117/a_114_74# sky130_fd_sc_hs__clkbuf_16
Xsky130_fd_sc_hs__clkbuf_16_128 DVSS: DVDD: DVDD: DVSS: osc_core_1/pi5_l[3] sky130_fd_sc_hs__clkbuf_4_137/X
+ sky130_fd_sc_hs__clkbuf_16_129/a_114_74# sky130_fd_sc_hs__clkbuf_16
Xsky130_fd_sc_hs__clkbuf_4_106 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__clkbuf_8_35/X
+ osc_core_1/pi2_l[0] sky130_fd_sc_hs__clkbuf_4_107/a_83_270# sky130_fd_sc_hs__clkbuf_4
Xsky130_fd_sc_hs__clkbuf_4_117 DVSS: DVDD: DVDD: DVSS: CTL_BUF_P[3] sky130_fd_sc_hs__clkbuf_8_75/A
+ sky130_fd_sc_hs__clkbuf_4_117/a_83_270# sky130_fd_sc_hs__clkbuf_4
Xsky130_fd_sc_hs__clkbuf_4_128 DVSS: DVDD: DVDD: DVSS: CTL_BUF_N[4] sky130_fd_sc_hs__clkbuf_8_77/A
+ sky130_fd_sc_hs__clkbuf_4_129/a_83_270# sky130_fd_sc_hs__clkbuf_4
Xsky130_fd_sc_hs__o21ai_2_8 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__inv_4_29/A sky130_fd_sc_hs__o21ai_2_9/A2
+ sky130_fd_sc_hs__nand2_2_5/B sky130_fd_sc_hs__buf_2_43/A sky130_fd_sc_hs__o21ai_2_9/a_116_368#
+ sky130_fd_sc_hs__o21ai_2_9/a_27_74# sky130_fd_sc_hs__o21ai_2
Xsky130_fd_sc_hs__clkbuf_4_13 DVSS: DVDD: DVDD: DVSS: pi1_con[3] sky130_fd_sc_hs__clkbuf_4_13/X
+ sky130_fd_sc_hs__clkbuf_4_13/a_83_270# sky130_fd_sc_hs__clkbuf_4
Xsky130_fd_sc_hs__clkbuf_4_24 DVSS: DVDD: DVDD: DVSS: manual_control_osc[7] sky130_fd_sc_hs__clkbuf_4_25/X
+ sky130_fd_sc_hs__clkbuf_4_25/a_83_270# sky130_fd_sc_hs__clkbuf_4
Xsky130_fd_sc_hs__clkbuf_4_35 DVSS: DVDD: DVDD: DVSS: manual_control_osc[4] sky130_fd_sc_hs__clkbuf_8_25/A
+ sky130_fd_sc_hs__clkbuf_4_35/a_83_270# sky130_fd_sc_hs__clkbuf_4
Xsky130_fd_sc_hs__clkbuf_8_0 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__clkbuf_8_1/X
+ pi2_con[3] sky130_fd_sc_hs__clkbuf_8_1/a_125_368# sky130_fd_sc_hs__clkbuf_8
Xsky130_fd_sc_hs__clkbuf_4_46 DVSS: DVDD: DVDD: DVSS: manual_control_osc[0] sky130_fd_sc_hs__clkbuf_4_47/X
+ sky130_fd_sc_hs__clkbuf_4_47/a_83_270# sky130_fd_sc_hs__clkbuf_4
Xsky130_fd_sc_hs__clkbuf_4_57 DVSS: DVDD: DVDD: DVSS: fine_con_step_size[2] sky130_fd_sc_hs__clkbuf_4_57/X
+ sky130_fd_sc_hs__clkbuf_4_57/a_83_270# sky130_fd_sc_hs__clkbuf_4
Xsky130_fd_sc_hs__clkbuf_4_68 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__inv_4_9/Y sky130_fd_sc_hs__einvp_2_65/A
+ sky130_fd_sc_hs__clkbuf_4_69/a_83_270# sky130_fd_sc_hs__clkbuf_4
Xsky130_fd_sc_hs__clkbuf_4_79 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__nand2_2_17/Y
+ sky130_fd_sc_hs__inv_4_21/A sky130_fd_sc_hs__clkbuf_4_79/a_83_270# sky130_fd_sc_hs__clkbuf_4
Xsky130_fd_sc_hs__clkinv_8_0 DVSS: DVDD: DVDD: DVSS: prbs_generator_syn_7/out hr_16t4_mux_top_3/din[11]
+ sky130_fd_sc_hs__clkinv_8
Xsky130_fd_sc_hs__clkinv_8_16 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__clkinv_8_19/Y
+ qr_4t1_mux_top_3/rst sky130_fd_sc_hs__clkinv_8
Xsky130_fd_sc_hs__buf_8_2 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__buf_8_3/X sky130_fd_sc_hs__buf_8_3/A
+ sky130_fd_sc_hs__buf_8_3/a_27_74# sky130_fd_sc_hs__buf_8
Xsky130_fd_sc_hs__conb_1_103 DVSS: DVDD: DVDD: DVSS: prbs_generator_syn_13/eqn[2]
+ prbs_generator_syn_13/eqn[1] sky130_fd_sc_hs__conb_1_103/a_165_290# sky130_fd_sc_hs__conb_1_103/a_21_290#
+ sky130_fd_sc_hs__conb_1
Xsky130_fd_sc_hs__conb_1_114 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__conb_1_115/LO
+ sky130_fd_sc_hs__conb_1_115/HI sky130_fd_sc_hs__conb_1_115/a_165_290# sky130_fd_sc_hs__conb_1_115/a_21_290#
+ sky130_fd_sc_hs__conb_1
Xsky130_fd_sc_hs__conb_1_125 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__conb_1_125/LO
+ sky130_fd_sc_hs__conb_1_125/HI sky130_fd_sc_hs__conb_1_125/a_165_290# sky130_fd_sc_hs__conb_1_125/a_21_290#
+ sky130_fd_sc_hs__conb_1
Xsky130_fd_sc_hs__conb_1_136 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__conb_1_137/LO
+ sky130_fd_sc_hs__conb_1_137/HI sky130_fd_sc_hs__conb_1_137/a_165_290# sky130_fd_sc_hs__conb_1_137/a_21_290#
+ sky130_fd_sc_hs__conb_1
Xsky130_fd_sc_hs__conb_1_147 DVSS: DVDD: DVDD: DVSS: prbs_generator_syn_17/eqn[13]
+ sky130_fd_sc_hs__conb_1_147/HI sky130_fd_sc_hs__conb_1_147/a_165_290# sky130_fd_sc_hs__conb_1_147/a_21_290#
+ sky130_fd_sc_hs__conb_1
Xsky130_fd_sc_hs__conb_1_158 DVSS: DVDD: DVDD: DVSS: prbs_generator_syn_17/eqn[31]
+ prbs_generator_syn_17/cke sky130_fd_sc_hs__conb_1_159/a_165_290# sky130_fd_sc_hs__conb_1_159/a_21_290#
+ sky130_fd_sc_hs__conb_1
Xsky130_fd_sc_hs__conb_1_169 DVSS: DVDD: DVDD: DVSS: prbs_generator_syn_21/eqn[22]
+ prbs_generator_syn_21/eqn[20] sky130_fd_sc_hs__conb_1_169/a_165_290# sky130_fd_sc_hs__conb_1_169/a_21_290#
+ sky130_fd_sc_hs__conb_1
Xsky130_fd_sc_hs__nand2_8_3 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__or4_2_1/C sky130_fd_sc_hs__or4_2_1/B
+ sky130_fd_sc_hs__or2b_4_5/A sky130_fd_sc_hs__nand2_8_3/a_27_74# sky130_fd_sc_hs__nand2_8
Xsky130_fd_sc_hs__or4_2_0 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__or4_2_1/X sky130_fd_sc_hs__or4_2_1/D
+ sky130_fd_sc_hs__or4_2_1/A sky130_fd_sc_hs__or4_2_1/B sky130_fd_sc_hs__or4_2_1/C
+ sky130_fd_sc_hs__or4_2_1/a_174_392# sky130_fd_sc_hs__or4_2_1/a_258_392# sky130_fd_sc_hs__or4_2_1/a_342_392#
+ sky130_fd_sc_hs__or4_2_1/a_85_392# sky130_fd_sc_hs__or4_2
Xsky130_fd_sc_hs__einvp_2_103 DVSS: DVDD: DVDD: DVSS: dout_p sky130_fd_sc_hs__einvp_2_97/A
+ sky130_fd_sc_hs__dlrtp_1_74/Q sky130_fd_sc_hs__einvp_2_103/a_263_323# sky130_fd_sc_hs__einvp_2_103/a_36_74#
+ sky130_fd_sc_hs__einvp_2_103/a_27_368# sky130_fd_sc_hs__einvp_2
Xsky130_fd_sc_hs__einvp_2_114 DVSS: DVDD: DVDD: DVSS: dout_n sky130_fd_sc_hs__einvp_2_9/A
+ sky130_fd_sc_hs__dlrtp_1_105/Q sky130_fd_sc_hs__einvp_2_115/a_263_323# sky130_fd_sc_hs__einvp_2_115/a_36_74#
+ sky130_fd_sc_hs__einvp_2_115/a_27_368# sky130_fd_sc_hs__einvp_2
Xsky130_fd_sc_hs__einvp_2_125 DVSS: DVDD: DVDD: DVSS: dout_n sky130_fd_sc_hs__buf_8_1/X
+ sky130_fd_sc_hs__dlrtp_1_121/Q sky130_fd_sc_hs__einvp_2_125/a_263_323# sky130_fd_sc_hs__einvp_2_125/a_36_74#
+ sky130_fd_sc_hs__einvp_2_125/a_27_368# sky130_fd_sc_hs__einvp_2
Xsky130_fd_sc_hs__einvp_2_136 DVSS: DVDD: DVDD: DVSS: dout_p sky130_fd_sc_hs__einvp_2_99/A
+ sky130_fd_sc_hs__dlrtp_1_55/Q sky130_fd_sc_hs__einvp_2_137/a_263_323# sky130_fd_sc_hs__einvp_2_137/a_36_74#
+ sky130_fd_sc_hs__einvp_2_137/a_27_368# sky130_fd_sc_hs__einvp_2
Xsky130_fd_sc_hs__einvp_2_147 DVSS: DVDD: DVDD: DVSS: dout_p sky130_fd_sc_hs__einvp_2_99/A
+ sky130_fd_sc_hs__dlrtp_1_149/Q sky130_fd_sc_hs__einvp_2_147/a_263_323# sky130_fd_sc_hs__einvp_2_147/a_36_74#
+ sky130_fd_sc_hs__einvp_2_147/a_27_368# sky130_fd_sc_hs__einvp_2
Xsky130_fd_sc_hs__einvp_2_158 DVSS: DVDD: DVDD: DVSS: dout_p sky130_fd_sc_hs__einvp_2_97/A
+ sky130_fd_sc_hs__dlrtp_1_151/Q sky130_fd_sc_hs__einvp_2_159/a_263_323# sky130_fd_sc_hs__einvp_2_159/a_36_74#
+ sky130_fd_sc_hs__einvp_2_159/a_27_368# sky130_fd_sc_hs__einvp_2
Xsky130_fd_sc_hs__clkbuf_16_19 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__clkbuf_16_19/X
+ sky130_fd_sc_hs__clkbuf_4_25/X sky130_fd_sc_hs__clkbuf_16_19/a_114_74# sky130_fd_sc_hs__clkbuf_16
Xsky130_fd_sc_hs__clkbuf_16_3 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__clkbuf_16_3/X
+ pi2_con[1] sky130_fd_sc_hs__clkbuf_16_3/a_114_74# sky130_fd_sc_hs__clkbuf_16
Xsky130_fd_sc_hs__clkbuf_16_107 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__einvp_8_3/TE
+ test_mux_clk_Q_select[0] sky130_fd_sc_hs__clkbuf_16_107/a_114_74# sky130_fd_sc_hs__clkbuf_16
Xsky130_fd_sc_hs__clkbuf_16_118 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__clkbuf_8_69/A
+ sky130_fd_sc_hs__clkbuf_8_97/X sky130_fd_sc_hs__clkbuf_16_119/a_114_74# sky130_fd_sc_hs__clkbuf_16
Xsky130_fd_sc_hs__clkbuf_16_129 DVSS: DVDD: DVDD: DVSS: osc_core_1/pi5_l[3] sky130_fd_sc_hs__clkbuf_4_137/X
+ sky130_fd_sc_hs__clkbuf_16_129/a_114_74# sky130_fd_sc_hs__clkbuf_16
Xsky130_fd_sc_hs__clkbuf_4_107 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__clkbuf_8_35/X
+ osc_core_1/pi2_l[0] sky130_fd_sc_hs__clkbuf_4_107/a_83_270# sky130_fd_sc_hs__clkbuf_4
Xsky130_fd_sc_hs__clkbuf_4_118 DVSS: DVDD: DVDD: DVSS: CTL_BUF_P[1] sky130_fd_sc_hs__clkbuf_4_119/X
+ sky130_fd_sc_hs__clkbuf_4_119/a_83_270# sky130_fd_sc_hs__clkbuf_4
Xsky130_fd_sc_hs__clkbuf_4_129 DVSS: DVDD: DVDD: DVSS: CTL_BUF_N[4] sky130_fd_sc_hs__clkbuf_8_77/A
+ sky130_fd_sc_hs__clkbuf_4_129/a_83_270# sky130_fd_sc_hs__clkbuf_4
Xsky130_fd_sc_hs__o21ai_2_9 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__inv_4_29/A sky130_fd_sc_hs__o21ai_2_9/A2
+ sky130_fd_sc_hs__nand2_2_5/B sky130_fd_sc_hs__buf_2_43/A sky130_fd_sc_hs__o21ai_2_9/a_116_368#
+ sky130_fd_sc_hs__o21ai_2_9/a_27_74# sky130_fd_sc_hs__o21ai_2
Xsky130_fd_sc_hs__clkbuf_4_14 DVSS: DVDD: DVDD: DVSS: manual_control_osc[10] sky130_fd_sc_hs__clkbuf_8_19/A
+ sky130_fd_sc_hs__clkbuf_4_15/a_83_270# sky130_fd_sc_hs__clkbuf_4
Xsky130_fd_sc_hs__clkbuf_4_25 DVSS: DVDD: DVDD: DVSS: manual_control_osc[7] sky130_fd_sc_hs__clkbuf_4_25/X
+ sky130_fd_sc_hs__clkbuf_4_25/a_83_270# sky130_fd_sc_hs__clkbuf_4
Xsky130_fd_sc_hs__clkbuf_8_1 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__clkbuf_8_1/X
+ pi2_con[3] sky130_fd_sc_hs__clkbuf_8_1/a_125_368# sky130_fd_sc_hs__clkbuf_8
Xsky130_fd_sc_hs__clkbuf_4_36 DVSS: DVDD: DVDD: DVSS: ref_clk_ext_p sky130_fd_sc_hs__clkbuf_4_37/X
+ sky130_fd_sc_hs__clkbuf_4_37/a_83_270# sky130_fd_sc_hs__clkbuf_4
Xsky130_fd_sc_hs__clkbuf_4_47 DVSS: DVDD: DVDD: DVSS: manual_control_osc[0] sky130_fd_sc_hs__clkbuf_4_47/X
+ sky130_fd_sc_hs__clkbuf_4_47/a_83_270# sky130_fd_sc_hs__clkbuf_4
Xsky130_fd_sc_hs__clkbuf_4_58 DVSS: DVDD: DVDD: DVSS: fine_con_step_size[1] sky130_fd_sc_hs__clkbuf_4_59/X
+ sky130_fd_sc_hs__clkbuf_4_59/a_83_270# sky130_fd_sc_hs__clkbuf_4
Xsky130_fd_sc_hs__clkbuf_4_69 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__inv_4_9/Y sky130_fd_sc_hs__einvp_2_65/A
+ sky130_fd_sc_hs__clkbuf_4_69/a_83_270# sky130_fd_sc_hs__clkbuf_4
Xsky130_fd_sc_hs__clkinv_8_1 DVSS: DVDD: DVDD: DVSS: prbs_generator_syn_7/out hr_16t4_mux_top_3/din[11]
+ sky130_fd_sc_hs__clkinv_8
Xsky130_fd_sc_hs__clkinv_8_17 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__clkinv_8_19/Y
+ qr_4t1_mux_top_3/rst sky130_fd_sc_hs__clkinv_8
Xsky130_fd_sc_hs__buf_8_3 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__buf_8_3/X sky130_fd_sc_hs__buf_8_3/A
+ sky130_fd_sc_hs__buf_8_3/a_27_74# sky130_fd_sc_hs__buf_8
Xsky130_fd_sc_hs__conb_1_104 DVSS: DVDD: DVDD: DVSS: prbs_generator_syn_13/eqn[30]
+ sky130_fd_sc_hs__conb_1_105/HI sky130_fd_sc_hs__conb_1_105/a_165_290# sky130_fd_sc_hs__conb_1_105/a_21_290#
+ sky130_fd_sc_hs__conb_1
Xsky130_fd_sc_hs__conb_1_115 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__conb_1_115/LO
+ sky130_fd_sc_hs__conb_1_115/HI sky130_fd_sc_hs__conb_1_115/a_165_290# sky130_fd_sc_hs__conb_1_115/a_21_290#
+ sky130_fd_sc_hs__conb_1
Xsky130_fd_sc_hs__conb_1_126 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__conb_1_127/LO
+ sky130_fd_sc_hs__conb_1_127/HI sky130_fd_sc_hs__conb_1_127/a_165_290# sky130_fd_sc_hs__conb_1_127/a_21_290#
+ sky130_fd_sc_hs__conb_1
Xsky130_fd_sc_hs__conb_1_137 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__conb_1_137/LO
+ sky130_fd_sc_hs__conb_1_137/HI sky130_fd_sc_hs__conb_1_137/a_165_290# sky130_fd_sc_hs__conb_1_137/a_21_290#
+ sky130_fd_sc_hs__conb_1
Xsky130_fd_sc_hs__conb_1_148 DVSS: DVDD: DVDD: DVSS: prbs_generator_syn_15/eqn[2]
+ prbs_generator_syn_15/eqn[1] sky130_fd_sc_hs__conb_1_149/a_165_290# sky130_fd_sc_hs__conb_1_149/a_21_290#
+ sky130_fd_sc_hs__conb_1
Xsky130_fd_sc_hs__conb_1_159 DVSS: DVDD: DVDD: DVSS: prbs_generator_syn_17/eqn[31]
+ prbs_generator_syn_17/cke sky130_fd_sc_hs__conb_1_159/a_165_290# sky130_fd_sc_hs__conb_1_159/a_21_290#
+ sky130_fd_sc_hs__conb_1
Xsky130_fd_sc_hs__nand2_8_4 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__nor2_4_3/B sky130_fd_sc_hs__or2b_4_3/A
+ sky130_fd_sc_hs__buf_2_77/A sky130_fd_sc_hs__nand2_8_6/a_27_74# sky130_fd_sc_hs__nand2_8
Xsky130_fd_sc_hs__or4_2_1 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__or4_2_1/X sky130_fd_sc_hs__or4_2_1/D
+ sky130_fd_sc_hs__or4_2_1/A sky130_fd_sc_hs__or4_2_1/B sky130_fd_sc_hs__or4_2_1/C
+ sky130_fd_sc_hs__or4_2_1/a_174_392# sky130_fd_sc_hs__or4_2_1/a_258_392# sky130_fd_sc_hs__or4_2_1/a_342_392#
+ sky130_fd_sc_hs__or4_2_1/a_85_392# sky130_fd_sc_hs__or4_2
Xsky130_fd_sc_hs__einvp_2_104 DVSS: DVDD: DVDD: DVSS: dout_n sky130_fd_sc_hs__einvp_2_9/A
+ sky130_fd_sc_hs__buf_2_93/X sky130_fd_sc_hs__einvp_2_105/a_263_323# sky130_fd_sc_hs__einvp_2_105/a_36_74#
+ sky130_fd_sc_hs__einvp_2_105/a_27_368# sky130_fd_sc_hs__einvp_2
Xsky130_fd_sc_hs__einvp_2_115 DVSS: DVDD: DVDD: DVSS: dout_n sky130_fd_sc_hs__einvp_2_9/A
+ sky130_fd_sc_hs__dlrtp_1_105/Q sky130_fd_sc_hs__einvp_2_115/a_263_323# sky130_fd_sc_hs__einvp_2_115/a_36_74#
+ sky130_fd_sc_hs__einvp_2_115/a_27_368# sky130_fd_sc_hs__einvp_2
Xsky130_fd_sc_hs__einvp_2_126 DVSS: DVDD: DVDD: DVSS: dout_n sky130_fd_sc_hs__buf_8_1/X
+ sky130_fd_sc_hs__dlrtp_1_123/Q sky130_fd_sc_hs__einvp_2_127/a_263_323# sky130_fd_sc_hs__einvp_2_127/a_36_74#
+ sky130_fd_sc_hs__einvp_2_127/a_27_368# sky130_fd_sc_hs__einvp_2
Xsky130_fd_sc_hs__einvp_2_137 DVSS: DVDD: DVDD: DVSS: dout_p sky130_fd_sc_hs__einvp_2_99/A
+ sky130_fd_sc_hs__dlrtp_1_55/Q sky130_fd_sc_hs__einvp_2_137/a_263_323# sky130_fd_sc_hs__einvp_2_137/a_36_74#
+ sky130_fd_sc_hs__einvp_2_137/a_27_368# sky130_fd_sc_hs__einvp_2
Xsky130_fd_sc_hs__einvp_2_148 DVSS: DVDD: DVDD: DVSS: dout_p sky130_fd_sc_hs__einvp_2_99/A
+ sky130_fd_sc_hs__buf_2_159/X sky130_fd_sc_hs__einvp_2_149/a_263_323# sky130_fd_sc_hs__einvp_2_149/a_36_74#
+ sky130_fd_sc_hs__einvp_2_149/a_27_368# sky130_fd_sc_hs__einvp_2
Xsky130_fd_sc_hs__einvp_2_159 DVSS: DVDD: DVDD: DVSS: dout_p sky130_fd_sc_hs__einvp_2_97/A
+ sky130_fd_sc_hs__dlrtp_1_151/Q sky130_fd_sc_hs__einvp_2_159/a_263_323# sky130_fd_sc_hs__einvp_2_159/a_36_74#
+ sky130_fd_sc_hs__einvp_2_159/a_27_368# sky130_fd_sc_hs__einvp_2
Xsky130_fd_sc_hs__clkbuf_16_4 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__clkbuf_8_35/A
+ sky130_fd_sc_hs__clkbuf_4_7/X sky130_fd_sc_hs__clkbuf_16_5/a_114_74# sky130_fd_sc_hs__clkbuf_16
Xsky130_fd_sc_hs__clkbuf_16_108 DVSS: DVDD: DVDD: DVSS: osc_core_1/pi4_l[0] pi4_con[0]
+ sky130_fd_sc_hs__clkbuf_16_109/a_114_74# sky130_fd_sc_hs__clkbuf_16
Xsky130_fd_sc_hs__clkbuf_16_119 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__clkbuf_8_69/A
+ sky130_fd_sc_hs__clkbuf_8_97/X sky130_fd_sc_hs__clkbuf_16_119/a_114_74# sky130_fd_sc_hs__clkbuf_16
Xsky130_fd_sc_hs__clkbuf_4_108 DVSS: DVDD: DVDD: DVSS: fftl_en sky130_fd_sc_hs__clkbuf_4_109/X
+ sky130_fd_sc_hs__clkbuf_4_109/a_83_270# sky130_fd_sc_hs__clkbuf_4
Xsky130_fd_sc_hs__clkbuf_4_119 DVSS: DVDD: DVDD: DVSS: CTL_BUF_P[1] sky130_fd_sc_hs__clkbuf_4_119/X
+ sky130_fd_sc_hs__clkbuf_4_119/a_83_270# sky130_fd_sc_hs__clkbuf_4
Xsky130_fd_sc_hs__clkbuf_8_90 DVSS: DVDD: DVDD: DVSS: prbs_generator_syn_27/inj_err
+ sky130_fd_sc_hs__clkbuf_8_91/A sky130_fd_sc_hs__clkbuf_8_91/a_125_368# sky130_fd_sc_hs__clkbuf_8
Xsky130_fd_sc_hs__clkbuf_4_15 DVSS: DVDD: DVDD: DVSS: manual_control_osc[10] sky130_fd_sc_hs__clkbuf_8_19/A
+ sky130_fd_sc_hs__clkbuf_4_15/a_83_270# sky130_fd_sc_hs__clkbuf_4
Xsky130_fd_sc_hs__clkbuf_4_26 DVSS: DVDD: DVDD: DVSS: manual_control_osc[6] sky130_fd_sc_hs__clkbuf_4_27/X
+ sky130_fd_sc_hs__clkbuf_4_27/a_83_270# sky130_fd_sc_hs__clkbuf_4
Xsky130_fd_sc_hs__clkbuf_4_37 DVSS: DVDD: DVDD: DVSS: ref_clk_ext_p sky130_fd_sc_hs__clkbuf_4_37/X
+ sky130_fd_sc_hs__clkbuf_4_37/a_83_270# sky130_fd_sc_hs__clkbuf_4
Xsky130_fd_sc_hs__clkbuf_8_2 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__clkbuf_8_3/X
+ pi2_con[2] sky130_fd_sc_hs__clkbuf_8_3/a_125_368# sky130_fd_sc_hs__clkbuf_8
Xsky130_fd_sc_hs__clkbuf_4_48 DVSS: DVDD: DVDD: DVSS: prbs_generator_syn_19/inj_err
+ sky130_fd_sc_hs__clkbuf_4_49/X sky130_fd_sc_hs__clkbuf_4_49/a_83_270# sky130_fd_sc_hs__clkbuf_4
Xsky130_fd_sc_hs__clkbuf_4_59 DVSS: DVDD: DVDD: DVSS: fine_con_step_size[1] sky130_fd_sc_hs__clkbuf_4_59/X
+ sky130_fd_sc_hs__clkbuf_4_59/a_83_270# sky130_fd_sc_hs__clkbuf_4
Xsky130_fd_sc_hs__clkinv_8_2 DVSS: DVDD: DVDD: DVSS: prbs_generator_syn_3/out hr_16t4_mux_top_3/din[13]
+ sky130_fd_sc_hs__clkinv_8
Xsky130_fd_sc_hs__clkinv_8_18 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__clkinv_8_19/A
+ sky130_fd_sc_hs__clkinv_8_19/Y sky130_fd_sc_hs__clkinv_8
Xsky130_fd_sc_hs__conb_1_105 DVSS: DVDD: DVDD: DVSS: prbs_generator_syn_13/eqn[30]
+ sky130_fd_sc_hs__conb_1_105/HI sky130_fd_sc_hs__conb_1_105/a_165_290# sky130_fd_sc_hs__conb_1_105/a_21_290#
+ sky130_fd_sc_hs__conb_1
Xsky130_fd_sc_hs__conb_1_116 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__conb_1_117/LO
+ sky130_fd_sc_hs__conb_1_117/HI sky130_fd_sc_hs__conb_1_117/a_165_290# sky130_fd_sc_hs__conb_1_117/a_21_290#
+ sky130_fd_sc_hs__conb_1
Xsky130_fd_sc_hs__conb_1_127 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__conb_1_127/LO
+ sky130_fd_sc_hs__conb_1_127/HI sky130_fd_sc_hs__conb_1_127/a_165_290# sky130_fd_sc_hs__conb_1_127/a_21_290#
+ sky130_fd_sc_hs__conb_1
Xsky130_fd_sc_hs__conb_1_138 DVSS: DVDD: DVDD: DVSS: prbs_generator_syn_15/eqn[22]
+ prbs_generator_syn_15/eqn[20] sky130_fd_sc_hs__conb_1_139/a_165_290# sky130_fd_sc_hs__conb_1_139/a_21_290#
+ sky130_fd_sc_hs__conb_1
Xsky130_fd_sc_hs__conb_1_149 DVSS: DVDD: DVDD: DVSS: prbs_generator_syn_15/eqn[2]
+ prbs_generator_syn_15/eqn[1] sky130_fd_sc_hs__conb_1_149/a_165_290# sky130_fd_sc_hs__conb_1_149/a_21_290#
+ sky130_fd_sc_hs__conb_1
Xsky130_fd_sc_hs__dlrtp_1_150 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__dlrtp_1_151/Q
+ sky130_fd_sc_hs__clkbuf_16_53/X sky130_fd_sc_hs__conb_1_127/HI sky130_fd_sc_hs__o21bai_2_69/Y
+ sky130_fd_sc_hs__dlrtp_1_151/a_216_424# sky130_fd_sc_hs__dlrtp_1_151/a_759_508#
+ sky130_fd_sc_hs__dlrtp_1_151/a_565_74# sky130_fd_sc_hs__dlrtp_1_151/a_27_424# sky130_fd_sc_hs__dlrtp_1_151/a_1045_74#
+ sky130_fd_sc_hs__dlrtp_1_151/a_643_74# sky130_fd_sc_hs__dlrtp_1_151/a_817_48# sky130_fd_sc_hs__dlrtp_1_151/a_568_392#
+ sky130_fd_sc_hs__dlrtp_1_151/a_363_74# sky130_fd_sc_hs__dlrtp_1_151/a_769_74# sky130_fd_sc_hs__dlrtp_1
Xsky130_fd_sc_hs__nand2_8_5 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__nor2_4_3/B sky130_fd_sc_hs__nor2_4_3/A
+ sky130_fd_sc_hs__or2b_2_5/A sky130_fd_sc_hs__nand2_8_7/a_27_74# sky130_fd_sc_hs__nand2_8
Xsky130_fd_sc_hs__clkbuf_2_70 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__buf_4_1/A sky130_fd_sc_hs__buf_1_1/A
+ sky130_fd_sc_hs__clkbuf_2_71/a_43_192# sky130_fd_sc_hs__clkbuf_2
Xsky130_fd_sc_hs__einvp_2_105 DVSS: DVDD: DVDD: DVSS: dout_n sky130_fd_sc_hs__einvp_2_9/A
+ sky130_fd_sc_hs__buf_2_93/X sky130_fd_sc_hs__einvp_2_105/a_263_323# sky130_fd_sc_hs__einvp_2_105/a_36_74#
+ sky130_fd_sc_hs__einvp_2_105/a_27_368# sky130_fd_sc_hs__einvp_2
Xsky130_fd_sc_hs__einvp_2_116 DVSS: DVDD: DVDD: DVSS: dout_n sky130_fd_sc_hs__einvp_2_9/A
+ sky130_fd_sc_hs__buf_2_115/X sky130_fd_sc_hs__einvp_2_117/a_263_323# sky130_fd_sc_hs__einvp_2_117/a_36_74#
+ sky130_fd_sc_hs__einvp_2_117/a_27_368# sky130_fd_sc_hs__einvp_2
Xsky130_fd_sc_hs__einvp_2_127 DVSS: DVDD: DVDD: DVSS: dout_n sky130_fd_sc_hs__buf_8_1/X
+ sky130_fd_sc_hs__dlrtp_1_123/Q sky130_fd_sc_hs__einvp_2_127/a_263_323# sky130_fd_sc_hs__einvp_2_127/a_36_74#
+ sky130_fd_sc_hs__einvp_2_127/a_27_368# sky130_fd_sc_hs__einvp_2
Xsky130_fd_sc_hs__einvp_2_138 DVSS: DVDD: DVDD: DVSS: dout_p sky130_fd_sc_hs__einvp_2_99/A
+ sky130_fd_sc_hs__dlrtp_1_137/Q sky130_fd_sc_hs__einvp_2_139/a_263_323# sky130_fd_sc_hs__einvp_2_139/a_36_74#
+ sky130_fd_sc_hs__einvp_2_139/a_27_368# sky130_fd_sc_hs__einvp_2
Xsky130_fd_sc_hs__einvp_2_149 DVSS: DVDD: DVDD: DVSS: dout_p sky130_fd_sc_hs__einvp_2_99/A
+ sky130_fd_sc_hs__buf_2_159/X sky130_fd_sc_hs__einvp_2_149/a_263_323# sky130_fd_sc_hs__einvp_2_149/a_36_74#
+ sky130_fd_sc_hs__einvp_2_149/a_27_368# sky130_fd_sc_hs__einvp_2
Xsky130_fd_sc_hs__clkbuf_16_5 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__clkbuf_8_35/A
+ sky130_fd_sc_hs__clkbuf_4_7/X sky130_fd_sc_hs__clkbuf_16_5/a_114_74# sky130_fd_sc_hs__clkbuf_16
Xsky130_fd_sc_hs__clkbuf_16_109 DVSS: DVDD: DVDD: DVSS: osc_core_1/pi4_l[0] pi4_con[0]
+ sky130_fd_sc_hs__clkbuf_16_109/a_114_74# sky130_fd_sc_hs__clkbuf_16
Xsky130_fd_sc_hs__clkbuf_4_109 DVSS: DVDD: DVDD: DVSS: fftl_en sky130_fd_sc_hs__clkbuf_4_109/X
+ sky130_fd_sc_hs__clkbuf_4_109/a_83_270# sky130_fd_sc_hs__clkbuf_4
Xsky130_fd_sc_hs__clkbuf_8_80 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__clkbuf_8_81/X
+ CTL_BUF_P[2] sky130_fd_sc_hs__clkbuf_8_81/a_125_368# sky130_fd_sc_hs__clkbuf_8
Xsky130_fd_sc_hs__clkbuf_8_91 DVSS: DVDD: DVDD: DVSS: prbs_generator_syn_27/inj_err
+ sky130_fd_sc_hs__clkbuf_8_91/A sky130_fd_sc_hs__clkbuf_8_91/a_125_368# sky130_fd_sc_hs__clkbuf_8
Xsky130_fd_sc_hs__clkbuf_4_16 DVSS: DVDD: DVDD: DVSS: manual_control_osc[9] sky130_fd_sc_hs__clkbuf_8_13/A
+ sky130_fd_sc_hs__clkbuf_4_17/a_83_270# sky130_fd_sc_hs__clkbuf_4
Xsky130_fd_sc_hs__einvp_8_0 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__einvp_8_3/Z sky130_fd_sc_hs__einvp_8_1/TE
+ osc_core_1/p1 sky130_fd_sc_hs__einvp_8_1/a_802_323# sky130_fd_sc_hs__einvp_8_1/a_27_74#
+ sky130_fd_sc_hs__einvp_8_1/a_27_368# sky130_fd_sc_hs__einvp_8
Xsky130_fd_sc_hs__clkbuf_4_27 DVSS: DVDD: DVDD: DVSS: manual_control_osc[6] sky130_fd_sc_hs__clkbuf_4_27/X
+ sky130_fd_sc_hs__clkbuf_4_27/a_83_270# sky130_fd_sc_hs__clkbuf_4
Xsky130_fd_sc_hs__clkbuf_4_38 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__clkbuf_4_49/X
+ sky130_fd_sc_hs__clkbuf_4_39/X sky130_fd_sc_hs__clkbuf_4_39/a_83_270# sky130_fd_sc_hs__clkbuf_4
Xsky130_fd_sc_hs__clkbuf_8_3 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__clkbuf_8_3/X
+ pi2_con[2] sky130_fd_sc_hs__clkbuf_8_3/a_125_368# sky130_fd_sc_hs__clkbuf_8
Xsky130_fd_sc_hs__clkbuf_4_49 DVSS: DVDD: DVDD: DVSS: prbs_generator_syn_19/inj_err
+ sky130_fd_sc_hs__clkbuf_4_49/X sky130_fd_sc_hs__clkbuf_4_49/a_83_270# sky130_fd_sc_hs__clkbuf_4
Xsky130_fd_sc_hs__clkinv_8_3 DVSS: DVDD: DVDD: DVSS: prbs_generator_syn_3/out hr_16t4_mux_top_3/din[13]
+ sky130_fd_sc_hs__clkinv_8
Xsky130_fd_sc_hs__clkinv_8_19 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__clkinv_8_19/A
+ sky130_fd_sc_hs__clkinv_8_19/Y sky130_fd_sc_hs__clkinv_8
Xsky130_fd_sc_hs__conb_1_106 DVSS: DVDD: DVDD: DVSS: prbs_generator_syn_13/eqn[31]
+ prbs_generator_syn_13/cke sky130_fd_sc_hs__conb_1_107/a_165_290# sky130_fd_sc_hs__conb_1_107/a_21_290#
+ sky130_fd_sc_hs__conb_1
Xsky130_fd_sc_hs__conb_1_117 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__conb_1_117/LO
+ sky130_fd_sc_hs__conb_1_117/HI sky130_fd_sc_hs__conb_1_117/a_165_290# sky130_fd_sc_hs__conb_1_117/a_21_290#
+ sky130_fd_sc_hs__conb_1
Xsky130_fd_sc_hs__conb_1_128 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__conb_1_129/LO
+ sky130_fd_sc_hs__conb_1_129/HI sky130_fd_sc_hs__conb_1_129/a_165_290# sky130_fd_sc_hs__conb_1_129/a_21_290#
+ sky130_fd_sc_hs__conb_1
Xsky130_fd_sc_hs__conb_1_139 DVSS: DVDD: DVDD: DVSS: prbs_generator_syn_15/eqn[22]
+ prbs_generator_syn_15/eqn[20] sky130_fd_sc_hs__conb_1_139/a_165_290# sky130_fd_sc_hs__conb_1_139/a_21_290#
+ sky130_fd_sc_hs__conb_1
Xsky130_fd_sc_hs__dlrtp_1_140 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__einvp_2_75/TE
+ sky130_fd_sc_hs__clkbuf_16_53/X sky130_fd_sc_hs__conb_1_127/HI sky130_fd_sc_hs__buf_2_143/X
+ sky130_fd_sc_hs__dlrtp_1_141/a_216_424# sky130_fd_sc_hs__dlrtp_1_141/a_759_508#
+ sky130_fd_sc_hs__dlrtp_1_141/a_565_74# sky130_fd_sc_hs__dlrtp_1_141/a_27_424# sky130_fd_sc_hs__dlrtp_1_141/a_1045_74#
+ sky130_fd_sc_hs__dlrtp_1_141/a_643_74# sky130_fd_sc_hs__dlrtp_1_141/a_817_48# sky130_fd_sc_hs__dlrtp_1_141/a_568_392#
+ sky130_fd_sc_hs__dlrtp_1_141/a_363_74# sky130_fd_sc_hs__dlrtp_1_141/a_769_74# sky130_fd_sc_hs__dlrtp_1
Xsky130_fd_sc_hs__dlrtp_1_151 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__dlrtp_1_151/Q
+ sky130_fd_sc_hs__clkbuf_16_53/X sky130_fd_sc_hs__conb_1_127/HI sky130_fd_sc_hs__o21bai_2_69/Y
+ sky130_fd_sc_hs__dlrtp_1_151/a_216_424# sky130_fd_sc_hs__dlrtp_1_151/a_759_508#
+ sky130_fd_sc_hs__dlrtp_1_151/a_565_74# sky130_fd_sc_hs__dlrtp_1_151/a_27_424# sky130_fd_sc_hs__dlrtp_1_151/a_1045_74#
+ sky130_fd_sc_hs__dlrtp_1_151/a_643_74# sky130_fd_sc_hs__dlrtp_1_151/a_817_48# sky130_fd_sc_hs__dlrtp_1_151/a_568_392#
+ sky130_fd_sc_hs__dlrtp_1_151/a_363_74# sky130_fd_sc_hs__dlrtp_1_151/a_769_74# sky130_fd_sc_hs__dlrtp_1
Xsky130_fd_sc_hs__nand2_8_6 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__nor2_4_3/B sky130_fd_sc_hs__or2b_4_3/A
+ sky130_fd_sc_hs__buf_2_77/A sky130_fd_sc_hs__nand2_8_6/a_27_74# sky130_fd_sc_hs__nand2_8
Xsky130_fd_sc_hs__clkbuf_2_60 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__dlrtp_1_133/D
+ sky130_fd_sc_hs__o21ai_2_51/Y sky130_fd_sc_hs__clkbuf_2_61/a_43_192# sky130_fd_sc_hs__clkbuf_2
Xsky130_fd_sc_hs__clkbuf_2_71 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__buf_4_1/A sky130_fd_sc_hs__buf_1_1/A
+ sky130_fd_sc_hs__clkbuf_2_71/a_43_192# sky130_fd_sc_hs__clkbuf_2
Xsky130_fd_sc_hs__einvp_2_106 DVSS: DVDD: DVDD: DVSS: dout_n sky130_fd_sc_hs__einvp_2_9/A
+ sky130_fd_sc_hs__dlrtp_1_98/Q sky130_fd_sc_hs__einvp_2_107/a_263_323# sky130_fd_sc_hs__einvp_2_107/a_36_74#
+ sky130_fd_sc_hs__einvp_2_107/a_27_368# sky130_fd_sc_hs__einvp_2
Xsky130_fd_sc_hs__einvp_2_117 DVSS: DVDD: DVDD: DVSS: dout_n sky130_fd_sc_hs__einvp_2_9/A
+ sky130_fd_sc_hs__buf_2_115/X sky130_fd_sc_hs__einvp_2_117/a_263_323# sky130_fd_sc_hs__einvp_2_117/a_36_74#
+ sky130_fd_sc_hs__einvp_2_117/a_27_368# sky130_fd_sc_hs__einvp_2
Xsky130_fd_sc_hs__einvp_2_128 DVSS: DVDD: DVDD: DVSS: dout_n sky130_fd_sc_hs__buf_8_1/X
+ sky130_fd_sc_hs__dlrtp_1_133/Q sky130_fd_sc_hs__einvp_2_129/a_263_323# sky130_fd_sc_hs__einvp_2_129/a_36_74#
+ sky130_fd_sc_hs__einvp_2_129/a_27_368# sky130_fd_sc_hs__einvp_2
Xsky130_fd_sc_hs__einvp_2_139 DVSS: DVDD: DVDD: DVSS: dout_p sky130_fd_sc_hs__einvp_2_99/A
+ sky130_fd_sc_hs__dlrtp_1_137/Q sky130_fd_sc_hs__einvp_2_139/a_263_323# sky130_fd_sc_hs__einvp_2_139/a_36_74#
+ sky130_fd_sc_hs__einvp_2_139/a_27_368# sky130_fd_sc_hs__einvp_2
Xsky130_fd_sc_hs__clkbuf_16_6 DVSS: DVDD: DVDD: DVSS: prbs_generator_syn_9/rst prbs_generator_syn_13/rst
+ sky130_fd_sc_hs__clkbuf_16_7/a_114_74# sky130_fd_sc_hs__clkbuf_16
Xsky130_fd_sc_hs__clkbuf_8_70 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__or2b_4_3/A
+ sky130_fd_sc_hs__clkbuf_8_71/A sky130_fd_sc_hs__clkbuf_8_71/a_125_368# sky130_fd_sc_hs__clkbuf_8
Xsky130_fd_sc_hs__clkbuf_8_81 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__clkbuf_8_81/X
+ CTL_BUF_P[2] sky130_fd_sc_hs__clkbuf_8_81/a_125_368# sky130_fd_sc_hs__clkbuf_8
Xsky130_fd_sc_hs__clkbuf_8_92 DVSS: DVDD: DVDD: DVSS: prbs_generator_syn_27/rst sky130_fd_sc_hs__clkbuf_8_93/A
+ sky130_fd_sc_hs__clkbuf_8_93/a_125_368# sky130_fd_sc_hs__clkbuf_8
Xsky130_fd_sc_hs__clkbuf_4_17 DVSS: DVDD: DVDD: DVSS: manual_control_osc[9] sky130_fd_sc_hs__clkbuf_8_13/A
+ sky130_fd_sc_hs__clkbuf_4_17/a_83_270# sky130_fd_sc_hs__clkbuf_4
Xsky130_fd_sc_hs__einvp_8_1 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__einvp_8_3/Z sky130_fd_sc_hs__einvp_8_1/TE
+ osc_core_1/p1 sky130_fd_sc_hs__einvp_8_1/a_802_323# sky130_fd_sc_hs__einvp_8_1/a_27_74#
+ sky130_fd_sc_hs__einvp_8_1/a_27_368# sky130_fd_sc_hs__einvp_8
Xsky130_fd_sc_hs__clkbuf_4_28 DVSS: DVDD: DVDD: DVSS: manual_control_osc[2] sky130_fd_sc_hs__clkbuf_4_51/A
+ sky130_fd_sc_hs__clkbuf_4_29/a_83_270# sky130_fd_sc_hs__clkbuf_4
Xsky130_fd_sc_hs__clkbuf_4_39 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__clkbuf_4_49/X
+ sky130_fd_sc_hs__clkbuf_4_39/X sky130_fd_sc_hs__clkbuf_4_39/a_83_270# sky130_fd_sc_hs__clkbuf_4
Xsky130_fd_sc_hs__clkbuf_8_4 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__clkbuf_8_5/X
+ sky130_fd_sc_hs__clkbuf_8_5/A sky130_fd_sc_hs__clkbuf_8_5/a_125_368# sky130_fd_sc_hs__clkbuf_8
Xsky130_fd_sc_hs__clkinv_8_4 DVSS: DVDD: DVDD: DVSS: prbs_generator_syn_11/out hr_16t4_mux_top_3/din[15]
+ sky130_fd_sc_hs__clkinv_8
Xsky130_fd_sc_hs__conb_1_107 DVSS: DVDD: DVDD: DVSS: prbs_generator_syn_13/eqn[31]
+ prbs_generator_syn_13/cke sky130_fd_sc_hs__conb_1_107/a_165_290# sky130_fd_sc_hs__conb_1_107/a_21_290#
+ sky130_fd_sc_hs__conb_1
Xsky130_fd_sc_hs__conb_1_118 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__conb_1_119/LO
+ sky130_fd_sc_hs__conb_1_119/HI sky130_fd_sc_hs__conb_1_119/a_165_290# sky130_fd_sc_hs__conb_1_119/a_21_290#
+ sky130_fd_sc_hs__conb_1
Xsky130_fd_sc_hs__conb_1_129 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__conb_1_129/LO
+ sky130_fd_sc_hs__conb_1_129/HI sky130_fd_sc_hs__conb_1_129/a_165_290# sky130_fd_sc_hs__conb_1_129/a_21_290#
+ sky130_fd_sc_hs__conb_1
Xsky130_fd_sc_hs__buf_4_0 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__buf_4_1/A hr_16t4_mux_top_3/clk
+ sky130_fd_sc_hs__buf_4_1/a_86_260# sky130_fd_sc_hs__buf_4
Xsky130_fd_sc_hs__dlrtp_1_130 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__dlrtp_1_131/Q
+ sky130_fd_sc_hs__clkbuf_16_53/X sky130_fd_sc_hs__conb_1_135/HI sky130_fd_sc_hs__clkbuf_2_7/X
+ sky130_fd_sc_hs__dlrtp_1_131/a_216_424# sky130_fd_sc_hs__dlrtp_1_131/a_759_508#
+ sky130_fd_sc_hs__dlrtp_1_131/a_565_74# sky130_fd_sc_hs__dlrtp_1_131/a_27_424# sky130_fd_sc_hs__dlrtp_1_131/a_1045_74#
+ sky130_fd_sc_hs__dlrtp_1_131/a_643_74# sky130_fd_sc_hs__dlrtp_1_131/a_817_48# sky130_fd_sc_hs__dlrtp_1_131/a_568_392#
+ sky130_fd_sc_hs__dlrtp_1_131/a_363_74# sky130_fd_sc_hs__dlrtp_1_131/a_769_74# sky130_fd_sc_hs__dlrtp_1
Xsky130_fd_sc_hs__dlrtp_1_141 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__einvp_2_75/TE
+ sky130_fd_sc_hs__clkbuf_16_53/X sky130_fd_sc_hs__conb_1_127/HI sky130_fd_sc_hs__buf_2_143/X
+ sky130_fd_sc_hs__dlrtp_1_141/a_216_424# sky130_fd_sc_hs__dlrtp_1_141/a_759_508#
+ sky130_fd_sc_hs__dlrtp_1_141/a_565_74# sky130_fd_sc_hs__dlrtp_1_141/a_27_424# sky130_fd_sc_hs__dlrtp_1_141/a_1045_74#
+ sky130_fd_sc_hs__dlrtp_1_141/a_643_74# sky130_fd_sc_hs__dlrtp_1_141/a_817_48# sky130_fd_sc_hs__dlrtp_1_141/a_568_392#
+ sky130_fd_sc_hs__dlrtp_1_141/a_363_74# sky130_fd_sc_hs__dlrtp_1_141/a_769_74# sky130_fd_sc_hs__dlrtp_1
Xsky130_fd_sc_hs__dlrtp_1_152 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__dlrtp_1_153/Q
+ sky130_fd_sc_hs__clkbuf_16_53/X sky130_fd_sc_hs__conb_1_127/HI sky130_fd_sc_hs__dlrtp_1_153/D
+ sky130_fd_sc_hs__dlrtp_1_153/a_216_424# sky130_fd_sc_hs__dlrtp_1_153/a_759_508#
+ sky130_fd_sc_hs__dlrtp_1_153/a_565_74# sky130_fd_sc_hs__dlrtp_1_153/a_27_424# sky130_fd_sc_hs__dlrtp_1_153/a_1045_74#
+ sky130_fd_sc_hs__dlrtp_1_153/a_643_74# sky130_fd_sc_hs__dlrtp_1_153/a_817_48# sky130_fd_sc_hs__dlrtp_1_153/a_568_392#
+ sky130_fd_sc_hs__dlrtp_1_153/a_363_74# sky130_fd_sc_hs__dlrtp_1_153/a_769_74# sky130_fd_sc_hs__dlrtp_1
Xsky130_fd_sc_hs__nand2_8_7 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__nor2_4_3/B sky130_fd_sc_hs__nor2_4_3/A
+ sky130_fd_sc_hs__or2b_2_5/A sky130_fd_sc_hs__nand2_8_7/a_27_74# sky130_fd_sc_hs__nand2_8
Xsky130_fd_sc_hs__inv_4_0 DVSS: DVDD: DVDD: DVSS: test_mux_clk_Q sky130_fd_sc_hs__inv_4_1/A
+ sky130_fd_sc_hs__inv_4
Xsky130_fd_sc_hs__clkbuf_2_50 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__dlrtp_1_115/D
+ sky130_fd_sc_hs__o21ai_2_41/Y sky130_fd_sc_hs__clkbuf_2_51/a_43_192# sky130_fd_sc_hs__clkbuf_2
Xsky130_fd_sc_hs__clkbuf_2_61 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__dlrtp_1_133/D
+ sky130_fd_sc_hs__o21ai_2_51/Y sky130_fd_sc_hs__clkbuf_2_61/a_43_192# sky130_fd_sc_hs__clkbuf_2
Xsky130_fd_sc_hs__einvp_2_107 DVSS: DVDD: DVDD: DVSS: dout_n sky130_fd_sc_hs__einvp_2_9/A
+ sky130_fd_sc_hs__dlrtp_1_98/Q sky130_fd_sc_hs__einvp_2_107/a_263_323# sky130_fd_sc_hs__einvp_2_107/a_36_74#
+ sky130_fd_sc_hs__einvp_2_107/a_27_368# sky130_fd_sc_hs__einvp_2
Xsky130_fd_sc_hs__einvp_2_118 DVSS: DVDD: DVDD: DVSS: dout_n sky130_fd_sc_hs__einvp_2_9/A
+ sky130_fd_sc_hs__dlrtp_1_111/Q sky130_fd_sc_hs__einvp_2_119/a_263_323# sky130_fd_sc_hs__einvp_2_119/a_36_74#
+ sky130_fd_sc_hs__einvp_2_119/a_27_368# sky130_fd_sc_hs__einvp_2
Xsky130_fd_sc_hs__einvp_2_129 DVSS: DVDD: DVDD: DVSS: dout_n sky130_fd_sc_hs__buf_8_1/X
+ sky130_fd_sc_hs__dlrtp_1_133/Q sky130_fd_sc_hs__einvp_2_129/a_263_323# sky130_fd_sc_hs__einvp_2_129/a_36_74#
+ sky130_fd_sc_hs__einvp_2_129/a_27_368# sky130_fd_sc_hs__einvp_2
Xsky130_fd_sc_hs__clkbuf_16_7 DVSS: DVDD: DVDD: DVSS: prbs_generator_syn_9/rst prbs_generator_syn_13/rst
+ sky130_fd_sc_hs__clkbuf_16_7/a_114_74# sky130_fd_sc_hs__clkbuf_16
Xsky130_fd_sc_hs__buf_2_90 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__buf_2_91/A sky130_fd_sc_hs__buf_2_91/X
+ sky130_fd_sc_hs__buf_2_91/a_21_260# sky130_fd_sc_hs__buf_2
Xsky130_fd_sc_hs__o21bai_2_70 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__buf_2_77/A
+ sky130_fd_sc_hs__o21bai_4_7/A1 sky130_fd_sc_hs__dlrtp_1_157/D sky130_fd_sc_hs__buf_2_75/A
+ sky130_fd_sc_hs__o21bai_2_71/a_27_74# sky130_fd_sc_hs__o21bai_2_71/a_225_74# sky130_fd_sc_hs__o21bai_2_71/a_507_368#
+ sky130_fd_sc_hs__o21bai_2
Xsky130_fd_sc_hs__clkbuf_8_60 DVSS: DVDD: DVDD: DVSS: osc_core_1/con_perb_5[3] con_perb[3]
+ sky130_fd_sc_hs__clkbuf_8_61/a_125_368# sky130_fd_sc_hs__clkbuf_8
Xsky130_fd_sc_hs__clkbuf_8_71 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__or2b_4_3/A
+ sky130_fd_sc_hs__clkbuf_8_71/A sky130_fd_sc_hs__clkbuf_8_71/a_125_368# sky130_fd_sc_hs__clkbuf_8
Xsky130_fd_sc_hs__clkbuf_8_82 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__einvp_8_9/TE
+ test_mux_select[0] sky130_fd_sc_hs__clkbuf_8_83/a_125_368# sky130_fd_sc_hs__clkbuf_8
Xsky130_fd_sc_hs__clkbuf_8_93 DVSS: DVDD: DVDD: DVSS: prbs_generator_syn_27/rst sky130_fd_sc_hs__clkbuf_8_93/A
+ sky130_fd_sc_hs__clkbuf_8_93/a_125_368# sky130_fd_sc_hs__clkbuf_8
Xsky130_fd_sc_hs__clkbuf_4_18 DVSS: DVDD: DVDD: DVSS: pi1_con[1] sky130_fd_sc_hs__clkbuf_4_19/X
+ sky130_fd_sc_hs__clkbuf_4_19/a_83_270# sky130_fd_sc_hs__clkbuf_4
Xsky130_fd_sc_hs__einvp_8_2 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__einvp_8_3/Z sky130_fd_sc_hs__einvp_8_3/TE
+ osc_core_1/p5 sky130_fd_sc_hs__einvp_8_3/a_802_323# sky130_fd_sc_hs__einvp_8_3/a_27_74#
+ sky130_fd_sc_hs__einvp_8_3/a_27_368# sky130_fd_sc_hs__einvp_8
Xsky130_fd_sc_hs__clkbuf_4_29 DVSS: DVDD: DVDD: DVSS: manual_control_osc[2] sky130_fd_sc_hs__clkbuf_4_51/A
+ sky130_fd_sc_hs__clkbuf_4_29/a_83_270# sky130_fd_sc_hs__clkbuf_4
Xsky130_fd_sc_hs__clkbuf_8_5 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__clkbuf_8_5/X
+ sky130_fd_sc_hs__clkbuf_8_5/A sky130_fd_sc_hs__clkbuf_8_5/a_125_368# sky130_fd_sc_hs__clkbuf_8
Xsky130_fd_sc_hs__clkinv_8_5 DVSS: DVDD: DVDD: DVSS: prbs_generator_syn_11/out hr_16t4_mux_top_3/din[15]
+ sky130_fd_sc_hs__clkinv_8
Xsky130_fd_sc_hs__conb_1_108 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__conb_1_109/LO
+ sky130_fd_sc_hs__conb_1_109/HI sky130_fd_sc_hs__conb_1_109/a_165_290# sky130_fd_sc_hs__conb_1_109/a_21_290#
+ sky130_fd_sc_hs__conb_1
Xsky130_fd_sc_hs__conb_1_119 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__conb_1_119/LO
+ sky130_fd_sc_hs__conb_1_119/HI sky130_fd_sc_hs__conb_1_119/a_165_290# sky130_fd_sc_hs__conb_1_119/a_21_290#
+ sky130_fd_sc_hs__conb_1
Xsky130_fd_sc_hs__buf_4_1 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__buf_4_1/A hr_16t4_mux_top_3/clk
+ sky130_fd_sc_hs__buf_4_1/a_86_260# sky130_fd_sc_hs__buf_4
Xsky130_fd_sc_hs__dlrtp_1_120 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__dlrtp_1_121/Q
+ sky130_fd_sc_hs__dlrtp_1_9/GATE sky130_fd_sc_hs__conb_1_131/HI sky130_fd_sc_hs__dlrtp_1_121/D
+ sky130_fd_sc_hs__dlrtp_1_121/a_216_424# sky130_fd_sc_hs__dlrtp_1_121/a_759_508#
+ sky130_fd_sc_hs__dlrtp_1_121/a_565_74# sky130_fd_sc_hs__dlrtp_1_121/a_27_424# sky130_fd_sc_hs__dlrtp_1_121/a_1045_74#
+ sky130_fd_sc_hs__dlrtp_1_121/a_643_74# sky130_fd_sc_hs__dlrtp_1_121/a_817_48# sky130_fd_sc_hs__dlrtp_1_121/a_568_392#
+ sky130_fd_sc_hs__dlrtp_1_121/a_363_74# sky130_fd_sc_hs__dlrtp_1_121/a_769_74# sky130_fd_sc_hs__dlrtp_1
Xsky130_fd_sc_hs__dlrtp_1_131 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__dlrtp_1_131/Q
+ sky130_fd_sc_hs__clkbuf_16_53/X sky130_fd_sc_hs__conb_1_135/HI sky130_fd_sc_hs__clkbuf_2_7/X
+ sky130_fd_sc_hs__dlrtp_1_131/a_216_424# sky130_fd_sc_hs__dlrtp_1_131/a_759_508#
+ sky130_fd_sc_hs__dlrtp_1_131/a_565_74# sky130_fd_sc_hs__dlrtp_1_131/a_27_424# sky130_fd_sc_hs__dlrtp_1_131/a_1045_74#
+ sky130_fd_sc_hs__dlrtp_1_131/a_643_74# sky130_fd_sc_hs__dlrtp_1_131/a_817_48# sky130_fd_sc_hs__dlrtp_1_131/a_568_392#
+ sky130_fd_sc_hs__dlrtp_1_131/a_363_74# sky130_fd_sc_hs__dlrtp_1_131/a_769_74# sky130_fd_sc_hs__dlrtp_1
Xsky130_fd_sc_hs__dlrtp_1_142 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__dlrtp_1_143/Q
+ sky130_fd_sc_hs__clkbuf_16_53/X sky130_fd_sc_hs__conb_1_127/HI sky130_fd_sc_hs__dlrtp_1_143/D
+ sky130_fd_sc_hs__dlrtp_1_143/a_216_424# sky130_fd_sc_hs__dlrtp_1_143/a_759_508#
+ sky130_fd_sc_hs__dlrtp_1_143/a_565_74# sky130_fd_sc_hs__dlrtp_1_143/a_27_424# sky130_fd_sc_hs__dlrtp_1_143/a_1045_74#
+ sky130_fd_sc_hs__dlrtp_1_143/a_643_74# sky130_fd_sc_hs__dlrtp_1_143/a_817_48# sky130_fd_sc_hs__dlrtp_1_143/a_568_392#
+ sky130_fd_sc_hs__dlrtp_1_143/a_363_74# sky130_fd_sc_hs__dlrtp_1_143/a_769_74# sky130_fd_sc_hs__dlrtp_1
Xsky130_fd_sc_hs__dlrtp_1_153 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__dlrtp_1_153/Q
+ sky130_fd_sc_hs__clkbuf_16_53/X sky130_fd_sc_hs__conb_1_127/HI sky130_fd_sc_hs__dlrtp_1_153/D
+ sky130_fd_sc_hs__dlrtp_1_153/a_216_424# sky130_fd_sc_hs__dlrtp_1_153/a_759_508#
+ sky130_fd_sc_hs__dlrtp_1_153/a_565_74# sky130_fd_sc_hs__dlrtp_1_153/a_27_424# sky130_fd_sc_hs__dlrtp_1_153/a_1045_74#
+ sky130_fd_sc_hs__dlrtp_1_153/a_643_74# sky130_fd_sc_hs__dlrtp_1_153/a_817_48# sky130_fd_sc_hs__dlrtp_1_153/a_568_392#
+ sky130_fd_sc_hs__dlrtp_1_153/a_363_74# sky130_fd_sc_hs__dlrtp_1_153/a_769_74# sky130_fd_sc_hs__dlrtp_1
Xsky130_fd_sc_hs__inv_4_1 DVSS: DVDD: DVDD: DVSS: test_mux_clk_Q sky130_fd_sc_hs__inv_4_1/A
+ sky130_fd_sc_hs__inv_4
Xsky130_fd_sc_hs__clkbuf_2_40 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__dlrtp_1_107/D
+ sky130_fd_sc_hs__buf_2_113/X sky130_fd_sc_hs__clkbuf_2_41/a_43_192# sky130_fd_sc_hs__clkbuf_2
Xsky130_fd_sc_hs__clkbuf_2_51 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__dlrtp_1_115/D
+ sky130_fd_sc_hs__o21ai_2_41/Y sky130_fd_sc_hs__clkbuf_2_51/a_43_192# sky130_fd_sc_hs__clkbuf_2
Xsky130_fd_sc_hs__clkbuf_2_62 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__einvp_8_1/TE
+ sky130_fd_sc_hs__einvp_8_3/TE sky130_fd_sc_hs__clkbuf_2_63/a_43_192# sky130_fd_sc_hs__clkbuf_2
Xsky130_fd_sc_hs__einvp_2_108 DVSS: DVDD: DVDD: DVSS: dout_n sky130_fd_sc_hs__einvp_2_9/A
+ sky130_fd_sc_hs__dlrtp_1_95/Q sky130_fd_sc_hs__einvp_2_109/a_263_323# sky130_fd_sc_hs__einvp_2_109/a_36_74#
+ sky130_fd_sc_hs__einvp_2_109/a_27_368# sky130_fd_sc_hs__einvp_2
Xsky130_fd_sc_hs__einvp_2_119 DVSS: DVDD: DVDD: DVSS: dout_n sky130_fd_sc_hs__einvp_2_9/A
+ sky130_fd_sc_hs__dlrtp_1_111/Q sky130_fd_sc_hs__einvp_2_119/a_263_323# sky130_fd_sc_hs__einvp_2_119/a_36_74#
+ sky130_fd_sc_hs__einvp_2_119/a_27_368# sky130_fd_sc_hs__einvp_2
Xsky130_fd_sc_hs__clkbuf_16_8 DVSS: DVDD: DVDD: DVSS: prbs_generator_syn_9/inj_err
+ sky130_fd_sc_hs__clkbuf_4_39/X sky130_fd_sc_hs__clkbuf_16_9/a_114_74# sky130_fd_sc_hs__clkbuf_16
Xsky130_fd_sc_hs__dlrtp_1_0 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__dlrtp_1_1/Q sky130_fd_sc_hs__dlrtp_1_9/GATE
+ sky130_fd_sc_hs__conb_1_117/HI sky130_fd_sc_hs__buf_2_81/X sky130_fd_sc_hs__dlrtp_1_1/a_216_424#
+ sky130_fd_sc_hs__dlrtp_1_1/a_759_508# sky130_fd_sc_hs__dlrtp_1_1/a_565_74# sky130_fd_sc_hs__dlrtp_1_1/a_27_424#
+ sky130_fd_sc_hs__dlrtp_1_1/a_1045_74# sky130_fd_sc_hs__dlrtp_1_1/a_643_74# sky130_fd_sc_hs__dlrtp_1_1/a_817_48#
+ sky130_fd_sc_hs__dlrtp_1_1/a_568_392# sky130_fd_sc_hs__dlrtp_1_1/a_363_74# sky130_fd_sc_hs__dlrtp_1_1/a_769_74#
+ sky130_fd_sc_hs__dlrtp_1
Xsky130_fd_sc_hs__buf_2_80 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__buf_2_83/X sky130_fd_sc_hs__buf_2_81/X
+ sky130_fd_sc_hs__buf_2_81/a_21_260# sky130_fd_sc_hs__buf_2
Xsky130_fd_sc_hs__buf_2_91 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__buf_2_91/A sky130_fd_sc_hs__buf_2_91/X
+ sky130_fd_sc_hs__buf_2_91/a_21_260# sky130_fd_sc_hs__buf_2
Xsky130_fd_sc_hs__o21bai_2_60 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__inv_8_1/Y sky130_fd_sc_hs__nand2_2_5/B
+ sky130_fd_sc_hs__dlrtp_1_143/D sky130_fd_sc_hs__o21bai_2_61/Y sky130_fd_sc_hs__o21bai_2_61/a_27_74#
+ sky130_fd_sc_hs__o21bai_2_61/a_225_74# sky130_fd_sc_hs__o21bai_2_61/a_507_368# sky130_fd_sc_hs__o21bai_2
Xsky130_fd_sc_hs__o21bai_2_71 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__buf_2_77/A
+ sky130_fd_sc_hs__o21bai_4_7/A1 sky130_fd_sc_hs__dlrtp_1_157/D sky130_fd_sc_hs__buf_2_75/A
+ sky130_fd_sc_hs__o21bai_2_71/a_27_74# sky130_fd_sc_hs__o21bai_2_71/a_225_74# sky130_fd_sc_hs__o21bai_2_71/a_507_368#
+ sky130_fd_sc_hs__o21bai_2
Xsky130_fd_sc_hs__clkbuf_8_50 DVSS: DVDD: DVDD: DVSS: qr_4t1_mux_top_3/clk_Q sky130_fd_sc_hs__einvn_8_1/Z
+ sky130_fd_sc_hs__clkbuf_8_51/a_125_368# sky130_fd_sc_hs__clkbuf_8
Xsky130_fd_sc_hs__clkbuf_8_61 DVSS: DVDD: DVDD: DVSS: osc_core_1/con_perb_5[3] con_perb[3]
+ sky130_fd_sc_hs__clkbuf_8_61/a_125_368# sky130_fd_sc_hs__clkbuf_8
Xsky130_fd_sc_hs__clkbuf_8_72 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__nor2_4_3/A
+ sky130_fd_sc_hs__clkbuf_8_77/X sky130_fd_sc_hs__clkbuf_8_73/a_125_368# sky130_fd_sc_hs__clkbuf_8
Xsky130_fd_sc_hs__clkbuf_8_83 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__einvp_8_9/TE
+ test_mux_select[0] sky130_fd_sc_hs__clkbuf_8_83/a_125_368# sky130_fd_sc_hs__clkbuf_8
Xsky130_fd_sc_hs__clkbuf_8_94 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__clkbuf_8_95/X
+ CTL_BUF_N[3] sky130_fd_sc_hs__clkbuf_8_95/a_125_368# sky130_fd_sc_hs__clkbuf_8
Xsky130_fd_sc_hs__clkbuf_4_19 DVSS: DVDD: DVDD: DVSS: pi1_con[1] sky130_fd_sc_hs__clkbuf_4_19/X
+ sky130_fd_sc_hs__clkbuf_4_19/a_83_270# sky130_fd_sc_hs__clkbuf_4
Xsky130_fd_sc_hs__einvp_8_3 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__einvp_8_3/Z sky130_fd_sc_hs__einvp_8_3/TE
+ osc_core_1/p5 sky130_fd_sc_hs__einvp_8_3/a_802_323# sky130_fd_sc_hs__einvp_8_3/a_27_74#
+ sky130_fd_sc_hs__einvp_8_3/a_27_368# sky130_fd_sc_hs__einvp_8
Xsky130_fd_sc_hs__clkbuf_8_6 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__clkbuf_8_7/X
+ sky130_fd_sc_hs__clkbuf_8_7/A sky130_fd_sc_hs__clkbuf_8_7/a_125_368# sky130_fd_sc_hs__clkbuf_8
Xhr_16t4_mux_top_0 hr_16t4_mux_top_1/clk prbs_generator_syn_11/out prbs_generator_syn_17/out
+ prbs_generator_syn_3/out prbs_generator_syn_21/out prbs_generator_syn_7/out prbs_generator_syn_19/out
+ prbs_generator_syn_1/out hr_16t4_mux_top_1/din[8] prbs_generator_syn_5/out hr_16t4_mux_top_1/din[6]
+ hr_16t4_mux_top_1/din[5] hr_16t4_mux_top_1/din[4] prbs_generator_syn_9/out hr_16t4_mux_top_1/din[2]
+ hr_16t4_mux_top_1/din[1] hr_16t4_mux_top_1/din[0] qr_4t1_mux_top_1/rst hr_16t4_mux_top_1/clk_prbs
+ qr_4t1_mux_top_1/din[3] qr_4t1_mux_top_1/din[2] qr_4t1_mux_top_1/din[1] qr_4t1_mux_top_1/din[0]
+ DVSS: DVDD: hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_31/D hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_15/a_735_102#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_23/Q hr_16t4_mux_top_1/sky130_fd_sc_hs__clkbuf_4_1/X
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__inv_4_11/A hr_16t4_mux_top_1/sky130_fd_sc_hs__clkbuf_2_25/a_43_192#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__inv_4_19/A hr_16t4_mux_top_1/sky130_fd_sc_hs__dfrtp_4_3/a_890_138#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__buf_2_11/a_21_260# hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_1/a_1141_508#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_5/Q hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_29/a_544_485#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_39/a_696_458# hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_46/a_735_102#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_47/a_1034_424# hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_24/D
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__a22o_1_9/A2 hr_16t4_mux_top_1/sky130_fd_sc_hs__a22o_1_9/B1
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_8/a_27_74# hr_16t4_mux_top_1/sky130_fd_sc_hs__a22o_1_5/X
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_19/a_651_503# hr_16t4_mux_top_1/sky130_fd_sc_hs__a22o_1_7/X
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_33/a_735_102# hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_31/a_27_74#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_46/a_1034_424# hr_16t4_mux_top_1/sky130_fd_sc_hs__clkinv_4_1/Y
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_25/a_1141_508# hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_46/Q
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_46/D hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_35/a_1226_296#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_5/a_696_458# hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_41/Q
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_45/a_1034_424# hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_24/a_1141_508#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__clkbuf_2_11/a_43_192# hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_33/a_1226_296#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__a22o_1_15/a_230_79# hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_47/a_206_368#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_39/a_544_485# hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_13/a_735_102#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_33/Q hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_23/a_1141_508#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__clkbuf_2_15/a_43_192# hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_45/D
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_29/Q hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_35/a_206_368#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_47/a_437_503# hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_27/a_651_503#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__inv_4_1/Y hr_16t4_mux_top_1/sky130_fd_sc_hs__a22o_1_17/X
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_45/a_735_102# hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_37/a_696_458#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_41/a_1034_424# hr_16t4_mux_top_1/sky130_fd_sc_hs__a22o_1_15/a_222_392#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_39/a_1141_508# hr_16t4_mux_top_1/sky130_fd_sc_hs__a22o_1_15/a_52_123#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_3/a_651_503# hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_15/D
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_5/a_544_485# hr_16t4_mux_top_1/sky130_fd_sc_hs__clkbuf_2_19/a_43_192#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_19/a_1178_124# hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_35/a_437_503#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_18/a_651_503# hr_16t4_mux_top_1/sky130_fd_sc_hs__inv_4_5/Y
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_37/a_1141_508# hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_31/a_1226_296#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_47/D hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_1/a_206_368#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_33/a_27_74# hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_18/a_1178_124#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_15/a_206_368# hr_16t4_mux_top_1/sky130_fd_sc_hs__a22o_1_23/a_132_392#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_5/D hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_19/a_696_458#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfrtp_4_3/a_313_74# hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_25/a_735_102#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__buf_2_5/X hr_16t4_mux_top_1/sky130_fd_sc_hs__a22o_1_5/B2
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_35/Q hr_16t4_mux_top_1/sky130_fd_sc_hs__dfrtp_4_3/a_494_366#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_1/a_437_503# hr_16t4_mux_top_1/sky130_fd_sc_hs__clkbuf_4_3/a_83_270#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__clkbuf_2_9/a_43_192# hr_16t4_mux_top_1/sky130_fd_sc_hs__a22o_1_19/X
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_9/a_735_102# hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_15/a_437_503#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_46/a_206_368# hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_37/a_544_485#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfrtp_4_1/a_1647_81# hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_8/Q
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfrtp_4_1/a_890_138# hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_15/a_1178_124#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__a22o_1_21/a_230_79# hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_33/a_206_368#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__a22o_1_1/a_222_392# hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_46/a_437_503#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__clkinv_2_1/Y hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_45/a_27_74#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__a22o_1_14/a_222_392# hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_35/a_1141_508#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_9/a_1178_124# hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_13/a_1178_124#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_33/a_437_503# hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_19/a_544_485#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_27/D hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_27/a_696_458#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_33/a_1141_508# hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_8/a_1178_124#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_5/a_27_74# hr_16t4_mux_top_1/sky130_fd_sc_hs__buf_2_15/X
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__inv_4_11/Y hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_18/Q
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_3/a_696_458# hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_13/a_206_368#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__a22o_1_21/a_52_123# hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_47/a_651_503#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_3/D hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_18/a_696_458#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_24/a_735_102# hr_16t4_mux_top_1/sky130_fd_sc_hs__clkbuf_2_23/a_43_192#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_7/a_1178_124# hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_47/a_1226_296#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__a22o_1_9/a_132_392# hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_8/a_735_102#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_45/a_206_368# hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_13/a_437_503#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_35/a_651_503# hr_16t4_mux_top_1/sky130_fd_sc_hs__dfrtp_4_3/a_2010_409#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_46/a_1226_296# hr_16t4_mux_top_1/sky130_fd_sc_hs__a22o_1_1/a_230_79#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_45/Q hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_23/a_27_74#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__a22o_1_11/a_230_79# hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_29/a_1178_124#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_45/a_437_503# hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_27/a_544_485#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_37/Q hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_41/a_735_102#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_31/a_1141_508# hr_16t4_mux_top_1/sky130_fd_sc_hs__inv_4_9/Y
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_45/a_1226_296# hr_16t4_mux_top_1/sky130_fd_sc_hs__dfrtp_4_1/a_37_78#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_1/a_651_503# hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_3/a_544_485#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__a22o_1_1/X hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_25/a_206_368#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__a22o_1_5/a_230_79# hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_15/a_651_503#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_18/a_544_485# hr_16t4_mux_top_1/sky130_fd_sc_hs__a22o_1_14/a_230_79#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfrtp_4_1/a_2010_409# hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_31/a_735_102#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__a22o_1_23/X hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_5/a_1178_124#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__buf_2_11/X hr_16t4_mux_top_1/sky130_fd_sc_hs__inv_4_19/Y
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_9/a_206_368# hr_16t4_mux_top_1/sky130_fd_sc_hs__a22o_1_1/a_52_123#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_15/a_27_74# hr_16t4_mux_top_1/sky130_fd_sc_hs__a22o_1_21/a_132_392#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_7/a_27_74# hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_1/D
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__a22o_1_11/a_52_123# hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_25/a_437_503#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_46/a_651_503# hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_23/a_735_102#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__a22o_1_9/a_230_79# hr_16t4_mux_top_1/sky130_fd_sc_hs__clkbuf_2_13/a_43_192#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_31/Q hr_16t4_mux_top_1/sky130_fd_sc_hs__a22o_1_19/a_230_79#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_41/a_1226_296# hr_16t4_mux_top_1/sky130_fd_sc_hs__dfrtp_4_1/a_494_366#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_19/a_1034_424# hr_16t4_mux_top_1/sky130_fd_sc_hs__a22o_1_21/X
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_9/a_437_503# hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_7/a_735_102#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_27/a_1178_124# hr_16t4_mux_top_1/sky130_fd_sc_hs__a22o_1_11/a_132_392#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__clkbuf_2_1/a_43_192# hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_33/a_651_503#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__a22o_1_5/a_52_123# hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_47/a_696_458#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__a22o_1_14/a_52_123# hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_3/a_1178_124#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__a22o_1_23/a_222_392# hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_39/D
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_18/a_1034_424# hr_16t4_mux_top_1/sky130_fd_sc_hs__clkbuf_2_17/a_43_192#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfrtp_4_1/Q hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_35/a_696_458#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__clkbuf_2_5/a_43_192# hr_16t4_mux_top_1/sky130_fd_sc_hs__inv_4_7/Y
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__a22o_1_9/a_52_123# hr_16t4_mux_top_1/sky130_fd_sc_hs__a22o_1_19/a_52_123#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfrtp_4_3/a_699_463# hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_24/a_206_368#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_13/a_651_503# hr_16t4_mux_top_1/sky130_fd_sc_hs__inv_4_21/Y
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_47/a_1141_508# hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_1/a_1178_124#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__inv_4_13/Y hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_15/a_1034_424#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_8/a_206_368# hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_1/a_696_458#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_19/Q hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_9/a_1034_424#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_24/a_437_503# hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_1/a_27_74#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_45/a_651_503# hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_47/a_544_485#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_15/a_696_458# hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_46/a_1141_508#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__buf_2_14/X hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_9/D
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_13/a_1034_424# hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_19/a_27_74#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__a22o_1_7/a_132_392# hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_8/a_437_503#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_27/Q hr_16t4_mux_top_1/sky130_fd_sc_hs__buf_2_9/X
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_25/a_1178_124# hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_8/a_1034_424#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_41/a_206_368# hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_35/a_544_485#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_46/a_696_458# hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_45/a_1141_508#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_24/a_1178_124# hr_16t4_mux_top_1/sky130_fd_sc_hs__a22o_1_9/a_222_392#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_7/a_1034_424# hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_31/a_206_368#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_25/a_651_503# hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_41/a_437_503#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_33/a_696_458# hr_16t4_mux_top_1/sky130_fd_sc_hs__buf_2_3/a_21_260#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_25/D hr_16t4_mux_top_1/sky130_fd_sc_hs__a22o_1_7/A2
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_9/a_651_503# hr_16t4_mux_top_1/sky130_fd_sc_hs__clkbuf_1_1/a_27_74#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_1/a_544_485# hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_23/a_1178_124#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_27/a_27_74# hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_23/a_206_368#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_31/a_437_503# hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_15/a_544_485#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_41/a_1141_508# hr_16t4_mux_top_1/sky130_fd_sc_hs__dfrtp_4_3/a_124_78#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_47/Q hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_29/a_1034_424#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__buf_2_7/a_21_260# hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_7/a_206_368#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_39/a_1178_124# hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_23/a_437_503#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_7/Q hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_46/a_544_485#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_13/a_696_458# hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_29/a_735_102#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__clkbuf_2_27/a_43_192# hr_16t4_mux_top_1/sky130_fd_sc_hs__a22o_1_3/X
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__buf_2_15/a_21_260# hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_7/a_437_503#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_37/a_1178_124# hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_5/a_1034_424#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_33/a_544_485# hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_45/a_696_458#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfrtp_4_3/a_1827_81# hr_16t4_mux_top_1/sky130_fd_sc_hs__a22o_1_21/a_222_392#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__a22o_1_3/a_230_79# hr_16t4_mux_top_1/sky130_fd_sc_hs__inv_4_17/Y
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_24/a_651_503# hr_16t4_mux_top_1/sky130_fd_sc_hs__inv_4_3/Y
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__a22o_1_11/a_222_392# hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_27/a_1034_424#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_19/a_1226_296# hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_8/a_651_503#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfrtp_4_1/a_699_463# hr_16t4_mux_top_1/sky130_fd_sc_hs__buf_2_7/X
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_3/a_1034_424# hr_16t4_mux_top_1/sky130_fd_sc_hs__a22o_1_17/a_230_79#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_13/a_544_485# hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_25/a_696_458#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_39/a_735_102# hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_29/a_27_74#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_18/a_1226_296# hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_9/a_696_458#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__a22o_1_3/a_52_123# hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_35/a_1178_124#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_47/a_27_74# hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_3/Q
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_41/a_651_503# hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_45/a_544_485#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_35/D hr_16t4_mux_top_1/sky130_fd_sc_hs__dfrtp_4_3/a_789_463#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__a22o_1_5/a_132_392# hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_33/a_1178_124#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_5/a_735_102# hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_1/a_1034_424#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__a22o_1_19/a_132_392# hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_13/a_27_74#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_31/a_651_503# hr_16t4_mux_top_1/sky130_fd_sc_hs__a22o_1_17/a_52_123#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfrtp_4_1/a_313_74# hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_23/D
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_15/a_1226_296# hr_16t4_mux_top_1/sky130_fd_sc_hs__clkbuf_2_31/a_43_192#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__inv_4_15/Y hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_39/a_27_74#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__a22o_1_7/a_222_392# hr_16t4_mux_top_1/sky130_fd_sc_hs__clkbuf_4_1/a_83_270#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_23/a_651_503# hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_25/a_544_485#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__clkbuf_2_7/a_43_192# hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_9/a_1226_296#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_8/D hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_25/a_1034_424#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfrtp_4_3/a_834_355# hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_13/a_1226_296#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_7/a_651_503# hr_16t4_mux_top_1/sky130_fd_sc_hs__dfrtp_4_3/a_1627_493#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_9/a_544_485# hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_29/a_206_368#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfrtp_4_3/a_812_138# hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_24/a_696_458#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_8/a_1226_296# hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_37/a_735_102#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_24/a_1034_424# hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_25/a_27_74#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_31/a_1178_124# hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_8/a_696_458#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_1/Q hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_29/a_437_503#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_7/a_1226_296# hr_16t4_mux_top_1/sky130_fd_sc_hs__dfrtp_4_3/a_37_78#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_23/a_1034_424# hr_16t4_mux_top_1/sky130_fd_sc_hs__a22o_1_23/a_230_79#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__a22o_1_3/a_132_392# hr_16t4_mux_top_1/sky130_fd_sc_hs__dfrtp_4_1/a_1627_493#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__a22o_1_17/a_132_392# hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_19/a_735_102#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_41/a_696_458# hr_16t4_mux_top_1/sky130_fd_sc_hs__dfrtp_4_1/a_1827_81#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_39/a_1034_424# hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_19/a_1141_508#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_9/a_27_74# hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_29/a_1226_296#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_18/a_27_74# hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_39/a_206_368#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_24/a_544_485# hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_31/a_696_458#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_37/a_1034_424# hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_18/a_1141_508#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_9/Q hr_16t4_mux_top_1/sky130_fd_sc_hs__a22o_1_23/a_52_123#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_8/a_544_485# hr_16t4_mux_top_1/sky130_fd_sc_hs__buf_2_3/X
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__buf_2_14/a_21_260# hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_5/a_1226_296#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_39/a_437_503# hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_23/a_696_458#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__buf_2_9/a_21_260# hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_5/a_206_368#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_7/a_696_458# hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_39/Q
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfrtp_4_3/a_1678_395# hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_41/a_544_485#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__clkbuf_2_29/a_43_192# hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_27/a_735_102#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfrtp_4_1/a_789_463# hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_15/a_1141_508#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__buf_2_1/X hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_41/a_27_74#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_5/a_437_503# hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_27/a_1226_296#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_3/a_735_102# hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_47/a_1178_124#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_9/a_1141_508# hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_3/a_1226_296#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_18/a_735_102# hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_31/a_544_485#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_35/a_1034_424# hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_13/a_1141_508#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__a22o_1_7/a_230_79# hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_3/a_27_74#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_46/a_1178_124# hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_8/a_1141_508#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfrtp_4_1/a_1678_395# hr_16t4_mux_top_1/sky130_fd_sc_hs__a22o_1_5/a_222_392#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_37/a_206_368# hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_23/a_544_485#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_29/a_651_503# hr_16t4_mux_top_1/sky130_fd_sc_hs__a22o_1_7/B2
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__a22o_1_19/a_222_392# hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_33/a_1034_424#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfrtp_4_1/a_834_355# hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_35/a_27_74#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_7/a_544_485# hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_45/a_1178_124#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_7/a_1141_508# hr_16t4_mux_top_1/sky130_fd_sc_hs__dfrtp_4_1/a_812_138#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_1/a_1226_296# hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_37/a_437_503#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__clkbuf_2_3/a_43_192# hr_16t4_mux_top_1/sky130_fd_sc_hs__a22o_1_7/a_52_123#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfrtp_4_3/a_1350_392# hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_19/a_206_368#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_29/a_1141_508# hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_25/a_1226_296#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_41/a_1178_124# hr_16t4_mux_top_1/sky130_fd_sc_hs__a22o_1_15/a_132_392#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_19/a_437_503# hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_46/a_27_74#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_39/a_651_503# hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_31/a_1034_424#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_24/a_1226_296# hr_16t4_mux_top_1/sky130_fd_sc_hs__dfrtp_4_1/a_1350_392#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_5/a_1141_508# hr_16t4_mux_top_1/sky130_fd_sc_hs__a22o_1_3/a_222_392#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__clkbuf_16_1/a_114_74# hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_47/a_735_102#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__a22o_1_17/a_222_392# hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_23/a_1226_296#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_5/a_651_503# hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_27/a_206_368#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_37/a_27_74# hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_29/a_696_458#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_35/a_735_102# hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_27/a_1141_508#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_3/a_206_368# hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_39/a_1226_296#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__buf_2_1/a_21_260# hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_3/a_1141_508#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_18/a_206_368# hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_27/a_437_503#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__clkbuf_2_21/a_43_192# hr_16t4_mux_top_1/sky130_fd_sc_hs__a22o_1_1/a_132_392#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_3/a_437_503# hr_16t4_mux_top_1/sky130_fd_sc_hs__dfrtp_4_1/a_124_78#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_37/a_1226_296# hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_24/a_27_74#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_1/a_735_102# hr_16t4_mux_top_1/sky130_fd_sc_hs__buf_2_5/a_21_260#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__a22o_1_14/a_132_392# hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_37/a_651_503#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_18/a_437_503# hr_16t4_mux_top_1/sky130_fd_sc_hs__dfrtp_4_3/a_1647_81#
+ hr_16t4_mux_top
Xsky130_fd_sc_hs__clkinv_8_6 DVSS: DVDD: DVDD: DVSS: hr_16t4_mux_top_1/din[5] hr_16t4_mux_top_3/din[5]
+ sky130_fd_sc_hs__clkinv_8
Xsky130_fd_sc_hs__clkbuf_4_0 DVSS: DVDD: DVDD: DVSS: pi3_con[3] sky130_fd_sc_hs__clkbuf_4_1/X
+ sky130_fd_sc_hs__clkbuf_4_1/a_83_270# sky130_fd_sc_hs__clkbuf_4
Xsky130_fd_sc_hs__clkinv_4_0 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__nand2_2_27/B
+ sky130_fd_sc_hs__dlrtp_1_24/D sky130_fd_sc_hs__clkinv_4
Xsky130_fd_sc_hs__conb_1_109 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__conb_1_109/LO
+ sky130_fd_sc_hs__conb_1_109/HI sky130_fd_sc_hs__conb_1_109/a_165_290# sky130_fd_sc_hs__conb_1_109/a_21_290#
+ sky130_fd_sc_hs__conb_1
Xsky130_fd_sc_hs__dlrtp_1_110 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__dlrtp_1_111/Q
+ sky130_fd_sc_hs__dlrtp_1_9/GATE sky130_fd_sc_hs__conb_1_131/HI sky130_fd_sc_hs__o21ai_2_39/Y
+ sky130_fd_sc_hs__dlrtp_1_111/a_216_424# sky130_fd_sc_hs__dlrtp_1_111/a_759_508#
+ sky130_fd_sc_hs__dlrtp_1_111/a_565_74# sky130_fd_sc_hs__dlrtp_1_111/a_27_424# sky130_fd_sc_hs__dlrtp_1_111/a_1045_74#
+ sky130_fd_sc_hs__dlrtp_1_111/a_643_74# sky130_fd_sc_hs__dlrtp_1_111/a_817_48# sky130_fd_sc_hs__dlrtp_1_111/a_568_392#
+ sky130_fd_sc_hs__dlrtp_1_111/a_363_74# sky130_fd_sc_hs__dlrtp_1_111/a_769_74# sky130_fd_sc_hs__dlrtp_1
Xsky130_fd_sc_hs__dlrtp_1_121 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__dlrtp_1_121/Q
+ sky130_fd_sc_hs__dlrtp_1_9/GATE sky130_fd_sc_hs__conb_1_131/HI sky130_fd_sc_hs__dlrtp_1_121/D
+ sky130_fd_sc_hs__dlrtp_1_121/a_216_424# sky130_fd_sc_hs__dlrtp_1_121/a_759_508#
+ sky130_fd_sc_hs__dlrtp_1_121/a_565_74# sky130_fd_sc_hs__dlrtp_1_121/a_27_424# sky130_fd_sc_hs__dlrtp_1_121/a_1045_74#
+ sky130_fd_sc_hs__dlrtp_1_121/a_643_74# sky130_fd_sc_hs__dlrtp_1_121/a_817_48# sky130_fd_sc_hs__dlrtp_1_121/a_568_392#
+ sky130_fd_sc_hs__dlrtp_1_121/a_363_74# sky130_fd_sc_hs__dlrtp_1_121/a_769_74# sky130_fd_sc_hs__dlrtp_1
Xsky130_fd_sc_hs__dlrtp_1_132 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__dlrtp_1_133/Q
+ sky130_fd_sc_hs__clkbuf_2_3/A sky130_fd_sc_hs__conb_1_135/HI sky130_fd_sc_hs__dlrtp_1_133/D
+ sky130_fd_sc_hs__dlrtp_1_133/a_216_424# sky130_fd_sc_hs__dlrtp_1_133/a_759_508#
+ sky130_fd_sc_hs__dlrtp_1_133/a_565_74# sky130_fd_sc_hs__dlrtp_1_133/a_27_424# sky130_fd_sc_hs__dlrtp_1_133/a_1045_74#
+ sky130_fd_sc_hs__dlrtp_1_133/a_643_74# sky130_fd_sc_hs__dlrtp_1_133/a_817_48# sky130_fd_sc_hs__dlrtp_1_133/a_568_392#
+ sky130_fd_sc_hs__dlrtp_1_133/a_363_74# sky130_fd_sc_hs__dlrtp_1_133/a_769_74# sky130_fd_sc_hs__dlrtp_1
Xsky130_fd_sc_hs__dlrtp_1_143 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__dlrtp_1_143/Q
+ sky130_fd_sc_hs__clkbuf_16_53/X sky130_fd_sc_hs__conb_1_127/HI sky130_fd_sc_hs__dlrtp_1_143/D
+ sky130_fd_sc_hs__dlrtp_1_143/a_216_424# sky130_fd_sc_hs__dlrtp_1_143/a_759_508#
+ sky130_fd_sc_hs__dlrtp_1_143/a_565_74# sky130_fd_sc_hs__dlrtp_1_143/a_27_424# sky130_fd_sc_hs__dlrtp_1_143/a_1045_74#
+ sky130_fd_sc_hs__dlrtp_1_143/a_643_74# sky130_fd_sc_hs__dlrtp_1_143/a_817_48# sky130_fd_sc_hs__dlrtp_1_143/a_568_392#
+ sky130_fd_sc_hs__dlrtp_1_143/a_363_74# sky130_fd_sc_hs__dlrtp_1_143/a_769_74# sky130_fd_sc_hs__dlrtp_1
Xsky130_fd_sc_hs__dlrtp_1_154 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__buf_2_155/A
+ sky130_fd_sc_hs__clkbuf_16_53/X sky130_fd_sc_hs__conb_1_137/HI sky130_fd_sc_hs__buf_2_163/X
+ sky130_fd_sc_hs__dlrtp_1_156/a_216_424# sky130_fd_sc_hs__dlrtp_1_156/a_759_508#
+ sky130_fd_sc_hs__dlrtp_1_156/a_565_74# sky130_fd_sc_hs__dlrtp_1_156/a_27_424# sky130_fd_sc_hs__dlrtp_1_156/a_1045_74#
+ sky130_fd_sc_hs__dlrtp_1_156/a_643_74# sky130_fd_sc_hs__dlrtp_1_156/a_817_48# sky130_fd_sc_hs__dlrtp_1_156/a_568_392#
+ sky130_fd_sc_hs__dlrtp_1_156/a_363_74# sky130_fd_sc_hs__dlrtp_1_156/a_769_74# sky130_fd_sc_hs__dlrtp_1
Xsky130_fd_sc_hs__inv_4_2 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__inv_4_3/Y ref_clk_ext_n
+ sky130_fd_sc_hs__inv_4
Xsky130_fd_sc_hs__clkbuf_2_30 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__einvp_2_3/TE
+ sky130_fd_sc_hs__dlrtp_1_91/Q sky130_fd_sc_hs__clkbuf_2_31/a_43_192# sky130_fd_sc_hs__clkbuf_2
Xsky130_fd_sc_hs__clkbuf_2_41 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__dlrtp_1_107/D
+ sky130_fd_sc_hs__buf_2_113/X sky130_fd_sc_hs__clkbuf_2_41/a_43_192# sky130_fd_sc_hs__clkbuf_2
Xsky130_fd_sc_hs__clkbuf_2_52 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__dlrtp_1_29/D
+ sky130_fd_sc_hs__o21bai_2_53/Y sky130_fd_sc_hs__clkbuf_2_53/a_43_192# sky130_fd_sc_hs__clkbuf_2
Xsky130_fd_sc_hs__clkbuf_2_63 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__einvp_8_1/TE
+ sky130_fd_sc_hs__einvp_8_3/TE sky130_fd_sc_hs__clkbuf_2_63/a_43_192# sky130_fd_sc_hs__clkbuf_2
Xsky130_fd_sc_hs__einvp_2_109 DVSS: DVDD: DVDD: DVSS: dout_n sky130_fd_sc_hs__einvp_2_9/A
+ sky130_fd_sc_hs__dlrtp_1_95/Q sky130_fd_sc_hs__einvp_2_109/a_263_323# sky130_fd_sc_hs__einvp_2_109/a_36_74#
+ sky130_fd_sc_hs__einvp_2_109/a_27_368# sky130_fd_sc_hs__einvp_2
Xsky130_fd_sc_hs__clkbuf_16_9 DVSS: DVDD: DVDD: DVSS: prbs_generator_syn_9/inj_err
+ sky130_fd_sc_hs__clkbuf_4_39/X sky130_fd_sc_hs__clkbuf_16_9/a_114_74# sky130_fd_sc_hs__clkbuf_16
Xsky130_fd_sc_hs__dlrtp_1_1 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__dlrtp_1_1/Q sky130_fd_sc_hs__dlrtp_1_9/GATE
+ sky130_fd_sc_hs__conb_1_117/HI sky130_fd_sc_hs__buf_2_81/X sky130_fd_sc_hs__dlrtp_1_1/a_216_424#
+ sky130_fd_sc_hs__dlrtp_1_1/a_759_508# sky130_fd_sc_hs__dlrtp_1_1/a_565_74# sky130_fd_sc_hs__dlrtp_1_1/a_27_424#
+ sky130_fd_sc_hs__dlrtp_1_1/a_1045_74# sky130_fd_sc_hs__dlrtp_1_1/a_643_74# sky130_fd_sc_hs__dlrtp_1_1/a_817_48#
+ sky130_fd_sc_hs__dlrtp_1_1/a_568_392# sky130_fd_sc_hs__dlrtp_1_1/a_363_74# sky130_fd_sc_hs__dlrtp_1_1/a_769_74#
+ sky130_fd_sc_hs__dlrtp_1
Xsky130_fd_sc_hs__buf_2_70 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__buf_2_71/A sky130_fd_sc_hs__buf_2_71/X
+ sky130_fd_sc_hs__buf_2_71/a_21_260# sky130_fd_sc_hs__buf_2
Xsky130_fd_sc_hs__buf_2_81 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__buf_2_83/X sky130_fd_sc_hs__buf_2_81/X
+ sky130_fd_sc_hs__buf_2_81/a_21_260# sky130_fd_sc_hs__buf_2
Xsky130_fd_sc_hs__buf_2_92 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__buf_2_93/A sky130_fd_sc_hs__buf_2_93/X
+ sky130_fd_sc_hs__buf_2_93/a_21_260# sky130_fd_sc_hs__buf_2
Xsky130_fd_sc_hs__o21bai_2_50 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__clkinv_4_5/Y
+ sky130_fd_sc_hs__nand2_2_21/B sky130_fd_sc_hs__dlrtp_1_29/D sky130_fd_sc_hs__buf_2_127/A
+ sky130_fd_sc_hs__o21bai_2_51/a_27_74# sky130_fd_sc_hs__o21bai_2_51/a_225_74# sky130_fd_sc_hs__o21bai_2_51/a_507_368#
+ sky130_fd_sc_hs__o21bai_2
Xsky130_fd_sc_hs__o21bai_2_61 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__inv_8_1/Y sky130_fd_sc_hs__nand2_2_5/B
+ sky130_fd_sc_hs__dlrtp_1_143/D sky130_fd_sc_hs__o21bai_2_61/Y sky130_fd_sc_hs__o21bai_2_61/a_27_74#
+ sky130_fd_sc_hs__o21bai_2_61/a_225_74# sky130_fd_sc_hs__o21bai_2_61/a_507_368# sky130_fd_sc_hs__o21bai_2
Xsky130_fd_sc_hs__conb_1_270 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__conb_1_271/LO
+ sky130_fd_sc_hs__conb_1_271/HI sky130_fd_sc_hs__conb_1_271/a_165_290# sky130_fd_sc_hs__conb_1_271/a_21_290#
+ sky130_fd_sc_hs__conb_1
Xsky130_fd_sc_hs__clkbuf_8_40 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__or2b_4_1/A
+ sky130_fd_sc_hs__nand2_2_23/Y sky130_fd_sc_hs__clkbuf_8_41/a_125_368# sky130_fd_sc_hs__clkbuf_8
Xsky130_fd_sc_hs__clkbuf_8_51 DVSS: DVDD: DVDD: DVSS: qr_4t1_mux_top_3/clk_Q sky130_fd_sc_hs__einvn_8_1/Z
+ sky130_fd_sc_hs__clkbuf_8_51/a_125_368# sky130_fd_sc_hs__clkbuf_8
Xsky130_fd_sc_hs__clkbuf_8_62 DVSS: DVDD: DVDD: DVSS: osc_core_1/con_perb_5[2] con_perb[2]
+ sky130_fd_sc_hs__clkbuf_8_63/a_125_368# sky130_fd_sc_hs__clkbuf_8
Xsky130_fd_sc_hs__clkbuf_8_73 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__nor2_4_3/A
+ sky130_fd_sc_hs__clkbuf_8_77/X sky130_fd_sc_hs__clkbuf_8_73/a_125_368# sky130_fd_sc_hs__clkbuf_8
Xsky130_fd_sc_hs__clkbuf_8_84 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__einvp_8_11/TE
+ test_mux_select[1] sky130_fd_sc_hs__clkbuf_8_85/a_125_368# sky130_fd_sc_hs__clkbuf_8
Xsky130_fd_sc_hs__clkbuf_8_95 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__clkbuf_8_95/X
+ CTL_BUF_N[3] sky130_fd_sc_hs__clkbuf_8_95/a_125_368# sky130_fd_sc_hs__clkbuf_8
Xsky130_fd_sc_hs__einvp_8_4 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__inv_4_39/A sky130_fd_sc_hs__einvp_8_5/TE
+ sky130_fd_sc_hs__einvp_8_5/A sky130_fd_sc_hs__einvp_8_5/a_802_323# sky130_fd_sc_hs__einvp_8_5/a_27_74#
+ sky130_fd_sc_hs__einvp_8_5/a_27_368# sky130_fd_sc_hs__einvp_8
Xsky130_fd_sc_hs__clkbuf_8_7 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__clkbuf_8_7/X
+ sky130_fd_sc_hs__clkbuf_8_7/A sky130_fd_sc_hs__clkbuf_8_7/a_125_368# sky130_fd_sc_hs__clkbuf_8
Xhr_16t4_mux_top_1 hr_16t4_mux_top_1/clk prbs_generator_syn_11/out prbs_generator_syn_17/out
+ prbs_generator_syn_3/out prbs_generator_syn_21/out prbs_generator_syn_7/out prbs_generator_syn_19/out
+ prbs_generator_syn_1/out hr_16t4_mux_top_1/din[8] prbs_generator_syn_5/out hr_16t4_mux_top_1/din[6]
+ hr_16t4_mux_top_1/din[5] hr_16t4_mux_top_1/din[4] prbs_generator_syn_9/out hr_16t4_mux_top_1/din[2]
+ hr_16t4_mux_top_1/din[1] hr_16t4_mux_top_1/din[0] qr_4t1_mux_top_1/rst hr_16t4_mux_top_1/clk_prbs
+ qr_4t1_mux_top_1/din[3] qr_4t1_mux_top_1/din[2] qr_4t1_mux_top_1/din[1] qr_4t1_mux_top_1/din[0]
+ DVSS: DVDD: hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_31/D hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_15/a_735_102#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_23/Q hr_16t4_mux_top_1/sky130_fd_sc_hs__clkbuf_4_1/X
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__inv_4_11/A hr_16t4_mux_top_1/sky130_fd_sc_hs__clkbuf_2_25/a_43_192#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__inv_4_19/A hr_16t4_mux_top_1/sky130_fd_sc_hs__dfrtp_4_3/a_890_138#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__buf_2_11/a_21_260# hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_1/a_1141_508#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_5/Q hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_29/a_544_485#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_39/a_696_458# hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_46/a_735_102#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_47/a_1034_424# hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_24/D
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__a22o_1_9/A2 hr_16t4_mux_top_1/sky130_fd_sc_hs__a22o_1_9/B1
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_8/a_27_74# hr_16t4_mux_top_1/sky130_fd_sc_hs__a22o_1_5/X
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_19/a_651_503# hr_16t4_mux_top_1/sky130_fd_sc_hs__a22o_1_7/X
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_33/a_735_102# hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_31/a_27_74#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_46/a_1034_424# hr_16t4_mux_top_1/sky130_fd_sc_hs__clkinv_4_1/Y
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_25/a_1141_508# hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_46/Q
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_46/D hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_35/a_1226_296#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_5/a_696_458# hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_41/Q
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_45/a_1034_424# hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_24/a_1141_508#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__clkbuf_2_11/a_43_192# hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_33/a_1226_296#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__a22o_1_15/a_230_79# hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_47/a_206_368#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_39/a_544_485# hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_13/a_735_102#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_33/Q hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_23/a_1141_508#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__clkbuf_2_15/a_43_192# hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_45/D
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_29/Q hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_35/a_206_368#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_47/a_437_503# hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_27/a_651_503#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__inv_4_1/Y hr_16t4_mux_top_1/sky130_fd_sc_hs__a22o_1_17/X
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_45/a_735_102# hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_37/a_696_458#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_41/a_1034_424# hr_16t4_mux_top_1/sky130_fd_sc_hs__a22o_1_15/a_222_392#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_39/a_1141_508# hr_16t4_mux_top_1/sky130_fd_sc_hs__a22o_1_15/a_52_123#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_3/a_651_503# hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_15/D
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_5/a_544_485# hr_16t4_mux_top_1/sky130_fd_sc_hs__clkbuf_2_19/a_43_192#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_19/a_1178_124# hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_35/a_437_503#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_18/a_651_503# hr_16t4_mux_top_1/sky130_fd_sc_hs__inv_4_5/Y
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_37/a_1141_508# hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_31/a_1226_296#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_47/D hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_1/a_206_368#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_33/a_27_74# hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_18/a_1178_124#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_15/a_206_368# hr_16t4_mux_top_1/sky130_fd_sc_hs__a22o_1_23/a_132_392#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_5/D hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_19/a_696_458#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfrtp_4_3/a_313_74# hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_25/a_735_102#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__buf_2_5/X hr_16t4_mux_top_1/sky130_fd_sc_hs__a22o_1_5/B2
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_35/Q hr_16t4_mux_top_1/sky130_fd_sc_hs__dfrtp_4_3/a_494_366#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_1/a_437_503# hr_16t4_mux_top_1/sky130_fd_sc_hs__clkbuf_4_3/a_83_270#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__clkbuf_2_9/a_43_192# hr_16t4_mux_top_1/sky130_fd_sc_hs__a22o_1_19/X
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_9/a_735_102# hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_15/a_437_503#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_46/a_206_368# hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_37/a_544_485#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfrtp_4_1/a_1647_81# hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_8/Q
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfrtp_4_1/a_890_138# hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_15/a_1178_124#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__a22o_1_21/a_230_79# hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_33/a_206_368#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__a22o_1_1/a_222_392# hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_46/a_437_503#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__clkinv_2_1/Y hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_45/a_27_74#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__a22o_1_14/a_222_392# hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_35/a_1141_508#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_9/a_1178_124# hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_13/a_1178_124#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_33/a_437_503# hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_19/a_544_485#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_27/D hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_27/a_696_458#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_33/a_1141_508# hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_8/a_1178_124#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_5/a_27_74# hr_16t4_mux_top_1/sky130_fd_sc_hs__buf_2_15/X
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__inv_4_11/Y hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_18/Q
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_3/a_696_458# hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_13/a_206_368#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__a22o_1_21/a_52_123# hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_47/a_651_503#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_3/D hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_18/a_696_458#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_24/a_735_102# hr_16t4_mux_top_1/sky130_fd_sc_hs__clkbuf_2_23/a_43_192#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_7/a_1178_124# hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_47/a_1226_296#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__a22o_1_9/a_132_392# hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_8/a_735_102#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_45/a_206_368# hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_13/a_437_503#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_35/a_651_503# hr_16t4_mux_top_1/sky130_fd_sc_hs__dfrtp_4_3/a_2010_409#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_46/a_1226_296# hr_16t4_mux_top_1/sky130_fd_sc_hs__a22o_1_1/a_230_79#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_45/Q hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_23/a_27_74#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__a22o_1_11/a_230_79# hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_29/a_1178_124#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_45/a_437_503# hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_27/a_544_485#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_37/Q hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_41/a_735_102#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_31/a_1141_508# hr_16t4_mux_top_1/sky130_fd_sc_hs__inv_4_9/Y
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_45/a_1226_296# hr_16t4_mux_top_1/sky130_fd_sc_hs__dfrtp_4_1/a_37_78#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_1/a_651_503# hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_3/a_544_485#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__a22o_1_1/X hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_25/a_206_368#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__a22o_1_5/a_230_79# hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_15/a_651_503#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_18/a_544_485# hr_16t4_mux_top_1/sky130_fd_sc_hs__a22o_1_14/a_230_79#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfrtp_4_1/a_2010_409# hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_31/a_735_102#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__a22o_1_23/X hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_5/a_1178_124#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__buf_2_11/X hr_16t4_mux_top_1/sky130_fd_sc_hs__inv_4_19/Y
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_9/a_206_368# hr_16t4_mux_top_1/sky130_fd_sc_hs__a22o_1_1/a_52_123#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_15/a_27_74# hr_16t4_mux_top_1/sky130_fd_sc_hs__a22o_1_21/a_132_392#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_7/a_27_74# hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_1/D
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__a22o_1_11/a_52_123# hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_25/a_437_503#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_46/a_651_503# hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_23/a_735_102#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__a22o_1_9/a_230_79# hr_16t4_mux_top_1/sky130_fd_sc_hs__clkbuf_2_13/a_43_192#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_31/Q hr_16t4_mux_top_1/sky130_fd_sc_hs__a22o_1_19/a_230_79#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_41/a_1226_296# hr_16t4_mux_top_1/sky130_fd_sc_hs__dfrtp_4_1/a_494_366#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_19/a_1034_424# hr_16t4_mux_top_1/sky130_fd_sc_hs__a22o_1_21/X
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_9/a_437_503# hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_7/a_735_102#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_27/a_1178_124# hr_16t4_mux_top_1/sky130_fd_sc_hs__a22o_1_11/a_132_392#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__clkbuf_2_1/a_43_192# hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_33/a_651_503#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__a22o_1_5/a_52_123# hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_47/a_696_458#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__a22o_1_14/a_52_123# hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_3/a_1178_124#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__a22o_1_23/a_222_392# hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_39/D
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_18/a_1034_424# hr_16t4_mux_top_1/sky130_fd_sc_hs__clkbuf_2_17/a_43_192#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfrtp_4_1/Q hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_35/a_696_458#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__clkbuf_2_5/a_43_192# hr_16t4_mux_top_1/sky130_fd_sc_hs__inv_4_7/Y
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__a22o_1_9/a_52_123# hr_16t4_mux_top_1/sky130_fd_sc_hs__a22o_1_19/a_52_123#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfrtp_4_3/a_699_463# hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_24/a_206_368#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_13/a_651_503# hr_16t4_mux_top_1/sky130_fd_sc_hs__inv_4_21/Y
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_47/a_1141_508# hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_1/a_1178_124#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__inv_4_13/Y hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_15/a_1034_424#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_8/a_206_368# hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_1/a_696_458#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_19/Q hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_9/a_1034_424#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_24/a_437_503# hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_1/a_27_74#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_45/a_651_503# hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_47/a_544_485#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_15/a_696_458# hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_46/a_1141_508#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__buf_2_14/X hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_9/D
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_13/a_1034_424# hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_19/a_27_74#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__a22o_1_7/a_132_392# hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_8/a_437_503#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_27/Q hr_16t4_mux_top_1/sky130_fd_sc_hs__buf_2_9/X
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_25/a_1178_124# hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_8/a_1034_424#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_41/a_206_368# hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_35/a_544_485#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_46/a_696_458# hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_45/a_1141_508#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_24/a_1178_124# hr_16t4_mux_top_1/sky130_fd_sc_hs__a22o_1_9/a_222_392#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_7/a_1034_424# hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_31/a_206_368#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_25/a_651_503# hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_41/a_437_503#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_33/a_696_458# hr_16t4_mux_top_1/sky130_fd_sc_hs__buf_2_3/a_21_260#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_25/D hr_16t4_mux_top_1/sky130_fd_sc_hs__a22o_1_7/A2
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_9/a_651_503# hr_16t4_mux_top_1/sky130_fd_sc_hs__clkbuf_1_1/a_27_74#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_1/a_544_485# hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_23/a_1178_124#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_27/a_27_74# hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_23/a_206_368#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_31/a_437_503# hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_15/a_544_485#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_41/a_1141_508# hr_16t4_mux_top_1/sky130_fd_sc_hs__dfrtp_4_3/a_124_78#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_47/Q hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_29/a_1034_424#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__buf_2_7/a_21_260# hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_7/a_206_368#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_39/a_1178_124# hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_23/a_437_503#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_7/Q hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_46/a_544_485#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_13/a_696_458# hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_29/a_735_102#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__clkbuf_2_27/a_43_192# hr_16t4_mux_top_1/sky130_fd_sc_hs__a22o_1_3/X
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__buf_2_15/a_21_260# hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_7/a_437_503#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_37/a_1178_124# hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_5/a_1034_424#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_33/a_544_485# hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_45/a_696_458#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfrtp_4_3/a_1827_81# hr_16t4_mux_top_1/sky130_fd_sc_hs__a22o_1_21/a_222_392#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__a22o_1_3/a_230_79# hr_16t4_mux_top_1/sky130_fd_sc_hs__inv_4_17/Y
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_24/a_651_503# hr_16t4_mux_top_1/sky130_fd_sc_hs__inv_4_3/Y
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__a22o_1_11/a_222_392# hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_27/a_1034_424#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_19/a_1226_296# hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_8/a_651_503#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfrtp_4_1/a_699_463# hr_16t4_mux_top_1/sky130_fd_sc_hs__buf_2_7/X
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_3/a_1034_424# hr_16t4_mux_top_1/sky130_fd_sc_hs__a22o_1_17/a_230_79#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_13/a_544_485# hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_25/a_696_458#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_39/a_735_102# hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_29/a_27_74#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_18/a_1226_296# hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_9/a_696_458#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__a22o_1_3/a_52_123# hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_35/a_1178_124#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_47/a_27_74# hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_3/Q
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_41/a_651_503# hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_45/a_544_485#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_35/D hr_16t4_mux_top_1/sky130_fd_sc_hs__dfrtp_4_3/a_789_463#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__a22o_1_5/a_132_392# hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_33/a_1178_124#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_5/a_735_102# hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_1/a_1034_424#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__a22o_1_19/a_132_392# hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_13/a_27_74#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_31/a_651_503# hr_16t4_mux_top_1/sky130_fd_sc_hs__a22o_1_17/a_52_123#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfrtp_4_1/a_313_74# hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_23/D
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_15/a_1226_296# hr_16t4_mux_top_1/sky130_fd_sc_hs__clkbuf_2_31/a_43_192#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__inv_4_15/Y hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_39/a_27_74#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__a22o_1_7/a_222_392# hr_16t4_mux_top_1/sky130_fd_sc_hs__clkbuf_4_1/a_83_270#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_23/a_651_503# hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_25/a_544_485#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__clkbuf_2_7/a_43_192# hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_9/a_1226_296#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_8/D hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_25/a_1034_424#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfrtp_4_3/a_834_355# hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_13/a_1226_296#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_7/a_651_503# hr_16t4_mux_top_1/sky130_fd_sc_hs__dfrtp_4_3/a_1627_493#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_9/a_544_485# hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_29/a_206_368#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfrtp_4_3/a_812_138# hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_24/a_696_458#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_8/a_1226_296# hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_37/a_735_102#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_24/a_1034_424# hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_25/a_27_74#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_31/a_1178_124# hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_8/a_696_458#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_1/Q hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_29/a_437_503#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_7/a_1226_296# hr_16t4_mux_top_1/sky130_fd_sc_hs__dfrtp_4_3/a_37_78#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_23/a_1034_424# hr_16t4_mux_top_1/sky130_fd_sc_hs__a22o_1_23/a_230_79#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__a22o_1_3/a_132_392# hr_16t4_mux_top_1/sky130_fd_sc_hs__dfrtp_4_1/a_1627_493#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__a22o_1_17/a_132_392# hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_19/a_735_102#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_41/a_696_458# hr_16t4_mux_top_1/sky130_fd_sc_hs__dfrtp_4_1/a_1827_81#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_39/a_1034_424# hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_19/a_1141_508#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_9/a_27_74# hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_29/a_1226_296#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_18/a_27_74# hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_39/a_206_368#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_24/a_544_485# hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_31/a_696_458#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_37/a_1034_424# hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_18/a_1141_508#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_9/Q hr_16t4_mux_top_1/sky130_fd_sc_hs__a22o_1_23/a_52_123#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_8/a_544_485# hr_16t4_mux_top_1/sky130_fd_sc_hs__buf_2_3/X
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__buf_2_14/a_21_260# hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_5/a_1226_296#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_39/a_437_503# hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_23/a_696_458#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__buf_2_9/a_21_260# hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_5/a_206_368#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_7/a_696_458# hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_39/Q
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfrtp_4_3/a_1678_395# hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_41/a_544_485#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__clkbuf_2_29/a_43_192# hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_27/a_735_102#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfrtp_4_1/a_789_463# hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_15/a_1141_508#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__buf_2_1/X hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_41/a_27_74#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_5/a_437_503# hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_27/a_1226_296#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_3/a_735_102# hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_47/a_1178_124#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_9/a_1141_508# hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_3/a_1226_296#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_18/a_735_102# hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_31/a_544_485#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_35/a_1034_424# hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_13/a_1141_508#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__a22o_1_7/a_230_79# hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_3/a_27_74#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_46/a_1178_124# hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_8/a_1141_508#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfrtp_4_1/a_1678_395# hr_16t4_mux_top_1/sky130_fd_sc_hs__a22o_1_5/a_222_392#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_37/a_206_368# hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_23/a_544_485#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_29/a_651_503# hr_16t4_mux_top_1/sky130_fd_sc_hs__a22o_1_7/B2
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__a22o_1_19/a_222_392# hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_33/a_1034_424#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfrtp_4_1/a_834_355# hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_35/a_27_74#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_7/a_544_485# hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_45/a_1178_124#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_7/a_1141_508# hr_16t4_mux_top_1/sky130_fd_sc_hs__dfrtp_4_1/a_812_138#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_1/a_1226_296# hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_37/a_437_503#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__clkbuf_2_3/a_43_192# hr_16t4_mux_top_1/sky130_fd_sc_hs__a22o_1_7/a_52_123#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfrtp_4_3/a_1350_392# hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_19/a_206_368#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_29/a_1141_508# hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_25/a_1226_296#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_41/a_1178_124# hr_16t4_mux_top_1/sky130_fd_sc_hs__a22o_1_15/a_132_392#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_19/a_437_503# hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_46/a_27_74#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_39/a_651_503# hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_31/a_1034_424#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_24/a_1226_296# hr_16t4_mux_top_1/sky130_fd_sc_hs__dfrtp_4_1/a_1350_392#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_5/a_1141_508# hr_16t4_mux_top_1/sky130_fd_sc_hs__a22o_1_3/a_222_392#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__clkbuf_16_1/a_114_74# hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_47/a_735_102#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__a22o_1_17/a_222_392# hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_23/a_1226_296#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_5/a_651_503# hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_27/a_206_368#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_37/a_27_74# hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_29/a_696_458#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_35/a_735_102# hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_27/a_1141_508#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_3/a_206_368# hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_39/a_1226_296#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__buf_2_1/a_21_260# hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_3/a_1141_508#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_18/a_206_368# hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_27/a_437_503#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__clkbuf_2_21/a_43_192# hr_16t4_mux_top_1/sky130_fd_sc_hs__a22o_1_1/a_132_392#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_3/a_437_503# hr_16t4_mux_top_1/sky130_fd_sc_hs__dfrtp_4_1/a_124_78#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_37/a_1226_296# hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_24/a_27_74#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_1/a_735_102# hr_16t4_mux_top_1/sky130_fd_sc_hs__buf_2_5/a_21_260#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__a22o_1_14/a_132_392# hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_37/a_651_503#
+ hr_16t4_mux_top_1/sky130_fd_sc_hs__dfxtp_4_18/a_437_503# hr_16t4_mux_top_1/sky130_fd_sc_hs__dfrtp_4_3/a_1647_81#
+ hr_16t4_mux_top
Xsky130_fd_sc_hs__clkinv_8_7 DVSS: DVDD: DVDD: DVSS: hr_16t4_mux_top_1/din[5] hr_16t4_mux_top_3/din[5]
+ sky130_fd_sc_hs__clkinv_8
Xsky130_fd_sc_hs__nand2_2_0 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__nand2_2_1/Y sky130_fd_sc_hs__nand2_2_1/B
+ sky130_fd_sc_hs__nand2_2_1/A sky130_fd_sc_hs__nand2_2_1/a_27_74# sky130_fd_sc_hs__nand2_2
Xsky130_fd_sc_hs__clkbuf_4_1 DVSS: DVDD: DVDD: DVSS: pi3_con[3] sky130_fd_sc_hs__clkbuf_4_1/X
+ sky130_fd_sc_hs__clkbuf_4_1/a_83_270# sky130_fd_sc_hs__clkbuf_4
Xsky130_fd_sc_hs__clkinv_4_1 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__nand2_2_27/B
+ sky130_fd_sc_hs__dlrtp_1_24/D sky130_fd_sc_hs__clkinv_4
Xsky130_fd_sc_hs__dlrtp_1_100 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__dlrtp_1_98/Q
+ sky130_fd_sc_hs__dlrtp_1_9/GATE sky130_fd_sc_hs__conb_1_95/HI sky130_fd_sc_hs__dlrtp_1_98/D
+ sky130_fd_sc_hs__dlrtp_1_98/a_216_424# sky130_fd_sc_hs__dlrtp_1_98/a_759_508# sky130_fd_sc_hs__dlrtp_1_98/a_565_74#
+ sky130_fd_sc_hs__dlrtp_1_98/a_27_424# sky130_fd_sc_hs__dlrtp_1_98/a_1045_74# sky130_fd_sc_hs__dlrtp_1_98/a_643_74#
+ sky130_fd_sc_hs__dlrtp_1_98/a_817_48# sky130_fd_sc_hs__dlrtp_1_98/a_568_392# sky130_fd_sc_hs__dlrtp_1_98/a_363_74#
+ sky130_fd_sc_hs__dlrtp_1_98/a_769_74# sky130_fd_sc_hs__dlrtp_1
Xsky130_fd_sc_hs__dlrtp_1_111 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__dlrtp_1_111/Q
+ sky130_fd_sc_hs__dlrtp_1_9/GATE sky130_fd_sc_hs__conb_1_131/HI sky130_fd_sc_hs__o21ai_2_39/Y
+ sky130_fd_sc_hs__dlrtp_1_111/a_216_424# sky130_fd_sc_hs__dlrtp_1_111/a_759_508#
+ sky130_fd_sc_hs__dlrtp_1_111/a_565_74# sky130_fd_sc_hs__dlrtp_1_111/a_27_424# sky130_fd_sc_hs__dlrtp_1_111/a_1045_74#
+ sky130_fd_sc_hs__dlrtp_1_111/a_643_74# sky130_fd_sc_hs__dlrtp_1_111/a_817_48# sky130_fd_sc_hs__dlrtp_1_111/a_568_392#
+ sky130_fd_sc_hs__dlrtp_1_111/a_363_74# sky130_fd_sc_hs__dlrtp_1_111/a_769_74# sky130_fd_sc_hs__dlrtp_1
Xsky130_fd_sc_hs__dlrtp_1_122 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__dlrtp_1_123/Q
+ sky130_fd_sc_hs__dlrtp_1_9/GATE sky130_fd_sc_hs__conb_1_131/HI sky130_fd_sc_hs__o21bai_2_49/Y
+ sky130_fd_sc_hs__dlrtp_1_123/a_216_424# sky130_fd_sc_hs__dlrtp_1_123/a_759_508#
+ sky130_fd_sc_hs__dlrtp_1_123/a_565_74# sky130_fd_sc_hs__dlrtp_1_123/a_27_424# sky130_fd_sc_hs__dlrtp_1_123/a_1045_74#
+ sky130_fd_sc_hs__dlrtp_1_123/a_643_74# sky130_fd_sc_hs__dlrtp_1_123/a_817_48# sky130_fd_sc_hs__dlrtp_1_123/a_568_392#
+ sky130_fd_sc_hs__dlrtp_1_123/a_363_74# sky130_fd_sc_hs__dlrtp_1_123/a_769_74# sky130_fd_sc_hs__dlrtp_1
Xsky130_fd_sc_hs__dlrtp_1_133 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__dlrtp_1_133/Q
+ sky130_fd_sc_hs__clkbuf_2_3/A sky130_fd_sc_hs__conb_1_135/HI sky130_fd_sc_hs__dlrtp_1_133/D
+ sky130_fd_sc_hs__dlrtp_1_133/a_216_424# sky130_fd_sc_hs__dlrtp_1_133/a_759_508#
+ sky130_fd_sc_hs__dlrtp_1_133/a_565_74# sky130_fd_sc_hs__dlrtp_1_133/a_27_424# sky130_fd_sc_hs__dlrtp_1_133/a_1045_74#
+ sky130_fd_sc_hs__dlrtp_1_133/a_643_74# sky130_fd_sc_hs__dlrtp_1_133/a_817_48# sky130_fd_sc_hs__dlrtp_1_133/a_568_392#
+ sky130_fd_sc_hs__dlrtp_1_133/a_363_74# sky130_fd_sc_hs__dlrtp_1_133/a_769_74# sky130_fd_sc_hs__dlrtp_1
Xsky130_fd_sc_hs__dlrtp_1_144 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__buf_2_35/A
+ sky130_fd_sc_hs__clkbuf_16_53/X sky130_fd_sc_hs__conb_1_127/HI sky130_fd_sc_hs__buf_2_153/X
+ sky130_fd_sc_hs__dlrtp_1_145/a_216_424# sky130_fd_sc_hs__dlrtp_1_145/a_759_508#
+ sky130_fd_sc_hs__dlrtp_1_145/a_565_74# sky130_fd_sc_hs__dlrtp_1_145/a_27_424# sky130_fd_sc_hs__dlrtp_1_145/a_1045_74#
+ sky130_fd_sc_hs__dlrtp_1_145/a_643_74# sky130_fd_sc_hs__dlrtp_1_145/a_817_48# sky130_fd_sc_hs__dlrtp_1_145/a_568_392#
+ sky130_fd_sc_hs__dlrtp_1_145/a_363_74# sky130_fd_sc_hs__dlrtp_1_145/a_769_74# sky130_fd_sc_hs__dlrtp_1
Xsky130_fd_sc_hs__dlrtp_1_155 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__dlrtp_1_157/Q
+ sky130_fd_sc_hs__clkbuf_16_53/X sky130_fd_sc_hs__conb_1_137/HI sky130_fd_sc_hs__dlrtp_1_157/D
+ sky130_fd_sc_hs__dlrtp_1_157/a_216_424# sky130_fd_sc_hs__dlrtp_1_157/a_759_508#
+ sky130_fd_sc_hs__dlrtp_1_157/a_565_74# sky130_fd_sc_hs__dlrtp_1_157/a_27_424# sky130_fd_sc_hs__dlrtp_1_157/a_1045_74#
+ sky130_fd_sc_hs__dlrtp_1_157/a_643_74# sky130_fd_sc_hs__dlrtp_1_157/a_817_48# sky130_fd_sc_hs__dlrtp_1_157/a_568_392#
+ sky130_fd_sc_hs__dlrtp_1_157/a_363_74# sky130_fd_sc_hs__dlrtp_1_157/a_769_74# sky130_fd_sc_hs__dlrtp_1
Xsky130_fd_sc_hs__inv_4_3 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__inv_4_3/Y ref_clk_ext_n
+ sky130_fd_sc_hs__inv_4
Xsky130_fd_sc_hs__dlrtp_1_90 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__dlrtp_1_91/Q
+ sky130_fd_sc_hs__dlrtp_1_9/GATE sky130_fd_sc_hs__conb_1_95/HI sky130_fd_sc_hs__buf_2_105/X
+ sky130_fd_sc_hs__dlrtp_1_91/a_216_424# sky130_fd_sc_hs__dlrtp_1_91/a_759_508# sky130_fd_sc_hs__dlrtp_1_91/a_565_74#
+ sky130_fd_sc_hs__dlrtp_1_91/a_27_424# sky130_fd_sc_hs__dlrtp_1_91/a_1045_74# sky130_fd_sc_hs__dlrtp_1_91/a_643_74#
+ sky130_fd_sc_hs__dlrtp_1_91/a_817_48# sky130_fd_sc_hs__dlrtp_1_91/a_568_392# sky130_fd_sc_hs__dlrtp_1_91/a_363_74#
+ sky130_fd_sc_hs__dlrtp_1_91/a_769_74# sky130_fd_sc_hs__dlrtp_1
Xsky130_fd_sc_hs__clkbuf_2_20 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__dlrtp_1_87/D
+ sky130_fd_sc_hs__o21ai_2_19/Y sky130_fd_sc_hs__clkbuf_2_21/a_43_192# sky130_fd_sc_hs__clkbuf_2
Xsky130_fd_sc_hs__clkbuf_2_31 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__einvp_2_3/TE
+ sky130_fd_sc_hs__dlrtp_1_91/Q sky130_fd_sc_hs__clkbuf_2_31/a_43_192# sky130_fd_sc_hs__clkbuf_2
Xsky130_fd_sc_hs__clkbuf_2_42 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__o21ai_2_31/A2
+ sky130_fd_sc_hs__or2b_4_1/X sky130_fd_sc_hs__clkbuf_2_43/a_43_192# sky130_fd_sc_hs__clkbuf_2
Xsky130_fd_sc_hs__clkbuf_2_53 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__dlrtp_1_29/D
+ sky130_fd_sc_hs__o21bai_2_53/Y sky130_fd_sc_hs__clkbuf_2_53/a_43_192# sky130_fd_sc_hs__clkbuf_2
Xsky130_fd_sc_hs__clkbuf_2_64 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__dlrtp_1_139/D
+ sky130_fd_sc_hs__o21bai_2_61/Y sky130_fd_sc_hs__clkbuf_2_65/a_43_192# sky130_fd_sc_hs__clkbuf_2
Xsky130_fd_sc_hs__buf_2_0 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__buf_2_3/X sky130_fd_sc_hs__inv_4_1/A
+ sky130_fd_sc_hs__buf_2_1/a_21_260# sky130_fd_sc_hs__buf_2
Xsky130_fd_sc_hs__dlrtp_1_2 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__dlrtp_1_3/Q sky130_fd_sc_hs__dlrtp_1_9/GATE
+ sky130_fd_sc_hs__conb_1_117/HI sky130_fd_sc_hs__buf_2_85/X sky130_fd_sc_hs__dlrtp_1_3/a_216_424#
+ sky130_fd_sc_hs__dlrtp_1_3/a_759_508# sky130_fd_sc_hs__dlrtp_1_3/a_565_74# sky130_fd_sc_hs__dlrtp_1_3/a_27_424#
+ sky130_fd_sc_hs__dlrtp_1_3/a_1045_74# sky130_fd_sc_hs__dlrtp_1_3/a_643_74# sky130_fd_sc_hs__dlrtp_1_3/a_817_48#
+ sky130_fd_sc_hs__dlrtp_1_3/a_568_392# sky130_fd_sc_hs__dlrtp_1_3/a_363_74# sky130_fd_sc_hs__dlrtp_1_3/a_769_74#
+ sky130_fd_sc_hs__dlrtp_1
Xsky130_fd_sc_hs__buf_2_60 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__buf_2_61/A sky130_fd_sc_hs__buf_2_61/X
+ sky130_fd_sc_hs__buf_2_61/a_21_260# sky130_fd_sc_hs__buf_2
Xsky130_fd_sc_hs__buf_2_71 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__buf_2_71/A sky130_fd_sc_hs__buf_2_71/X
+ sky130_fd_sc_hs__buf_2_71/a_21_260# sky130_fd_sc_hs__buf_2
Xsky130_fd_sc_hs__buf_2_82 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__buf_2_83/A sky130_fd_sc_hs__buf_2_83/X
+ sky130_fd_sc_hs__buf_2_83/a_21_260# sky130_fd_sc_hs__buf_2
Xsky130_fd_sc_hs__buf_2_93 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__buf_2_93/A sky130_fd_sc_hs__buf_2_93/X
+ sky130_fd_sc_hs__buf_2_93/a_21_260# sky130_fd_sc_hs__buf_2
Xsky130_fd_sc_hs__o21bai_2_40 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__o21ai_4_1/A1
+ sky130_fd_sc_hs__nand2_8_1/Y sky130_fd_sc_hs__dlrtp_1_21/D sky130_fd_sc_hs__o21bai_2_41/Y
+ sky130_fd_sc_hs__o21bai_2_41/a_27_74# sky130_fd_sc_hs__o21bai_2_41/a_225_74# sky130_fd_sc_hs__o21bai_2_41/a_507_368#
+ sky130_fd_sc_hs__o21bai_2
Xsky130_fd_sc_hs__o21bai_2_51 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__clkinv_4_5/Y
+ sky130_fd_sc_hs__nand2_2_21/B sky130_fd_sc_hs__dlrtp_1_29/D sky130_fd_sc_hs__buf_2_127/A
+ sky130_fd_sc_hs__o21bai_2_51/a_27_74# sky130_fd_sc_hs__o21bai_2_51/a_225_74# sky130_fd_sc_hs__o21bai_2_51/a_507_368#
+ sky130_fd_sc_hs__o21bai_2
Xsky130_fd_sc_hs__o21bai_2_62 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__o21bai_2_5/A1
+ sky130_fd_sc_hs__nand2_2_5/B sky130_fd_sc_hs__buf_2_153/X sky130_fd_sc_hs__buf_2_147/A
+ sky130_fd_sc_hs__o21bai_2_63/a_27_74# sky130_fd_sc_hs__o21bai_2_63/a_225_74# sky130_fd_sc_hs__o21bai_2_63/a_507_368#
+ sky130_fd_sc_hs__o21bai_2
Xsky130_fd_sc_hs__conb_1_260 DVSS: DVDD: DVDD: DVSS: prbs_generator_syn_31/eqn[31]
+ prbs_generator_syn_31/cke sky130_fd_sc_hs__conb_1_261/a_165_290# sky130_fd_sc_hs__conb_1_261/a_21_290#
+ sky130_fd_sc_hs__conb_1
Xsky130_fd_sc_hs__conb_1_271 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__conb_1_271/LO
+ sky130_fd_sc_hs__conb_1_271/HI sky130_fd_sc_hs__conb_1_271/a_165_290# sky130_fd_sc_hs__conb_1_271/a_21_290#
+ sky130_fd_sc_hs__conb_1
Xsky130_fd_sc_hs__clkbuf_8_30 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__clkbuf_8_31/X
+ sky130_fd_sc_hs__clkbuf_8_31/A sky130_fd_sc_hs__clkbuf_8_31/a_125_368# sky130_fd_sc_hs__clkbuf_8
Xsky130_fd_sc_hs__clkbuf_8_41 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__or2b_4_1/A
+ sky130_fd_sc_hs__nand2_2_23/Y sky130_fd_sc_hs__clkbuf_8_41/a_125_368# sky130_fd_sc_hs__clkbuf_8
Xsky130_fd_sc_hs__clkbuf_8_52 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__o21bai_4_7/A1
+ sky130_fd_sc_hs__nand2_2_31/Y sky130_fd_sc_hs__clkbuf_8_53/a_125_368# sky130_fd_sc_hs__clkbuf_8
Xsky130_fd_sc_hs__clkbuf_8_63 DVSS: DVDD: DVDD: DVSS: osc_core_1/con_perb_5[2] con_perb[2]
+ sky130_fd_sc_hs__clkbuf_8_63/a_125_368# sky130_fd_sc_hs__clkbuf_8
Xsky130_fd_sc_hs__clkbuf_8_74 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__clkbuf_8_75/X
+ sky130_fd_sc_hs__clkbuf_8_75/A sky130_fd_sc_hs__clkbuf_8_75/a_125_368# sky130_fd_sc_hs__clkbuf_8
Xsky130_fd_sc_hs__clkbuf_8_85 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__einvp_8_11/TE
+ test_mux_select[1] sky130_fd_sc_hs__clkbuf_8_85/a_125_368# sky130_fd_sc_hs__clkbuf_8
Xsky130_fd_sc_hs__clkbuf_8_96 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__clkbuf_8_97/X
+ CTL_BUF_N[1] sky130_fd_sc_hs__clkbuf_8_97/a_125_368# sky130_fd_sc_hs__clkbuf_8
Xsky130_fd_sc_hs__nor2_4_0 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__nor2_4_1/Y sky130_fd_sc_hs__nor2_4_1/A
+ sky130_fd_sc_hs__nor2_4_1/B sky130_fd_sc_hs__nor2_4_1/a_27_368# sky130_fd_sc_hs__nor2_4
Xsky130_fd_sc_hs__einvp_8_5 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__inv_4_39/A sky130_fd_sc_hs__einvp_8_5/TE
+ sky130_fd_sc_hs__einvp_8_5/A sky130_fd_sc_hs__einvp_8_5/a_802_323# sky130_fd_sc_hs__einvp_8_5/a_27_74#
+ sky130_fd_sc_hs__einvp_8_5/a_27_368# sky130_fd_sc_hs__einvp_8
Xsky130_fd_sc_hs__clkbuf_8_8 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__clkbuf_8_9/X
+ sky130_fd_sc_hs__clkbuf_8_9/A sky130_fd_sc_hs__clkbuf_8_9/a_125_368# sky130_fd_sc_hs__clkbuf_8
Xhr_16t4_mux_top_2 hr_16t4_mux_top_3/clk hr_16t4_mux_top_3/din[15] hr_16t4_mux_top_3/din[14]
+ hr_16t4_mux_top_3/din[13] hr_16t4_mux_top_3/din[12] hr_16t4_mux_top_3/din[11] hr_16t4_mux_top_3/din[10]
+ hr_16t4_mux_top_3/din[9] hr_16t4_mux_top_3/din[8] hr_16t4_mux_top_3/din[7] hr_16t4_mux_top_3/din[6]
+ hr_16t4_mux_top_3/din[5] hr_16t4_mux_top_3/din[4] hr_16t4_mux_top_3/din[3] hr_16t4_mux_top_3/din[2]
+ hr_16t4_mux_top_3/din[1] hr_16t4_mux_top_3/din[0] qr_4t1_mux_top_3/rst hr_16t4_mux_top_3/clk_prbs
+ qr_4t1_mux_top_3/din[3] qr_4t1_mux_top_3/din[2] qr_4t1_mux_top_3/din[1] qr_4t1_mux_top_3/din[0]
+ DVSS: DVDD: hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_31/D hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_15/a_735_102#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_23/Q hr_16t4_mux_top_3/sky130_fd_sc_hs__clkbuf_4_1/X
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__inv_4_11/A hr_16t4_mux_top_3/sky130_fd_sc_hs__clkbuf_2_25/a_43_192#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__inv_4_19/A hr_16t4_mux_top_3/sky130_fd_sc_hs__dfrtp_4_3/a_890_138#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__buf_2_11/a_21_260# hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_1/a_1141_508#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_5/Q hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_29/a_544_485#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_39/a_696_458# hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_46/a_735_102#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_47/a_1034_424# hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_24/D
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__a22o_1_9/A2 hr_16t4_mux_top_3/sky130_fd_sc_hs__a22o_1_9/B1
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_8/a_27_74# hr_16t4_mux_top_3/sky130_fd_sc_hs__a22o_1_5/X
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_19/a_651_503# hr_16t4_mux_top_3/sky130_fd_sc_hs__a22o_1_7/X
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_33/a_735_102# hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_31/a_27_74#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_46/a_1034_424# hr_16t4_mux_top_3/sky130_fd_sc_hs__clkinv_4_1/Y
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_25/a_1141_508# hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_46/Q
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_46/D hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_35/a_1226_296#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_5/a_696_458# hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_41/Q
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_45/a_1034_424# hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_24/a_1141_508#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__clkbuf_2_11/a_43_192# hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_33/a_1226_296#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__a22o_1_15/a_230_79# hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_47/a_206_368#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_39/a_544_485# hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_13/a_735_102#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_33/Q hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_23/a_1141_508#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__clkbuf_2_15/a_43_192# hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_45/D
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_29/Q hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_35/a_206_368#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_47/a_437_503# hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_27/a_651_503#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__inv_4_1/Y hr_16t4_mux_top_3/sky130_fd_sc_hs__a22o_1_17/X
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_45/a_735_102# hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_37/a_696_458#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_41/a_1034_424# hr_16t4_mux_top_3/sky130_fd_sc_hs__a22o_1_15/a_222_392#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_39/a_1141_508# hr_16t4_mux_top_3/sky130_fd_sc_hs__a22o_1_15/a_52_123#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_3/a_651_503# hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_15/D
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_5/a_544_485# hr_16t4_mux_top_3/sky130_fd_sc_hs__clkbuf_2_19/a_43_192#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_19/a_1178_124# hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_35/a_437_503#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_18/a_651_503# hr_16t4_mux_top_3/sky130_fd_sc_hs__inv_4_5/Y
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_37/a_1141_508# hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_31/a_1226_296#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_47/D hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_1/a_206_368#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_33/a_27_74# hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_18/a_1178_124#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_15/a_206_368# hr_16t4_mux_top_3/sky130_fd_sc_hs__a22o_1_23/a_132_392#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_5/D hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_19/a_696_458#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfrtp_4_3/a_313_74# hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_25/a_735_102#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__buf_2_5/X hr_16t4_mux_top_3/sky130_fd_sc_hs__a22o_1_5/B2
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_35/Q hr_16t4_mux_top_3/sky130_fd_sc_hs__dfrtp_4_3/a_494_366#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_1/a_437_503# hr_16t4_mux_top_3/sky130_fd_sc_hs__clkbuf_4_3/a_83_270#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__clkbuf_2_9/a_43_192# hr_16t4_mux_top_3/sky130_fd_sc_hs__a22o_1_19/X
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_9/a_735_102# hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_15/a_437_503#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_46/a_206_368# hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_37/a_544_485#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfrtp_4_1/a_1647_81# hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_8/Q
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfrtp_4_1/a_890_138# hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_15/a_1178_124#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__a22o_1_21/a_230_79# hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_33/a_206_368#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__a22o_1_1/a_222_392# hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_46/a_437_503#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__clkinv_2_1/Y hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_45/a_27_74#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__a22o_1_14/a_222_392# hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_35/a_1141_508#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_9/a_1178_124# hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_13/a_1178_124#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_33/a_437_503# hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_19/a_544_485#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_27/D hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_27/a_696_458#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_33/a_1141_508# hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_8/a_1178_124#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_5/a_27_74# hr_16t4_mux_top_3/sky130_fd_sc_hs__buf_2_15/X
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__inv_4_11/Y hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_18/Q
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_3/a_696_458# hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_13/a_206_368#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__a22o_1_21/a_52_123# hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_47/a_651_503#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_3/D hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_18/a_696_458#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_24/a_735_102# hr_16t4_mux_top_3/sky130_fd_sc_hs__clkbuf_2_23/a_43_192#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_7/a_1178_124# hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_47/a_1226_296#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__a22o_1_9/a_132_392# hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_8/a_735_102#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_45/a_206_368# hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_13/a_437_503#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_35/a_651_503# hr_16t4_mux_top_3/sky130_fd_sc_hs__dfrtp_4_3/a_2010_409#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_46/a_1226_296# hr_16t4_mux_top_3/sky130_fd_sc_hs__a22o_1_1/a_230_79#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_45/Q hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_23/a_27_74#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__a22o_1_11/a_230_79# hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_29/a_1178_124#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_45/a_437_503# hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_27/a_544_485#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_37/Q hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_41/a_735_102#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_31/a_1141_508# hr_16t4_mux_top_3/sky130_fd_sc_hs__inv_4_9/Y
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_45/a_1226_296# hr_16t4_mux_top_3/sky130_fd_sc_hs__dfrtp_4_1/a_37_78#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_1/a_651_503# hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_3/a_544_485#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__a22o_1_1/X hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_25/a_206_368#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__a22o_1_5/a_230_79# hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_15/a_651_503#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_18/a_544_485# hr_16t4_mux_top_3/sky130_fd_sc_hs__a22o_1_14/a_230_79#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfrtp_4_1/a_2010_409# hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_31/a_735_102#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__a22o_1_23/X hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_5/a_1178_124#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__buf_2_11/X hr_16t4_mux_top_3/sky130_fd_sc_hs__inv_4_19/Y
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_9/a_206_368# hr_16t4_mux_top_3/sky130_fd_sc_hs__a22o_1_1/a_52_123#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_15/a_27_74# hr_16t4_mux_top_3/sky130_fd_sc_hs__a22o_1_21/a_132_392#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_7/a_27_74# hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_1/D
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__a22o_1_11/a_52_123# hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_25/a_437_503#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_46/a_651_503# hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_23/a_735_102#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__a22o_1_9/a_230_79# hr_16t4_mux_top_3/sky130_fd_sc_hs__clkbuf_2_13/a_43_192#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_31/Q hr_16t4_mux_top_3/sky130_fd_sc_hs__a22o_1_19/a_230_79#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_41/a_1226_296# hr_16t4_mux_top_3/sky130_fd_sc_hs__dfrtp_4_1/a_494_366#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_19/a_1034_424# hr_16t4_mux_top_3/sky130_fd_sc_hs__a22o_1_21/X
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_9/a_437_503# hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_7/a_735_102#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_27/a_1178_124# hr_16t4_mux_top_3/sky130_fd_sc_hs__a22o_1_11/a_132_392#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__clkbuf_2_1/a_43_192# hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_33/a_651_503#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__a22o_1_5/a_52_123# hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_47/a_696_458#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__a22o_1_14/a_52_123# hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_3/a_1178_124#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__a22o_1_23/a_222_392# hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_39/D
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_18/a_1034_424# hr_16t4_mux_top_3/sky130_fd_sc_hs__clkbuf_2_17/a_43_192#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfrtp_4_1/Q hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_35/a_696_458#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__clkbuf_2_5/a_43_192# hr_16t4_mux_top_3/sky130_fd_sc_hs__inv_4_7/Y
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__a22o_1_9/a_52_123# hr_16t4_mux_top_3/sky130_fd_sc_hs__a22o_1_19/a_52_123#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfrtp_4_3/a_699_463# hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_24/a_206_368#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_13/a_651_503# hr_16t4_mux_top_3/sky130_fd_sc_hs__inv_4_21/Y
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_47/a_1141_508# hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_1/a_1178_124#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__inv_4_13/Y hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_15/a_1034_424#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_8/a_206_368# hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_1/a_696_458#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_19/Q hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_9/a_1034_424#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_24/a_437_503# hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_1/a_27_74#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_45/a_651_503# hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_47/a_544_485#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_15/a_696_458# hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_46/a_1141_508#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__buf_2_14/X hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_9/D
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_13/a_1034_424# hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_19/a_27_74#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__a22o_1_7/a_132_392# hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_8/a_437_503#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_27/Q hr_16t4_mux_top_3/sky130_fd_sc_hs__buf_2_9/X
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_25/a_1178_124# hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_8/a_1034_424#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_41/a_206_368# hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_35/a_544_485#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_46/a_696_458# hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_45/a_1141_508#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_24/a_1178_124# hr_16t4_mux_top_3/sky130_fd_sc_hs__a22o_1_9/a_222_392#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_7/a_1034_424# hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_31/a_206_368#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_25/a_651_503# hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_41/a_437_503#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_33/a_696_458# hr_16t4_mux_top_3/sky130_fd_sc_hs__buf_2_3/a_21_260#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_25/D hr_16t4_mux_top_3/sky130_fd_sc_hs__a22o_1_7/A2
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_9/a_651_503# hr_16t4_mux_top_3/sky130_fd_sc_hs__clkbuf_1_1/a_27_74#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_1/a_544_485# hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_23/a_1178_124#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_27/a_27_74# hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_23/a_206_368#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_31/a_437_503# hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_15/a_544_485#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_41/a_1141_508# hr_16t4_mux_top_3/sky130_fd_sc_hs__dfrtp_4_3/a_124_78#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_47/Q hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_29/a_1034_424#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__buf_2_7/a_21_260# hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_7/a_206_368#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_39/a_1178_124# hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_23/a_437_503#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_7/Q hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_46/a_544_485#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_13/a_696_458# hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_29/a_735_102#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__clkbuf_2_27/a_43_192# hr_16t4_mux_top_3/sky130_fd_sc_hs__a22o_1_3/X
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__buf_2_15/a_21_260# hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_7/a_437_503#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_37/a_1178_124# hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_5/a_1034_424#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_33/a_544_485# hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_45/a_696_458#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfrtp_4_3/a_1827_81# hr_16t4_mux_top_3/sky130_fd_sc_hs__a22o_1_21/a_222_392#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__a22o_1_3/a_230_79# hr_16t4_mux_top_3/sky130_fd_sc_hs__inv_4_17/Y
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_24/a_651_503# hr_16t4_mux_top_3/sky130_fd_sc_hs__inv_4_3/Y
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__a22o_1_11/a_222_392# hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_27/a_1034_424#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_19/a_1226_296# hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_8/a_651_503#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfrtp_4_1/a_699_463# hr_16t4_mux_top_3/sky130_fd_sc_hs__buf_2_7/X
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_3/a_1034_424# hr_16t4_mux_top_3/sky130_fd_sc_hs__a22o_1_17/a_230_79#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_13/a_544_485# hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_25/a_696_458#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_39/a_735_102# hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_29/a_27_74#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_18/a_1226_296# hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_9/a_696_458#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__a22o_1_3/a_52_123# hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_35/a_1178_124#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_47/a_27_74# hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_3/Q
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_41/a_651_503# hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_45/a_544_485#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_35/D hr_16t4_mux_top_3/sky130_fd_sc_hs__dfrtp_4_3/a_789_463#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__a22o_1_5/a_132_392# hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_33/a_1178_124#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_5/a_735_102# hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_1/a_1034_424#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__a22o_1_19/a_132_392# hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_13/a_27_74#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_31/a_651_503# hr_16t4_mux_top_3/sky130_fd_sc_hs__a22o_1_17/a_52_123#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfrtp_4_1/a_313_74# hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_23/D
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_15/a_1226_296# hr_16t4_mux_top_3/sky130_fd_sc_hs__clkbuf_2_31/a_43_192#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__inv_4_15/Y hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_39/a_27_74#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__a22o_1_7/a_222_392# hr_16t4_mux_top_3/sky130_fd_sc_hs__clkbuf_4_1/a_83_270#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_23/a_651_503# hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_25/a_544_485#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__clkbuf_2_7/a_43_192# hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_9/a_1226_296#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_8/D hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_25/a_1034_424#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfrtp_4_3/a_834_355# hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_13/a_1226_296#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_7/a_651_503# hr_16t4_mux_top_3/sky130_fd_sc_hs__dfrtp_4_3/a_1627_493#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_9/a_544_485# hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_29/a_206_368#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfrtp_4_3/a_812_138# hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_24/a_696_458#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_8/a_1226_296# hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_37/a_735_102#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_24/a_1034_424# hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_25/a_27_74#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_31/a_1178_124# hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_8/a_696_458#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_1/Q hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_29/a_437_503#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_7/a_1226_296# hr_16t4_mux_top_3/sky130_fd_sc_hs__dfrtp_4_3/a_37_78#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_23/a_1034_424# hr_16t4_mux_top_3/sky130_fd_sc_hs__a22o_1_23/a_230_79#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__a22o_1_3/a_132_392# hr_16t4_mux_top_3/sky130_fd_sc_hs__dfrtp_4_1/a_1627_493#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__a22o_1_17/a_132_392# hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_19/a_735_102#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_41/a_696_458# hr_16t4_mux_top_3/sky130_fd_sc_hs__dfrtp_4_1/a_1827_81#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_39/a_1034_424# hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_19/a_1141_508#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_9/a_27_74# hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_29/a_1226_296#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_18/a_27_74# hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_39/a_206_368#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_24/a_544_485# hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_31/a_696_458#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_37/a_1034_424# hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_18/a_1141_508#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_9/Q hr_16t4_mux_top_3/sky130_fd_sc_hs__a22o_1_23/a_52_123#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_8/a_544_485# hr_16t4_mux_top_3/sky130_fd_sc_hs__buf_2_3/X
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__buf_2_14/a_21_260# hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_5/a_1226_296#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_39/a_437_503# hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_23/a_696_458#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__buf_2_9/a_21_260# hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_5/a_206_368#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_7/a_696_458# hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_39/Q
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfrtp_4_3/a_1678_395# hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_41/a_544_485#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__clkbuf_2_29/a_43_192# hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_27/a_735_102#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfrtp_4_1/a_789_463# hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_15/a_1141_508#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__buf_2_1/X hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_41/a_27_74#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_5/a_437_503# hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_27/a_1226_296#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_3/a_735_102# hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_47/a_1178_124#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_9/a_1141_508# hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_3/a_1226_296#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_18/a_735_102# hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_31/a_544_485#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_35/a_1034_424# hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_13/a_1141_508#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__a22o_1_7/a_230_79# hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_3/a_27_74#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_46/a_1178_124# hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_8/a_1141_508#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfrtp_4_1/a_1678_395# hr_16t4_mux_top_3/sky130_fd_sc_hs__a22o_1_5/a_222_392#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_37/a_206_368# hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_23/a_544_485#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_29/a_651_503# hr_16t4_mux_top_3/sky130_fd_sc_hs__a22o_1_7/B2
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__a22o_1_19/a_222_392# hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_33/a_1034_424#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfrtp_4_1/a_834_355# hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_35/a_27_74#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_7/a_544_485# hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_45/a_1178_124#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_7/a_1141_508# hr_16t4_mux_top_3/sky130_fd_sc_hs__dfrtp_4_1/a_812_138#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_1/a_1226_296# hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_37/a_437_503#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__clkbuf_2_3/a_43_192# hr_16t4_mux_top_3/sky130_fd_sc_hs__a22o_1_7/a_52_123#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfrtp_4_3/a_1350_392# hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_19/a_206_368#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_29/a_1141_508# hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_25/a_1226_296#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_41/a_1178_124# hr_16t4_mux_top_3/sky130_fd_sc_hs__a22o_1_15/a_132_392#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_19/a_437_503# hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_46/a_27_74#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_39/a_651_503# hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_31/a_1034_424#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_24/a_1226_296# hr_16t4_mux_top_3/sky130_fd_sc_hs__dfrtp_4_1/a_1350_392#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_5/a_1141_508# hr_16t4_mux_top_3/sky130_fd_sc_hs__a22o_1_3/a_222_392#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__clkbuf_16_1/a_114_74# hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_47/a_735_102#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__a22o_1_17/a_222_392# hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_23/a_1226_296#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_5/a_651_503# hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_27/a_206_368#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_37/a_27_74# hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_29/a_696_458#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_35/a_735_102# hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_27/a_1141_508#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_3/a_206_368# hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_39/a_1226_296#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__buf_2_1/a_21_260# hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_3/a_1141_508#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_18/a_206_368# hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_27/a_437_503#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__clkbuf_2_21/a_43_192# hr_16t4_mux_top_3/sky130_fd_sc_hs__a22o_1_1/a_132_392#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_3/a_437_503# hr_16t4_mux_top_3/sky130_fd_sc_hs__dfrtp_4_1/a_124_78#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_37/a_1226_296# hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_24/a_27_74#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_1/a_735_102# hr_16t4_mux_top_3/sky130_fd_sc_hs__buf_2_5/a_21_260#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__a22o_1_14/a_132_392# hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_37/a_651_503#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_18/a_437_503# hr_16t4_mux_top_3/sky130_fd_sc_hs__dfrtp_4_3/a_1647_81#
+ hr_16t4_mux_top
Xsky130_fd_sc_hs__clkinv_8_8 DVSS: DVDD: DVDD: DVSS: prbs_generator_syn_1/out hr_16t4_mux_top_3/din[9]
+ sky130_fd_sc_hs__clkinv_8
Xsky130_fd_sc_hs__nand2_2_1 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__nand2_2_1/Y sky130_fd_sc_hs__nand2_2_1/B
+ sky130_fd_sc_hs__nand2_2_1/A sky130_fd_sc_hs__nand2_2_1/a_27_74# sky130_fd_sc_hs__nand2_2
Xsky130_fd_sc_hs__clkbuf_4_2 DVSS: DVDD: DVDD: DVSS: pi3_con[1] sky130_fd_sc_hs__clkbuf_8_9/A
+ sky130_fd_sc_hs__clkbuf_4_3/a_83_270# sky130_fd_sc_hs__clkbuf_4
Xsky130_fd_sc_hs__einvp_2_90 DVSS: DVDD: DVDD: DVSS: dout_p sky130_fd_sc_hs__einvp_2_99/A
+ sky130_fd_sc_hs__buf_2_63/X sky130_fd_sc_hs__einvp_2_91/a_263_323# sky130_fd_sc_hs__einvp_2_91/a_36_74#
+ sky130_fd_sc_hs__einvp_2_91/a_27_368# sky130_fd_sc_hs__einvp_2
Xsky130_fd_sc_hs__clkinv_4_2 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__clkinv_4_3/Y
+ sky130_fd_sc_hs__nor4_2_1/C sky130_fd_sc_hs__clkinv_4
Xsky130_fd_sc_hs__dlrtp_1_101 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__buf_2_99/A
+ sky130_fd_sc_hs__dlrtp_1_9/GATE sky130_fd_sc_hs__conb_1_131/HI sky130_fd_sc_hs__dlrtp_1_99/D
+ sky130_fd_sc_hs__dlrtp_1_99/a_216_424# sky130_fd_sc_hs__dlrtp_1_99/a_759_508# sky130_fd_sc_hs__dlrtp_1_99/a_565_74#
+ sky130_fd_sc_hs__dlrtp_1_99/a_27_424# sky130_fd_sc_hs__dlrtp_1_99/a_1045_74# sky130_fd_sc_hs__dlrtp_1_99/a_643_74#
+ sky130_fd_sc_hs__dlrtp_1_99/a_817_48# sky130_fd_sc_hs__dlrtp_1_99/a_568_392# sky130_fd_sc_hs__dlrtp_1_99/a_363_74#
+ sky130_fd_sc_hs__dlrtp_1_99/a_769_74# sky130_fd_sc_hs__dlrtp_1
Xsky130_fd_sc_hs__dlrtp_1_112 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__buf_2_123/A
+ sky130_fd_sc_hs__dlrtp_1_9/GATE sky130_fd_sc_hs__conb_1_131/HI sky130_fd_sc_hs__o21bai_2_43/Y
+ sky130_fd_sc_hs__dlrtp_1_113/a_216_424# sky130_fd_sc_hs__dlrtp_1_113/a_759_508#
+ sky130_fd_sc_hs__dlrtp_1_113/a_565_74# sky130_fd_sc_hs__dlrtp_1_113/a_27_424# sky130_fd_sc_hs__dlrtp_1_113/a_1045_74#
+ sky130_fd_sc_hs__dlrtp_1_113/a_643_74# sky130_fd_sc_hs__dlrtp_1_113/a_817_48# sky130_fd_sc_hs__dlrtp_1_113/a_568_392#
+ sky130_fd_sc_hs__dlrtp_1_113/a_363_74# sky130_fd_sc_hs__dlrtp_1_113/a_769_74# sky130_fd_sc_hs__dlrtp_1
Xsky130_fd_sc_hs__dlrtp_1_123 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__dlrtp_1_123/Q
+ sky130_fd_sc_hs__dlrtp_1_9/GATE sky130_fd_sc_hs__conb_1_131/HI sky130_fd_sc_hs__o21bai_2_49/Y
+ sky130_fd_sc_hs__dlrtp_1_123/a_216_424# sky130_fd_sc_hs__dlrtp_1_123/a_759_508#
+ sky130_fd_sc_hs__dlrtp_1_123/a_565_74# sky130_fd_sc_hs__dlrtp_1_123/a_27_424# sky130_fd_sc_hs__dlrtp_1_123/a_1045_74#
+ sky130_fd_sc_hs__dlrtp_1_123/a_643_74# sky130_fd_sc_hs__dlrtp_1_123/a_817_48# sky130_fd_sc_hs__dlrtp_1_123/a_568_392#
+ sky130_fd_sc_hs__dlrtp_1_123/a_363_74# sky130_fd_sc_hs__dlrtp_1_123/a_769_74# sky130_fd_sc_hs__dlrtp_1
Xsky130_fd_sc_hs__dlrtp_1_134 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__dlrtp_1_135/Q
+ sky130_fd_sc_hs__clkbuf_16_53/X sky130_fd_sc_hs__conb_1_135/HI sky130_fd_sc_hs__buf_2_141/X
+ sky130_fd_sc_hs__dlrtp_1_135/a_216_424# sky130_fd_sc_hs__dlrtp_1_135/a_759_508#
+ sky130_fd_sc_hs__dlrtp_1_135/a_565_74# sky130_fd_sc_hs__dlrtp_1_135/a_27_424# sky130_fd_sc_hs__dlrtp_1_135/a_1045_74#
+ sky130_fd_sc_hs__dlrtp_1_135/a_643_74# sky130_fd_sc_hs__dlrtp_1_135/a_817_48# sky130_fd_sc_hs__dlrtp_1_135/a_568_392#
+ sky130_fd_sc_hs__dlrtp_1_135/a_363_74# sky130_fd_sc_hs__dlrtp_1_135/a_769_74# sky130_fd_sc_hs__dlrtp_1
Xsky130_fd_sc_hs__dlrtp_1_145 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__buf_2_35/A
+ sky130_fd_sc_hs__clkbuf_16_53/X sky130_fd_sc_hs__conb_1_127/HI sky130_fd_sc_hs__buf_2_153/X
+ sky130_fd_sc_hs__dlrtp_1_145/a_216_424# sky130_fd_sc_hs__dlrtp_1_145/a_759_508#
+ sky130_fd_sc_hs__dlrtp_1_145/a_565_74# sky130_fd_sc_hs__dlrtp_1_145/a_27_424# sky130_fd_sc_hs__dlrtp_1_145/a_1045_74#
+ sky130_fd_sc_hs__dlrtp_1_145/a_643_74# sky130_fd_sc_hs__dlrtp_1_145/a_817_48# sky130_fd_sc_hs__dlrtp_1_145/a_568_392#
+ sky130_fd_sc_hs__dlrtp_1_145/a_363_74# sky130_fd_sc_hs__dlrtp_1_145/a_769_74# sky130_fd_sc_hs__dlrtp_1
Xsky130_fd_sc_hs__dlrtp_1_156 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__buf_2_155/A
+ sky130_fd_sc_hs__clkbuf_16_53/X sky130_fd_sc_hs__conb_1_137/HI sky130_fd_sc_hs__buf_2_163/X
+ sky130_fd_sc_hs__dlrtp_1_156/a_216_424# sky130_fd_sc_hs__dlrtp_1_156/a_759_508#
+ sky130_fd_sc_hs__dlrtp_1_156/a_565_74# sky130_fd_sc_hs__dlrtp_1_156/a_27_424# sky130_fd_sc_hs__dlrtp_1_156/a_1045_74#
+ sky130_fd_sc_hs__dlrtp_1_156/a_643_74# sky130_fd_sc_hs__dlrtp_1_156/a_817_48# sky130_fd_sc_hs__dlrtp_1_156/a_568_392#
+ sky130_fd_sc_hs__dlrtp_1_156/a_363_74# sky130_fd_sc_hs__dlrtp_1_156/a_769_74# sky130_fd_sc_hs__dlrtp_1
Xsky130_fd_sc_hs__inv_4_4 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__inv_4_5/Y ref_clk_ext_n
+ sky130_fd_sc_hs__inv_4
Xsky130_fd_sc_hs__dlrtp_1_80 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__dlrtp_1_81/Q
+ sky130_fd_sc_hs__clkbuf_16_53/X sky130_fd_sc_hs__conb_1_137/HI sky130_fd_sc_hs__buf_2_73/X
+ sky130_fd_sc_hs__dlrtp_1_81/a_216_424# sky130_fd_sc_hs__dlrtp_1_81/a_759_508# sky130_fd_sc_hs__dlrtp_1_81/a_565_74#
+ sky130_fd_sc_hs__dlrtp_1_81/a_27_424# sky130_fd_sc_hs__dlrtp_1_81/a_1045_74# sky130_fd_sc_hs__dlrtp_1_81/a_643_74#
+ sky130_fd_sc_hs__dlrtp_1_81/a_817_48# sky130_fd_sc_hs__dlrtp_1_81/a_568_392# sky130_fd_sc_hs__dlrtp_1_81/a_363_74#
+ sky130_fd_sc_hs__dlrtp_1_81/a_769_74# sky130_fd_sc_hs__dlrtp_1
Xsky130_fd_sc_hs__dlrtp_1_91 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__dlrtp_1_91/Q
+ sky130_fd_sc_hs__dlrtp_1_9/GATE sky130_fd_sc_hs__conb_1_95/HI sky130_fd_sc_hs__buf_2_105/X
+ sky130_fd_sc_hs__dlrtp_1_91/a_216_424# sky130_fd_sc_hs__dlrtp_1_91/a_759_508# sky130_fd_sc_hs__dlrtp_1_91/a_565_74#
+ sky130_fd_sc_hs__dlrtp_1_91/a_27_424# sky130_fd_sc_hs__dlrtp_1_91/a_1045_74# sky130_fd_sc_hs__dlrtp_1_91/a_643_74#
+ sky130_fd_sc_hs__dlrtp_1_91/a_817_48# sky130_fd_sc_hs__dlrtp_1_91/a_568_392# sky130_fd_sc_hs__dlrtp_1_91/a_363_74#
+ sky130_fd_sc_hs__dlrtp_1_91/a_769_74# sky130_fd_sc_hs__dlrtp_1
Xsky130_fd_sc_hs__clkbuf_2_10 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__dlrtp_1_55/D
+ sky130_fd_sc_hs__o21ai_2_11/Y sky130_fd_sc_hs__clkbuf_2_11/a_43_192# sky130_fd_sc_hs__clkbuf_2
Xsky130_fd_sc_hs__clkbuf_2_21 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__dlrtp_1_87/D
+ sky130_fd_sc_hs__o21ai_2_19/Y sky130_fd_sc_hs__clkbuf_2_21/a_43_192# sky130_fd_sc_hs__clkbuf_2
Xsky130_fd_sc_hs__clkbuf_2_32 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__dlrtp_1_9/D
+ sky130_fd_sc_hs__buf_2_95/X sky130_fd_sc_hs__clkbuf_2_33/a_43_192# sky130_fd_sc_hs__clkbuf_2
Xsky130_fd_sc_hs__clkbuf_2_43 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__o21ai_2_31/A2
+ sky130_fd_sc_hs__or2b_4_1/X sky130_fd_sc_hs__clkbuf_2_43/a_43_192# sky130_fd_sc_hs__clkbuf_2
Xsky130_fd_sc_hs__clkbuf_2_54 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__dlrtp_1_121/D
+ sky130_fd_sc_hs__o21ai_2_47/Y sky130_fd_sc_hs__clkbuf_2_55/a_43_192# sky130_fd_sc_hs__clkbuf_2
Xsky130_fd_sc_hs__clkbuf_2_65 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__dlrtp_1_139/D
+ sky130_fd_sc_hs__o21bai_2_61/Y sky130_fd_sc_hs__clkbuf_2_65/a_43_192# sky130_fd_sc_hs__clkbuf_2
Xsky130_fd_sc_hs__buf_2_1 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__buf_2_3/X sky130_fd_sc_hs__inv_4_1/A
+ sky130_fd_sc_hs__buf_2_1/a_21_260# sky130_fd_sc_hs__buf_2
Xsky130_fd_sc_hs__dlrtp_1_3 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__dlrtp_1_3/Q sky130_fd_sc_hs__dlrtp_1_9/GATE
+ sky130_fd_sc_hs__conb_1_117/HI sky130_fd_sc_hs__buf_2_85/X sky130_fd_sc_hs__dlrtp_1_3/a_216_424#
+ sky130_fd_sc_hs__dlrtp_1_3/a_759_508# sky130_fd_sc_hs__dlrtp_1_3/a_565_74# sky130_fd_sc_hs__dlrtp_1_3/a_27_424#
+ sky130_fd_sc_hs__dlrtp_1_3/a_1045_74# sky130_fd_sc_hs__dlrtp_1_3/a_643_74# sky130_fd_sc_hs__dlrtp_1_3/a_817_48#
+ sky130_fd_sc_hs__dlrtp_1_3/a_568_392# sky130_fd_sc_hs__dlrtp_1_3/a_363_74# sky130_fd_sc_hs__dlrtp_1_3/a_769_74#
+ sky130_fd_sc_hs__dlrtp_1
Xsky130_fd_sc_hs__buf_2_50 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__buf_2_51/A sky130_fd_sc_hs__buf_2_51/X
+ sky130_fd_sc_hs__buf_2_51/a_21_260# sky130_fd_sc_hs__buf_2
Xsky130_fd_sc_hs__buf_2_61 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__buf_2_61/A sky130_fd_sc_hs__buf_2_61/X
+ sky130_fd_sc_hs__buf_2_61/a_21_260# sky130_fd_sc_hs__buf_2
Xsky130_fd_sc_hs__buf_2_72 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__buf_2_79/X sky130_fd_sc_hs__buf_2_73/X
+ sky130_fd_sc_hs__buf_2_73/a_21_260# sky130_fd_sc_hs__buf_2
Xsky130_fd_sc_hs__buf_2_83 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__buf_2_83/A sky130_fd_sc_hs__buf_2_83/X
+ sky130_fd_sc_hs__buf_2_83/a_21_260# sky130_fd_sc_hs__buf_2
Xsky130_fd_sc_hs__buf_2_94 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__buf_2_95/A sky130_fd_sc_hs__buf_2_95/X
+ sky130_fd_sc_hs__buf_2_95/a_21_260# sky130_fd_sc_hs__buf_2
Xsky130_fd_sc_hs__o21bai_2_30 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__o21ai_4_1/A1
+ sky130_fd_sc_hs__o21bai_4_3/A2 sky130_fd_sc_hs__dlrtp_1_103/D sky130_fd_sc_hs__o21bai_2_31/Y
+ sky130_fd_sc_hs__o21bai_2_31/a_27_74# sky130_fd_sc_hs__o21bai_2_31/a_225_74# sky130_fd_sc_hs__o21bai_2_31/a_507_368#
+ sky130_fd_sc_hs__o21bai_2
Xsky130_fd_sc_hs__o21bai_2_41 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__o21ai_4_1/A1
+ sky130_fd_sc_hs__nand2_8_1/Y sky130_fd_sc_hs__dlrtp_1_21/D sky130_fd_sc_hs__o21bai_2_41/Y
+ sky130_fd_sc_hs__o21bai_2_41/a_27_74# sky130_fd_sc_hs__o21bai_2_41/a_225_74# sky130_fd_sc_hs__o21bai_2_41/a_507_368#
+ sky130_fd_sc_hs__o21bai_2
Xsky130_fd_sc_hs__o21bai_2_52 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__clkinv_4_3/Y
+ sky130_fd_sc_hs__nand2_2_21/B sky130_fd_sc_hs__dlrtp_1_121/D sky130_fd_sc_hs__o21bai_2_53/Y
+ sky130_fd_sc_hs__o21bai_2_53/a_27_74# sky130_fd_sc_hs__o21bai_2_53/a_225_74# sky130_fd_sc_hs__o21bai_2_53/a_507_368#
+ sky130_fd_sc_hs__o21bai_2
Xsky130_fd_sc_hs__o21bai_2_63 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__o21bai_2_5/A1
+ sky130_fd_sc_hs__nand2_2_5/B sky130_fd_sc_hs__buf_2_153/X sky130_fd_sc_hs__buf_2_147/A
+ sky130_fd_sc_hs__o21bai_2_63/a_27_74# sky130_fd_sc_hs__o21bai_2_63/a_225_74# sky130_fd_sc_hs__o21bai_2_63/a_507_368#
+ sky130_fd_sc_hs__o21bai_2
Xsky130_fd_sc_hs__conb_1_250 DVSS: DVDD: DVDD: DVSS: prbs_generator_syn_27/eqn[28]
+ sky130_fd_sc_hs__conb_1_251/HI sky130_fd_sc_hs__conb_1_251/a_165_290# sky130_fd_sc_hs__conb_1_251/a_21_290#
+ sky130_fd_sc_hs__conb_1
Xsky130_fd_sc_hs__conb_1_261 DVSS: DVDD: DVDD: DVSS: prbs_generator_syn_31/eqn[31]
+ prbs_generator_syn_31/cke sky130_fd_sc_hs__conb_1_261/a_165_290# sky130_fd_sc_hs__conb_1_261/a_21_290#
+ sky130_fd_sc_hs__conb_1
Xsky130_fd_sc_hs__conb_1_272 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__conb_1_273/LO
+ sky130_fd_sc_hs__conb_1_273/HI sky130_fd_sc_hs__conb_1_273/a_165_290# sky130_fd_sc_hs__conb_1_273/a_21_290#
+ sky130_fd_sc_hs__conb_1
Xsky130_fd_sc_hs__clkbuf_8_20 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__clkbuf_8_21/X
+ sky130_fd_sc_hs__clkbuf_8_21/A sky130_fd_sc_hs__clkbuf_8_21/a_125_368# sky130_fd_sc_hs__clkbuf_8
Xsky130_fd_sc_hs__clkbuf_8_31 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__clkbuf_8_31/X
+ sky130_fd_sc_hs__clkbuf_8_31/A sky130_fd_sc_hs__clkbuf_8_31/a_125_368# sky130_fd_sc_hs__clkbuf_8
Xsky130_fd_sc_hs__clkbuf_8_42 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__o21bai_4_3/A2
+ sky130_fd_sc_hs__nand2_2_25/Y sky130_fd_sc_hs__clkbuf_8_43/a_125_368# sky130_fd_sc_hs__clkbuf_8
Xsky130_fd_sc_hs__clkbuf_8_53 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__o21bai_4_7/A1
+ sky130_fd_sc_hs__nand2_2_31/Y sky130_fd_sc_hs__clkbuf_8_53/a_125_368# sky130_fd_sc_hs__clkbuf_8
Xsky130_fd_sc_hs__clkbuf_8_64 DVSS: DVDD: DVDD: DVSS: fine_freq_track_1/aux_osc_en
+ aux_osc_en sky130_fd_sc_hs__clkbuf_8_65/a_125_368# sky130_fd_sc_hs__clkbuf_8
Xsky130_fd_sc_hs__clkbuf_8_75 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__clkbuf_8_75/X
+ sky130_fd_sc_hs__clkbuf_8_75/A sky130_fd_sc_hs__clkbuf_8_75/a_125_368# sky130_fd_sc_hs__clkbuf_8
Xsky130_fd_sc_hs__clkbuf_8_86 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__einvp_8_5/TE
+ test_mux_select[2] sky130_fd_sc_hs__clkbuf_8_87/a_125_368# sky130_fd_sc_hs__clkbuf_8
Xsky130_fd_sc_hs__clkbuf_8_97 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__clkbuf_8_97/X
+ CTL_BUF_N[1] sky130_fd_sc_hs__clkbuf_8_97/a_125_368# sky130_fd_sc_hs__clkbuf_8
Xsky130_fd_sc_hs__nor2_4_1 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__nor2_4_1/Y sky130_fd_sc_hs__nor2_4_1/A
+ sky130_fd_sc_hs__nor2_4_1/B sky130_fd_sc_hs__nor2_4_1/a_27_368# sky130_fd_sc_hs__nor2_4
Xsky130_fd_sc_hs__einvp_8_6 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__inv_4_39/A sky130_fd_sc_hs__einvp_8_7/TE
+ osc_core_1/osc_hold sky130_fd_sc_hs__einvp_8_7/a_802_323# sky130_fd_sc_hs__einvp_8_7/a_27_74#
+ sky130_fd_sc_hs__einvp_8_7/a_27_368# sky130_fd_sc_hs__einvp_8
Xsky130_fd_sc_hs__clkbuf_8_9 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__clkbuf_8_9/X
+ sky130_fd_sc_hs__clkbuf_8_9/A sky130_fd_sc_hs__clkbuf_8_9/a_125_368# sky130_fd_sc_hs__clkbuf_8
Xhr_16t4_mux_top_3 hr_16t4_mux_top_3/clk hr_16t4_mux_top_3/din[15] hr_16t4_mux_top_3/din[14]
+ hr_16t4_mux_top_3/din[13] hr_16t4_mux_top_3/din[12] hr_16t4_mux_top_3/din[11] hr_16t4_mux_top_3/din[10]
+ hr_16t4_mux_top_3/din[9] hr_16t4_mux_top_3/din[8] hr_16t4_mux_top_3/din[7] hr_16t4_mux_top_3/din[6]
+ hr_16t4_mux_top_3/din[5] hr_16t4_mux_top_3/din[4] hr_16t4_mux_top_3/din[3] hr_16t4_mux_top_3/din[2]
+ hr_16t4_mux_top_3/din[1] hr_16t4_mux_top_3/din[0] qr_4t1_mux_top_3/rst hr_16t4_mux_top_3/clk_prbs
+ qr_4t1_mux_top_3/din[3] qr_4t1_mux_top_3/din[2] qr_4t1_mux_top_3/din[1] qr_4t1_mux_top_3/din[0]
+ DVSS: DVDD: hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_31/D hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_15/a_735_102#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_23/Q hr_16t4_mux_top_3/sky130_fd_sc_hs__clkbuf_4_1/X
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__inv_4_11/A hr_16t4_mux_top_3/sky130_fd_sc_hs__clkbuf_2_25/a_43_192#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__inv_4_19/A hr_16t4_mux_top_3/sky130_fd_sc_hs__dfrtp_4_3/a_890_138#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__buf_2_11/a_21_260# hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_1/a_1141_508#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_5/Q hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_29/a_544_485#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_39/a_696_458# hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_46/a_735_102#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_47/a_1034_424# hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_24/D
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__a22o_1_9/A2 hr_16t4_mux_top_3/sky130_fd_sc_hs__a22o_1_9/B1
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_8/a_27_74# hr_16t4_mux_top_3/sky130_fd_sc_hs__a22o_1_5/X
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_19/a_651_503# hr_16t4_mux_top_3/sky130_fd_sc_hs__a22o_1_7/X
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_33/a_735_102# hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_31/a_27_74#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_46/a_1034_424# hr_16t4_mux_top_3/sky130_fd_sc_hs__clkinv_4_1/Y
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_25/a_1141_508# hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_46/Q
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_46/D hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_35/a_1226_296#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_5/a_696_458# hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_41/Q
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_45/a_1034_424# hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_24/a_1141_508#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__clkbuf_2_11/a_43_192# hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_33/a_1226_296#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__a22o_1_15/a_230_79# hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_47/a_206_368#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_39/a_544_485# hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_13/a_735_102#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_33/Q hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_23/a_1141_508#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__clkbuf_2_15/a_43_192# hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_45/D
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_29/Q hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_35/a_206_368#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_47/a_437_503# hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_27/a_651_503#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__inv_4_1/Y hr_16t4_mux_top_3/sky130_fd_sc_hs__a22o_1_17/X
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_45/a_735_102# hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_37/a_696_458#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_41/a_1034_424# hr_16t4_mux_top_3/sky130_fd_sc_hs__a22o_1_15/a_222_392#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_39/a_1141_508# hr_16t4_mux_top_3/sky130_fd_sc_hs__a22o_1_15/a_52_123#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_3/a_651_503# hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_15/D
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_5/a_544_485# hr_16t4_mux_top_3/sky130_fd_sc_hs__clkbuf_2_19/a_43_192#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_19/a_1178_124# hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_35/a_437_503#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_18/a_651_503# hr_16t4_mux_top_3/sky130_fd_sc_hs__inv_4_5/Y
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_37/a_1141_508# hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_31/a_1226_296#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_47/D hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_1/a_206_368#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_33/a_27_74# hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_18/a_1178_124#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_15/a_206_368# hr_16t4_mux_top_3/sky130_fd_sc_hs__a22o_1_23/a_132_392#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_5/D hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_19/a_696_458#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfrtp_4_3/a_313_74# hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_25/a_735_102#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__buf_2_5/X hr_16t4_mux_top_3/sky130_fd_sc_hs__a22o_1_5/B2
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_35/Q hr_16t4_mux_top_3/sky130_fd_sc_hs__dfrtp_4_3/a_494_366#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_1/a_437_503# hr_16t4_mux_top_3/sky130_fd_sc_hs__clkbuf_4_3/a_83_270#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__clkbuf_2_9/a_43_192# hr_16t4_mux_top_3/sky130_fd_sc_hs__a22o_1_19/X
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_9/a_735_102# hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_15/a_437_503#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_46/a_206_368# hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_37/a_544_485#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfrtp_4_1/a_1647_81# hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_8/Q
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfrtp_4_1/a_890_138# hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_15/a_1178_124#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__a22o_1_21/a_230_79# hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_33/a_206_368#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__a22o_1_1/a_222_392# hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_46/a_437_503#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__clkinv_2_1/Y hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_45/a_27_74#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__a22o_1_14/a_222_392# hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_35/a_1141_508#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_9/a_1178_124# hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_13/a_1178_124#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_33/a_437_503# hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_19/a_544_485#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_27/D hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_27/a_696_458#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_33/a_1141_508# hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_8/a_1178_124#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_5/a_27_74# hr_16t4_mux_top_3/sky130_fd_sc_hs__buf_2_15/X
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__inv_4_11/Y hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_18/Q
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_3/a_696_458# hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_13/a_206_368#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__a22o_1_21/a_52_123# hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_47/a_651_503#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_3/D hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_18/a_696_458#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_24/a_735_102# hr_16t4_mux_top_3/sky130_fd_sc_hs__clkbuf_2_23/a_43_192#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_7/a_1178_124# hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_47/a_1226_296#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__a22o_1_9/a_132_392# hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_8/a_735_102#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_45/a_206_368# hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_13/a_437_503#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_35/a_651_503# hr_16t4_mux_top_3/sky130_fd_sc_hs__dfrtp_4_3/a_2010_409#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_46/a_1226_296# hr_16t4_mux_top_3/sky130_fd_sc_hs__a22o_1_1/a_230_79#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_45/Q hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_23/a_27_74#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__a22o_1_11/a_230_79# hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_29/a_1178_124#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_45/a_437_503# hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_27/a_544_485#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_37/Q hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_41/a_735_102#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_31/a_1141_508# hr_16t4_mux_top_3/sky130_fd_sc_hs__inv_4_9/Y
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_45/a_1226_296# hr_16t4_mux_top_3/sky130_fd_sc_hs__dfrtp_4_1/a_37_78#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_1/a_651_503# hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_3/a_544_485#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__a22o_1_1/X hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_25/a_206_368#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__a22o_1_5/a_230_79# hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_15/a_651_503#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_18/a_544_485# hr_16t4_mux_top_3/sky130_fd_sc_hs__a22o_1_14/a_230_79#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfrtp_4_1/a_2010_409# hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_31/a_735_102#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__a22o_1_23/X hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_5/a_1178_124#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__buf_2_11/X hr_16t4_mux_top_3/sky130_fd_sc_hs__inv_4_19/Y
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_9/a_206_368# hr_16t4_mux_top_3/sky130_fd_sc_hs__a22o_1_1/a_52_123#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_15/a_27_74# hr_16t4_mux_top_3/sky130_fd_sc_hs__a22o_1_21/a_132_392#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_7/a_27_74# hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_1/D
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__a22o_1_11/a_52_123# hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_25/a_437_503#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_46/a_651_503# hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_23/a_735_102#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__a22o_1_9/a_230_79# hr_16t4_mux_top_3/sky130_fd_sc_hs__clkbuf_2_13/a_43_192#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_31/Q hr_16t4_mux_top_3/sky130_fd_sc_hs__a22o_1_19/a_230_79#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_41/a_1226_296# hr_16t4_mux_top_3/sky130_fd_sc_hs__dfrtp_4_1/a_494_366#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_19/a_1034_424# hr_16t4_mux_top_3/sky130_fd_sc_hs__a22o_1_21/X
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_9/a_437_503# hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_7/a_735_102#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_27/a_1178_124# hr_16t4_mux_top_3/sky130_fd_sc_hs__a22o_1_11/a_132_392#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__clkbuf_2_1/a_43_192# hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_33/a_651_503#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__a22o_1_5/a_52_123# hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_47/a_696_458#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__a22o_1_14/a_52_123# hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_3/a_1178_124#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__a22o_1_23/a_222_392# hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_39/D
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_18/a_1034_424# hr_16t4_mux_top_3/sky130_fd_sc_hs__clkbuf_2_17/a_43_192#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfrtp_4_1/Q hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_35/a_696_458#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__clkbuf_2_5/a_43_192# hr_16t4_mux_top_3/sky130_fd_sc_hs__inv_4_7/Y
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__a22o_1_9/a_52_123# hr_16t4_mux_top_3/sky130_fd_sc_hs__a22o_1_19/a_52_123#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfrtp_4_3/a_699_463# hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_24/a_206_368#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_13/a_651_503# hr_16t4_mux_top_3/sky130_fd_sc_hs__inv_4_21/Y
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_47/a_1141_508# hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_1/a_1178_124#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__inv_4_13/Y hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_15/a_1034_424#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_8/a_206_368# hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_1/a_696_458#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_19/Q hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_9/a_1034_424#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_24/a_437_503# hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_1/a_27_74#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_45/a_651_503# hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_47/a_544_485#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_15/a_696_458# hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_46/a_1141_508#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__buf_2_14/X hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_9/D
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_13/a_1034_424# hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_19/a_27_74#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__a22o_1_7/a_132_392# hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_8/a_437_503#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_27/Q hr_16t4_mux_top_3/sky130_fd_sc_hs__buf_2_9/X
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_25/a_1178_124# hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_8/a_1034_424#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_41/a_206_368# hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_35/a_544_485#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_46/a_696_458# hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_45/a_1141_508#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_24/a_1178_124# hr_16t4_mux_top_3/sky130_fd_sc_hs__a22o_1_9/a_222_392#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_7/a_1034_424# hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_31/a_206_368#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_25/a_651_503# hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_41/a_437_503#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_33/a_696_458# hr_16t4_mux_top_3/sky130_fd_sc_hs__buf_2_3/a_21_260#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_25/D hr_16t4_mux_top_3/sky130_fd_sc_hs__a22o_1_7/A2
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_9/a_651_503# hr_16t4_mux_top_3/sky130_fd_sc_hs__clkbuf_1_1/a_27_74#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_1/a_544_485# hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_23/a_1178_124#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_27/a_27_74# hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_23/a_206_368#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_31/a_437_503# hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_15/a_544_485#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_41/a_1141_508# hr_16t4_mux_top_3/sky130_fd_sc_hs__dfrtp_4_3/a_124_78#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_47/Q hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_29/a_1034_424#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__buf_2_7/a_21_260# hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_7/a_206_368#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_39/a_1178_124# hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_23/a_437_503#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_7/Q hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_46/a_544_485#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_13/a_696_458# hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_29/a_735_102#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__clkbuf_2_27/a_43_192# hr_16t4_mux_top_3/sky130_fd_sc_hs__a22o_1_3/X
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__buf_2_15/a_21_260# hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_7/a_437_503#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_37/a_1178_124# hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_5/a_1034_424#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_33/a_544_485# hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_45/a_696_458#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfrtp_4_3/a_1827_81# hr_16t4_mux_top_3/sky130_fd_sc_hs__a22o_1_21/a_222_392#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__a22o_1_3/a_230_79# hr_16t4_mux_top_3/sky130_fd_sc_hs__inv_4_17/Y
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_24/a_651_503# hr_16t4_mux_top_3/sky130_fd_sc_hs__inv_4_3/Y
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__a22o_1_11/a_222_392# hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_27/a_1034_424#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_19/a_1226_296# hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_8/a_651_503#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfrtp_4_1/a_699_463# hr_16t4_mux_top_3/sky130_fd_sc_hs__buf_2_7/X
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_3/a_1034_424# hr_16t4_mux_top_3/sky130_fd_sc_hs__a22o_1_17/a_230_79#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_13/a_544_485# hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_25/a_696_458#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_39/a_735_102# hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_29/a_27_74#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_18/a_1226_296# hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_9/a_696_458#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__a22o_1_3/a_52_123# hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_35/a_1178_124#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_47/a_27_74# hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_3/Q
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_41/a_651_503# hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_45/a_544_485#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_35/D hr_16t4_mux_top_3/sky130_fd_sc_hs__dfrtp_4_3/a_789_463#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__a22o_1_5/a_132_392# hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_33/a_1178_124#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_5/a_735_102# hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_1/a_1034_424#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__a22o_1_19/a_132_392# hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_13/a_27_74#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_31/a_651_503# hr_16t4_mux_top_3/sky130_fd_sc_hs__a22o_1_17/a_52_123#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfrtp_4_1/a_313_74# hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_23/D
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_15/a_1226_296# hr_16t4_mux_top_3/sky130_fd_sc_hs__clkbuf_2_31/a_43_192#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__inv_4_15/Y hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_39/a_27_74#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__a22o_1_7/a_222_392# hr_16t4_mux_top_3/sky130_fd_sc_hs__clkbuf_4_1/a_83_270#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_23/a_651_503# hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_25/a_544_485#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__clkbuf_2_7/a_43_192# hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_9/a_1226_296#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_8/D hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_25/a_1034_424#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfrtp_4_3/a_834_355# hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_13/a_1226_296#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_7/a_651_503# hr_16t4_mux_top_3/sky130_fd_sc_hs__dfrtp_4_3/a_1627_493#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_9/a_544_485# hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_29/a_206_368#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfrtp_4_3/a_812_138# hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_24/a_696_458#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_8/a_1226_296# hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_37/a_735_102#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_24/a_1034_424# hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_25/a_27_74#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_31/a_1178_124# hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_8/a_696_458#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_1/Q hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_29/a_437_503#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_7/a_1226_296# hr_16t4_mux_top_3/sky130_fd_sc_hs__dfrtp_4_3/a_37_78#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_23/a_1034_424# hr_16t4_mux_top_3/sky130_fd_sc_hs__a22o_1_23/a_230_79#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__a22o_1_3/a_132_392# hr_16t4_mux_top_3/sky130_fd_sc_hs__dfrtp_4_1/a_1627_493#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__a22o_1_17/a_132_392# hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_19/a_735_102#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_41/a_696_458# hr_16t4_mux_top_3/sky130_fd_sc_hs__dfrtp_4_1/a_1827_81#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_39/a_1034_424# hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_19/a_1141_508#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_9/a_27_74# hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_29/a_1226_296#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_18/a_27_74# hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_39/a_206_368#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_24/a_544_485# hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_31/a_696_458#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_37/a_1034_424# hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_18/a_1141_508#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_9/Q hr_16t4_mux_top_3/sky130_fd_sc_hs__a22o_1_23/a_52_123#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_8/a_544_485# hr_16t4_mux_top_3/sky130_fd_sc_hs__buf_2_3/X
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__buf_2_14/a_21_260# hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_5/a_1226_296#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_39/a_437_503# hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_23/a_696_458#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__buf_2_9/a_21_260# hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_5/a_206_368#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_7/a_696_458# hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_39/Q
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfrtp_4_3/a_1678_395# hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_41/a_544_485#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__clkbuf_2_29/a_43_192# hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_27/a_735_102#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfrtp_4_1/a_789_463# hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_15/a_1141_508#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__buf_2_1/X hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_41/a_27_74#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_5/a_437_503# hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_27/a_1226_296#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_3/a_735_102# hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_47/a_1178_124#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_9/a_1141_508# hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_3/a_1226_296#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_18/a_735_102# hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_31/a_544_485#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_35/a_1034_424# hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_13/a_1141_508#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__a22o_1_7/a_230_79# hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_3/a_27_74#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_46/a_1178_124# hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_8/a_1141_508#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfrtp_4_1/a_1678_395# hr_16t4_mux_top_3/sky130_fd_sc_hs__a22o_1_5/a_222_392#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_37/a_206_368# hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_23/a_544_485#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_29/a_651_503# hr_16t4_mux_top_3/sky130_fd_sc_hs__a22o_1_7/B2
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__a22o_1_19/a_222_392# hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_33/a_1034_424#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfrtp_4_1/a_834_355# hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_35/a_27_74#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_7/a_544_485# hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_45/a_1178_124#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_7/a_1141_508# hr_16t4_mux_top_3/sky130_fd_sc_hs__dfrtp_4_1/a_812_138#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_1/a_1226_296# hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_37/a_437_503#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__clkbuf_2_3/a_43_192# hr_16t4_mux_top_3/sky130_fd_sc_hs__a22o_1_7/a_52_123#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfrtp_4_3/a_1350_392# hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_19/a_206_368#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_29/a_1141_508# hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_25/a_1226_296#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_41/a_1178_124# hr_16t4_mux_top_3/sky130_fd_sc_hs__a22o_1_15/a_132_392#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_19/a_437_503# hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_46/a_27_74#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_39/a_651_503# hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_31/a_1034_424#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_24/a_1226_296# hr_16t4_mux_top_3/sky130_fd_sc_hs__dfrtp_4_1/a_1350_392#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_5/a_1141_508# hr_16t4_mux_top_3/sky130_fd_sc_hs__a22o_1_3/a_222_392#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__clkbuf_16_1/a_114_74# hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_47/a_735_102#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__a22o_1_17/a_222_392# hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_23/a_1226_296#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_5/a_651_503# hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_27/a_206_368#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_37/a_27_74# hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_29/a_696_458#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_35/a_735_102# hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_27/a_1141_508#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_3/a_206_368# hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_39/a_1226_296#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__buf_2_1/a_21_260# hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_3/a_1141_508#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_18/a_206_368# hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_27/a_437_503#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__clkbuf_2_21/a_43_192# hr_16t4_mux_top_3/sky130_fd_sc_hs__a22o_1_1/a_132_392#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_3/a_437_503# hr_16t4_mux_top_3/sky130_fd_sc_hs__dfrtp_4_1/a_124_78#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_37/a_1226_296# hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_24/a_27_74#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_1/a_735_102# hr_16t4_mux_top_3/sky130_fd_sc_hs__buf_2_5/a_21_260#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__a22o_1_14/a_132_392# hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_37/a_651_503#
+ hr_16t4_mux_top_3/sky130_fd_sc_hs__dfxtp_4_18/a_437_503# hr_16t4_mux_top_3/sky130_fd_sc_hs__dfrtp_4_3/a_1647_81#
+ hr_16t4_mux_top
Xsky130_fd_sc_hs__clkinv_8_9 DVSS: DVDD: DVDD: DVSS: prbs_generator_syn_1/out hr_16t4_mux_top_3/din[9]
+ sky130_fd_sc_hs__clkinv_8
Xsky130_fd_sc_hs__nand2_2_2 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__buf_2_33/A sky130_fd_sc_hs__nand2_2_3/B
+ sky130_fd_sc_hs__inv_4_11/Y sky130_fd_sc_hs__nand2_2_3/a_27_74# sky130_fd_sc_hs__nand2_2
Xsky130_fd_sc_hs__and2_4_0 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__and2_4_1/X hr_16t4_mux_top_3/clk_prbs
+ hr_16t4_mux_top_1/clk_prbs sky130_fd_sc_hs__and2_4_1/a_83_269# sky130_fd_sc_hs__and2_4_1/a_504_119#
+ sky130_fd_sc_hs__and2_4
Xsky130_fd_sc_hs__clkbuf_4_3 DVSS: DVDD: DVDD: DVSS: pi3_con[1] sky130_fd_sc_hs__clkbuf_8_9/A
+ sky130_fd_sc_hs__clkbuf_4_3/a_83_270# sky130_fd_sc_hs__clkbuf_4
Xsky130_fd_sc_hs__einvp_2_80 DVSS: DVDD: DVDD: DVSS: dout_p sky130_fd_sc_hs__einvp_2_97/A
+ sky130_fd_sc_hs__dlrtp_1_71/Q sky130_fd_sc_hs__einvp_2_81/a_263_323# sky130_fd_sc_hs__einvp_2_81/a_36_74#
+ sky130_fd_sc_hs__einvp_2_81/a_27_368# sky130_fd_sc_hs__einvp_2
Xsky130_fd_sc_hs__einvp_2_91 DVSS: DVDD: DVDD: DVSS: dout_p sky130_fd_sc_hs__einvp_2_99/A
+ sky130_fd_sc_hs__buf_2_63/X sky130_fd_sc_hs__einvp_2_91/a_263_323# sky130_fd_sc_hs__einvp_2_91/a_36_74#
+ sky130_fd_sc_hs__einvp_2_91/a_27_368# sky130_fd_sc_hs__einvp_2
Xsky130_fd_sc_hs__clkinv_4_3 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__clkinv_4_3/Y
+ sky130_fd_sc_hs__nor4_2_1/C sky130_fd_sc_hs__clkinv_4
Xsky130_fd_sc_hs__conb_1_90 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__conb_1_91/LO
+ sky130_fd_sc_hs__conb_1_91/HI sky130_fd_sc_hs__conb_1_91/a_165_290# sky130_fd_sc_hs__conb_1_91/a_21_290#
+ sky130_fd_sc_hs__conb_1
Xsky130_fd_sc_hs__dlrtp_1_102 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__dlrtp_1_103/Q
+ sky130_fd_sc_hs__dlrtp_1_9/GATE sky130_fd_sc_hs__conb_1_133/HI sky130_fd_sc_hs__dlrtp_1_103/D
+ sky130_fd_sc_hs__dlrtp_1_103/a_216_424# sky130_fd_sc_hs__dlrtp_1_103/a_759_508#
+ sky130_fd_sc_hs__dlrtp_1_103/a_565_74# sky130_fd_sc_hs__dlrtp_1_103/a_27_424# sky130_fd_sc_hs__dlrtp_1_103/a_1045_74#
+ sky130_fd_sc_hs__dlrtp_1_103/a_643_74# sky130_fd_sc_hs__dlrtp_1_103/a_817_48# sky130_fd_sc_hs__dlrtp_1_103/a_568_392#
+ sky130_fd_sc_hs__dlrtp_1_103/a_363_74# sky130_fd_sc_hs__dlrtp_1_103/a_769_74# sky130_fd_sc_hs__dlrtp_1
Xsky130_fd_sc_hs__dlrtp_1_113 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__buf_2_123/A
+ sky130_fd_sc_hs__dlrtp_1_9/GATE sky130_fd_sc_hs__conb_1_131/HI sky130_fd_sc_hs__o21bai_2_43/Y
+ sky130_fd_sc_hs__dlrtp_1_113/a_216_424# sky130_fd_sc_hs__dlrtp_1_113/a_759_508#
+ sky130_fd_sc_hs__dlrtp_1_113/a_565_74# sky130_fd_sc_hs__dlrtp_1_113/a_27_424# sky130_fd_sc_hs__dlrtp_1_113/a_1045_74#
+ sky130_fd_sc_hs__dlrtp_1_113/a_643_74# sky130_fd_sc_hs__dlrtp_1_113/a_817_48# sky130_fd_sc_hs__dlrtp_1_113/a_568_392#
+ sky130_fd_sc_hs__dlrtp_1_113/a_363_74# sky130_fd_sc_hs__dlrtp_1_113/a_769_74# sky130_fd_sc_hs__dlrtp_1
Xsky130_fd_sc_hs__dlrtp_1_124 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__einvp_2_49/TE
+ sky130_fd_sc_hs__clkbuf_2_3/A sky130_fd_sc_hs__conb_1_121/HI sky130_fd_sc_hs__inv_4_25/A
+ sky130_fd_sc_hs__dlrtp_1_125/a_216_424# sky130_fd_sc_hs__dlrtp_1_125/a_759_508#
+ sky130_fd_sc_hs__dlrtp_1_125/a_565_74# sky130_fd_sc_hs__dlrtp_1_125/a_27_424# sky130_fd_sc_hs__dlrtp_1_125/a_1045_74#
+ sky130_fd_sc_hs__dlrtp_1_125/a_643_74# sky130_fd_sc_hs__dlrtp_1_125/a_817_48# sky130_fd_sc_hs__dlrtp_1_125/a_568_392#
+ sky130_fd_sc_hs__dlrtp_1_125/a_363_74# sky130_fd_sc_hs__dlrtp_1_125/a_769_74# sky130_fd_sc_hs__dlrtp_1
Xsky130_fd_sc_hs__dlrtp_1_135 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__dlrtp_1_135/Q
+ sky130_fd_sc_hs__clkbuf_16_53/X sky130_fd_sc_hs__conb_1_135/HI sky130_fd_sc_hs__buf_2_141/X
+ sky130_fd_sc_hs__dlrtp_1_135/a_216_424# sky130_fd_sc_hs__dlrtp_1_135/a_759_508#
+ sky130_fd_sc_hs__dlrtp_1_135/a_565_74# sky130_fd_sc_hs__dlrtp_1_135/a_27_424# sky130_fd_sc_hs__dlrtp_1_135/a_1045_74#
+ sky130_fd_sc_hs__dlrtp_1_135/a_643_74# sky130_fd_sc_hs__dlrtp_1_135/a_817_48# sky130_fd_sc_hs__dlrtp_1_135/a_568_392#
+ sky130_fd_sc_hs__dlrtp_1_135/a_363_74# sky130_fd_sc_hs__dlrtp_1_135/a_769_74# sky130_fd_sc_hs__dlrtp_1
Xsky130_fd_sc_hs__dlrtp_1_146 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__dlrtp_1_147/Q
+ sky130_fd_sc_hs__clkbuf_16_53/X sky130_fd_sc_hs__conb_1_127/HI sky130_fd_sc_hs__inv_4_29/Y
+ sky130_fd_sc_hs__dlrtp_1_147/a_216_424# sky130_fd_sc_hs__dlrtp_1_147/a_759_508#
+ sky130_fd_sc_hs__dlrtp_1_147/a_565_74# sky130_fd_sc_hs__dlrtp_1_147/a_27_424# sky130_fd_sc_hs__dlrtp_1_147/a_1045_74#
+ sky130_fd_sc_hs__dlrtp_1_147/a_643_74# sky130_fd_sc_hs__dlrtp_1_147/a_817_48# sky130_fd_sc_hs__dlrtp_1_147/a_568_392#
+ sky130_fd_sc_hs__dlrtp_1_147/a_363_74# sky130_fd_sc_hs__dlrtp_1_147/a_769_74# sky130_fd_sc_hs__dlrtp_1
Xsky130_fd_sc_hs__dlrtp_1_157 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__dlrtp_1_157/Q
+ sky130_fd_sc_hs__clkbuf_16_53/X sky130_fd_sc_hs__conb_1_137/HI sky130_fd_sc_hs__dlrtp_1_157/D
+ sky130_fd_sc_hs__dlrtp_1_157/a_216_424# sky130_fd_sc_hs__dlrtp_1_157/a_759_508#
+ sky130_fd_sc_hs__dlrtp_1_157/a_565_74# sky130_fd_sc_hs__dlrtp_1_157/a_27_424# sky130_fd_sc_hs__dlrtp_1_157/a_1045_74#
+ sky130_fd_sc_hs__dlrtp_1_157/a_643_74# sky130_fd_sc_hs__dlrtp_1_157/a_817_48# sky130_fd_sc_hs__dlrtp_1_157/a_568_392#
+ sky130_fd_sc_hs__dlrtp_1_157/a_363_74# sky130_fd_sc_hs__dlrtp_1_157/a_769_74# sky130_fd_sc_hs__dlrtp_1
Xsky130_fd_sc_hs__inv_4_5 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__inv_4_5/Y ref_clk_ext_n
+ sky130_fd_sc_hs__inv_4
Xsky130_fd_sc_hs__dlrtp_1_70 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__dlrtp_1_71/Q
+ sky130_fd_sc_hs__clkbuf_16_53/A sky130_fd_sc_hs__conb_1_129/HI sky130_fd_sc_hs__dlrtp_1_71/D
+ sky130_fd_sc_hs__dlrtp_1_71/a_216_424# sky130_fd_sc_hs__dlrtp_1_71/a_759_508# sky130_fd_sc_hs__dlrtp_1_71/a_565_74#
+ sky130_fd_sc_hs__dlrtp_1_71/a_27_424# sky130_fd_sc_hs__dlrtp_1_71/a_1045_74# sky130_fd_sc_hs__dlrtp_1_71/a_643_74#
+ sky130_fd_sc_hs__dlrtp_1_71/a_817_48# sky130_fd_sc_hs__dlrtp_1_71/a_568_392# sky130_fd_sc_hs__dlrtp_1_71/a_363_74#
+ sky130_fd_sc_hs__dlrtp_1_71/a_769_74# sky130_fd_sc_hs__dlrtp_1
Xsky130_fd_sc_hs__dlrtp_1_81 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__dlrtp_1_81/Q
+ sky130_fd_sc_hs__clkbuf_16_53/X sky130_fd_sc_hs__conb_1_137/HI sky130_fd_sc_hs__buf_2_73/X
+ sky130_fd_sc_hs__dlrtp_1_81/a_216_424# sky130_fd_sc_hs__dlrtp_1_81/a_759_508# sky130_fd_sc_hs__dlrtp_1_81/a_565_74#
+ sky130_fd_sc_hs__dlrtp_1_81/a_27_424# sky130_fd_sc_hs__dlrtp_1_81/a_1045_74# sky130_fd_sc_hs__dlrtp_1_81/a_643_74#
+ sky130_fd_sc_hs__dlrtp_1_81/a_817_48# sky130_fd_sc_hs__dlrtp_1_81/a_568_392# sky130_fd_sc_hs__dlrtp_1_81/a_363_74#
+ sky130_fd_sc_hs__dlrtp_1_81/a_769_74# sky130_fd_sc_hs__dlrtp_1
Xsky130_fd_sc_hs__dlrtp_1_92 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__buf_2_93/A sky130_fd_sc_hs__dlrtp_1_9/GATE
+ sky130_fd_sc_hs__conb_1_95/HI sky130_fd_sc_hs__buf_2_107/X sky130_fd_sc_hs__dlrtp_1_93/a_216_424#
+ sky130_fd_sc_hs__dlrtp_1_93/a_759_508# sky130_fd_sc_hs__dlrtp_1_93/a_565_74# sky130_fd_sc_hs__dlrtp_1_93/a_27_424#
+ sky130_fd_sc_hs__dlrtp_1_93/a_1045_74# sky130_fd_sc_hs__dlrtp_1_93/a_643_74# sky130_fd_sc_hs__dlrtp_1_93/a_817_48#
+ sky130_fd_sc_hs__dlrtp_1_93/a_568_392# sky130_fd_sc_hs__dlrtp_1_93/a_363_74# sky130_fd_sc_hs__dlrtp_1_93/a_769_74#
+ sky130_fd_sc_hs__dlrtp_1
Xsky130_fd_sc_hs__clkbuf_2_0 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__dlrtp_1_27/D
+ sky130_fd_sc_hs__o21bai_4_3/Y sky130_fd_sc_hs__clkbuf_2_1/a_43_192# sky130_fd_sc_hs__clkbuf_2
Xsky130_fd_sc_hs__clkbuf_2_11 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__dlrtp_1_55/D
+ sky130_fd_sc_hs__o21ai_2_11/Y sky130_fd_sc_hs__clkbuf_2_11/a_43_192# sky130_fd_sc_hs__clkbuf_2
Xsky130_fd_sc_hs__clkbuf_2_22 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__dlrtp_1_157/D
+ sky130_fd_sc_hs__o21ai_2_25/Y sky130_fd_sc_hs__clkbuf_2_23/a_43_192# sky130_fd_sc_hs__clkbuf_2
Xsky130_fd_sc_hs__clkbuf_2_33 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__dlrtp_1_9/D
+ sky130_fd_sc_hs__buf_2_95/X sky130_fd_sc_hs__clkbuf_2_33/a_43_192# sky130_fd_sc_hs__clkbuf_2
Xsky130_fd_sc_hs__clkbuf_2_44 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__dlrtp_1_19/D
+ sky130_fd_sc_hs__o21bai_2_37/Y sky130_fd_sc_hs__clkbuf_2_45/a_43_192# sky130_fd_sc_hs__clkbuf_2
Xsky130_fd_sc_hs__clkbuf_2_55 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__dlrtp_1_121/D
+ sky130_fd_sc_hs__o21ai_2_47/Y sky130_fd_sc_hs__clkbuf_2_55/a_43_192# sky130_fd_sc_hs__clkbuf_2
Xsky130_fd_sc_hs__clkbuf_2_66 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__dlrtp_1_143/D
+ sky130_fd_sc_hs__buf_2_147/X sky130_fd_sc_hs__clkbuf_2_67/a_43_192# sky130_fd_sc_hs__clkbuf_2
Xsky130_fd_sc_hs__clkinv_2_0 DVSS: DVDD: DVDD: DVSS: test_mux_clk_I sky130_fd_sc_hs__buf_2_3/X
+ sky130_fd_sc_hs__clkinv_2
Xsky130_fd_sc_hs__buf_2_2 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__buf_2_3/A sky130_fd_sc_hs__buf_2_3/X
+ sky130_fd_sc_hs__buf_2_3/a_21_260# sky130_fd_sc_hs__buf_2
Xsky130_fd_sc_hs__dlrtp_1_4 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__dlrtp_1_5/Q sky130_fd_sc_hs__dlrtp_1_9/GATE
+ sky130_fd_sc_hs__conb_1_117/HI sky130_fd_sc_hs__buf_2_87/A sky130_fd_sc_hs__dlrtp_1_5/a_216_424#
+ sky130_fd_sc_hs__dlrtp_1_5/a_759_508# sky130_fd_sc_hs__dlrtp_1_5/a_565_74# sky130_fd_sc_hs__dlrtp_1_5/a_27_424#
+ sky130_fd_sc_hs__dlrtp_1_5/a_1045_74# sky130_fd_sc_hs__dlrtp_1_5/a_643_74# sky130_fd_sc_hs__dlrtp_1_5/a_817_48#
+ sky130_fd_sc_hs__dlrtp_1_5/a_568_392# sky130_fd_sc_hs__dlrtp_1_5/a_363_74# sky130_fd_sc_hs__dlrtp_1_5/a_769_74#
+ sky130_fd_sc_hs__dlrtp_1
Xsky130_fd_sc_hs__buf_2_40 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__buf_2_41/A sky130_fd_sc_hs__buf_2_41/X
+ sky130_fd_sc_hs__buf_2_41/a_21_260# sky130_fd_sc_hs__buf_2
Xsky130_fd_sc_hs__buf_2_51 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__buf_2_51/A sky130_fd_sc_hs__buf_2_51/X
+ sky130_fd_sc_hs__buf_2_51/a_21_260# sky130_fd_sc_hs__buf_2
Xsky130_fd_sc_hs__buf_2_62 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__buf_2_63/A sky130_fd_sc_hs__buf_2_63/X
+ sky130_fd_sc_hs__buf_2_63/a_21_260# sky130_fd_sc_hs__buf_2
Xsky130_fd_sc_hs__buf_2_73 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__buf_2_79/X sky130_fd_sc_hs__buf_2_73/X
+ sky130_fd_sc_hs__buf_2_73/a_21_260# sky130_fd_sc_hs__buf_2
Xsky130_fd_sc_hs__buf_2_84 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__buf_2_85/A sky130_fd_sc_hs__buf_2_85/X
+ sky130_fd_sc_hs__buf_2_85/a_21_260# sky130_fd_sc_hs__buf_2
Xsky130_fd_sc_hs__buf_2_95 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__buf_2_95/A sky130_fd_sc_hs__buf_2_95/X
+ sky130_fd_sc_hs__buf_2_95/a_21_260# sky130_fd_sc_hs__buf_2
Xsky130_fd_sc_hs__o21bai_2_20 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__buf_8_3/X sky130_fd_sc_hs__o21bai_4_3/A2
+ sky130_fd_sc_hs__dlrtp_1_9/D sky130_fd_sc_hs__dlrtp_1_8/D sky130_fd_sc_hs__o21bai_2_21/a_27_74#
+ sky130_fd_sc_hs__o21bai_2_21/a_225_74# sky130_fd_sc_hs__o21bai_2_21/a_507_368# sky130_fd_sc_hs__o21bai_2
Xsky130_fd_sc_hs__o21bai_2_31 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__o21ai_4_1/A1
+ sky130_fd_sc_hs__o21bai_4_3/A2 sky130_fd_sc_hs__dlrtp_1_103/D sky130_fd_sc_hs__o21bai_2_31/Y
+ sky130_fd_sc_hs__o21bai_2_31/a_27_74# sky130_fd_sc_hs__o21bai_2_31/a_225_74# sky130_fd_sc_hs__o21bai_2_31/a_507_368#
+ sky130_fd_sc_hs__o21bai_2
Xsky130_fd_sc_hs__o21bai_2_42 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__nand2_2_15/B
+ sky130_fd_sc_hs__clkbuf_4_81/X sky130_fd_sc_hs__dlrtp_1_115/D sky130_fd_sc_hs__o21bai_2_43/Y
+ sky130_fd_sc_hs__o21bai_2_43/a_27_74# sky130_fd_sc_hs__o21bai_2_43/a_225_74# sky130_fd_sc_hs__o21bai_2_43/a_507_368#
+ sky130_fd_sc_hs__o21bai_2
Xsky130_fd_sc_hs__o21bai_2_53 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__clkinv_4_3/Y
+ sky130_fd_sc_hs__nand2_2_21/B sky130_fd_sc_hs__dlrtp_1_121/D sky130_fd_sc_hs__o21bai_2_53/Y
+ sky130_fd_sc_hs__o21bai_2_53/a_27_74# sky130_fd_sc_hs__o21bai_2_53/a_225_74# sky130_fd_sc_hs__o21bai_2_53/a_507_368#
+ sky130_fd_sc_hs__o21bai_2
Xsky130_fd_sc_hs__o21bai_2_64 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__nand2_2_9/B
+ sky130_fd_sc_hs__o21bai_4_7/A1 sky130_fd_sc_hs__buf_2_47/X sky130_fd_sc_hs__dlrtp_1_74/D
+ sky130_fd_sc_hs__o21bai_2_66/a_27_74# sky130_fd_sc_hs__o21bai_2_66/a_225_74# sky130_fd_sc_hs__o21bai_2_66/a_507_368#
+ sky130_fd_sc_hs__o21bai_2
Xsky130_fd_sc_hs__conb_1_240 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__conb_1_241/LO
+ sky130_fd_sc_hs__conb_1_241/HI sky130_fd_sc_hs__conb_1_241/a_165_290# sky130_fd_sc_hs__conb_1_241/a_21_290#
+ sky130_fd_sc_hs__conb_1
Xsky130_fd_sc_hs__conb_1_251 DVSS: DVDD: DVDD: DVSS: prbs_generator_syn_27/eqn[28]
+ sky130_fd_sc_hs__conb_1_251/HI sky130_fd_sc_hs__conb_1_251/a_165_290# sky130_fd_sc_hs__conb_1_251/a_21_290#
+ sky130_fd_sc_hs__conb_1
Xsky130_fd_sc_hs__conb_1_262 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__conb_1_263/LO
+ sky130_fd_sc_hs__conb_1_263/HI sky130_fd_sc_hs__conb_1_263/a_165_290# sky130_fd_sc_hs__conb_1_263/a_21_290#
+ sky130_fd_sc_hs__conb_1
Xsky130_fd_sc_hs__conb_1_273 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__conb_1_273/LO
+ sky130_fd_sc_hs__conb_1_273/HI sky130_fd_sc_hs__conb_1_273/a_165_290# sky130_fd_sc_hs__conb_1_273/a_21_290#
+ sky130_fd_sc_hs__conb_1
Xsky130_fd_sc_hs__clkbuf_8_10 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__clkbuf_8_11/X
+ sky130_fd_sc_hs__clkbuf_4_1/X sky130_fd_sc_hs__clkbuf_8_11/a_125_368# sky130_fd_sc_hs__clkbuf_8
Xsky130_fd_sc_hs__clkbuf_8_21 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__clkbuf_8_21/X
+ sky130_fd_sc_hs__clkbuf_8_21/A sky130_fd_sc_hs__clkbuf_8_21/a_125_368# sky130_fd_sc_hs__clkbuf_8
Xsky130_fd_sc_hs__clkbuf_8_32 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__nand2_2_11/B
+ sky130_fd_sc_hs__buf_2_77/X sky130_fd_sc_hs__clkbuf_8_33/a_125_368# sky130_fd_sc_hs__clkbuf_8
Xsky130_fd_sc_hs__clkbuf_8_43 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__o21bai_4_3/A2
+ sky130_fd_sc_hs__nand2_2_25/Y sky130_fd_sc_hs__clkbuf_8_43/a_125_368# sky130_fd_sc_hs__clkbuf_8
Xsky130_fd_sc_hs__clkbuf_8_54 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__inv_4_29/A
+ sky130_fd_sc_hs__or4_2_1/X sky130_fd_sc_hs__clkbuf_8_55/a_125_368# sky130_fd_sc_hs__clkbuf_8
Xsky130_fd_sc_hs__clkbuf_8_65 DVSS: DVDD: DVDD: DVSS: fine_freq_track_1/aux_osc_en
+ aux_osc_en sky130_fd_sc_hs__clkbuf_8_65/a_125_368# sky130_fd_sc_hs__clkbuf_8
Xsky130_fd_sc_hs__clkbuf_8_76 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__clkbuf_8_77/X
+ sky130_fd_sc_hs__clkbuf_8_77/A sky130_fd_sc_hs__clkbuf_8_77/a_125_368# sky130_fd_sc_hs__clkbuf_8
Xsky130_fd_sc_hs__clkbuf_8_87 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__einvp_8_5/TE
+ test_mux_select[2] sky130_fd_sc_hs__clkbuf_8_87/a_125_368# sky130_fd_sc_hs__clkbuf_8
Xsky130_fd_sc_hs__clkbuf_8_98 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__clkbuf_8_99/X
+ CTL_BUF_N[0] sky130_fd_sc_hs__clkbuf_8_99/a_125_368# sky130_fd_sc_hs__clkbuf_8
Xsky130_fd_sc_hs__nor2_4_2 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__nor2_4_3/Y sky130_fd_sc_hs__nor2_4_3/A
+ sky130_fd_sc_hs__nor2_4_3/B sky130_fd_sc_hs__nor2_4_3/a_27_368# sky130_fd_sc_hs__nor2_4
Xsky130_fd_sc_hs__einvp_8_7 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__inv_4_39/A sky130_fd_sc_hs__einvp_8_7/TE
+ osc_core_1/osc_hold sky130_fd_sc_hs__einvp_8_7/a_802_323# sky130_fd_sc_hs__einvp_8_7/a_27_74#
+ sky130_fd_sc_hs__einvp_8_7/a_27_368# sky130_fd_sc_hs__einvp_8
Xsky130_fd_sc_hs__nand2_2_3 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__buf_2_33/A sky130_fd_sc_hs__nand2_2_3/B
+ sky130_fd_sc_hs__inv_4_11/Y sky130_fd_sc_hs__nand2_2_3/a_27_74# sky130_fd_sc_hs__nand2_2
Xsky130_fd_sc_hs__and2_4_1 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__and2_4_1/X hr_16t4_mux_top_3/clk_prbs
+ hr_16t4_mux_top_1/clk_prbs sky130_fd_sc_hs__and2_4_1/a_83_269# sky130_fd_sc_hs__and2_4_1/a_504_119#
+ sky130_fd_sc_hs__and2_4
Xsky130_fd_sc_hs__clkbuf_4_4 DVSS: DVDD: DVDD: DVSS: pi3_con[2] sky130_fd_sc_hs__clkbuf_8_7/A
+ sky130_fd_sc_hs__clkbuf_4_5/a_83_270# sky130_fd_sc_hs__clkbuf_4
Xsky130_fd_sc_hs__einvp_2_70 DVSS: DVDD: DVDD: DVSS: dout_p sky130_fd_sc_hs__einvp_2_97/A
+ sky130_fd_sc_hs__dlrtp_1_58/Q sky130_fd_sc_hs__einvp_2_71/a_263_323# sky130_fd_sc_hs__einvp_2_71/a_36_74#
+ sky130_fd_sc_hs__einvp_2_71/a_27_368# sky130_fd_sc_hs__einvp_2
Xsky130_fd_sc_hs__einvp_2_81 DVSS: DVDD: DVDD: DVSS: dout_p sky130_fd_sc_hs__einvp_2_97/A
+ sky130_fd_sc_hs__dlrtp_1_71/Q sky130_fd_sc_hs__einvp_2_81/a_263_323# sky130_fd_sc_hs__einvp_2_81/a_36_74#
+ sky130_fd_sc_hs__einvp_2_81/a_27_368# sky130_fd_sc_hs__einvp_2
Xsky130_fd_sc_hs__einvp_2_92 DVSS: DVDD: DVDD: DVSS: dout_p sky130_fd_sc_hs__einvp_2_97/A
+ sky130_fd_sc_hs__dlrtp_1_77/Q sky130_fd_sc_hs__einvp_2_93/a_263_323# sky130_fd_sc_hs__einvp_2_93/a_36_74#
+ sky130_fd_sc_hs__einvp_2_93/a_27_368# sky130_fd_sc_hs__einvp_2
Xsky130_fd_sc_hs__clkinv_4_4 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__clkinv_4_5/Y
+ sky130_fd_sc_hs__nor4_2_1/A sky130_fd_sc_hs__clkinv_4
Xsky130_fd_sc_hs__conb_1_80 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__conb_1_81/LO
+ prbs_generator_syn_11/cke sky130_fd_sc_hs__conb_1_81/a_165_290# sky130_fd_sc_hs__conb_1_81/a_21_290#
+ sky130_fd_sc_hs__conb_1
Xsky130_fd_sc_hs__conb_1_91 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__conb_1_91/LO
+ sky130_fd_sc_hs__conb_1_91/HI sky130_fd_sc_hs__conb_1_91/a_165_290# sky130_fd_sc_hs__conb_1_91/a_21_290#
+ sky130_fd_sc_hs__conb_1
Xsky130_fd_sc_hs__dlrtp_1_103 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__dlrtp_1_103/Q
+ sky130_fd_sc_hs__dlrtp_1_9/GATE sky130_fd_sc_hs__conb_1_133/HI sky130_fd_sc_hs__dlrtp_1_103/D
+ sky130_fd_sc_hs__dlrtp_1_103/a_216_424# sky130_fd_sc_hs__dlrtp_1_103/a_759_508#
+ sky130_fd_sc_hs__dlrtp_1_103/a_565_74# sky130_fd_sc_hs__dlrtp_1_103/a_27_424# sky130_fd_sc_hs__dlrtp_1_103/a_1045_74#
+ sky130_fd_sc_hs__dlrtp_1_103/a_643_74# sky130_fd_sc_hs__dlrtp_1_103/a_817_48# sky130_fd_sc_hs__dlrtp_1_103/a_568_392#
+ sky130_fd_sc_hs__dlrtp_1_103/a_363_74# sky130_fd_sc_hs__dlrtp_1_103/a_769_74# sky130_fd_sc_hs__dlrtp_1
Xsky130_fd_sc_hs__dlrtp_1_114 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__buf_2_125/A
+ sky130_fd_sc_hs__dlrtp_1_9/GATE sky130_fd_sc_hs__conb_1_131/HI sky130_fd_sc_hs__dlrtp_1_115/D
+ sky130_fd_sc_hs__dlrtp_1_115/a_216_424# sky130_fd_sc_hs__dlrtp_1_115/a_759_508#
+ sky130_fd_sc_hs__dlrtp_1_115/a_565_74# sky130_fd_sc_hs__dlrtp_1_115/a_27_424# sky130_fd_sc_hs__dlrtp_1_115/a_1045_74#
+ sky130_fd_sc_hs__dlrtp_1_115/a_643_74# sky130_fd_sc_hs__dlrtp_1_115/a_817_48# sky130_fd_sc_hs__dlrtp_1_115/a_568_392#
+ sky130_fd_sc_hs__dlrtp_1_115/a_363_74# sky130_fd_sc_hs__dlrtp_1_115/a_769_74# sky130_fd_sc_hs__dlrtp_1
Xsky130_fd_sc_hs__dlrtp_1_125 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__einvp_2_49/TE
+ sky130_fd_sc_hs__clkbuf_2_3/A sky130_fd_sc_hs__conb_1_121/HI sky130_fd_sc_hs__inv_4_25/A
+ sky130_fd_sc_hs__dlrtp_1_125/a_216_424# sky130_fd_sc_hs__dlrtp_1_125/a_759_508#
+ sky130_fd_sc_hs__dlrtp_1_125/a_565_74# sky130_fd_sc_hs__dlrtp_1_125/a_27_424# sky130_fd_sc_hs__dlrtp_1_125/a_1045_74#
+ sky130_fd_sc_hs__dlrtp_1_125/a_643_74# sky130_fd_sc_hs__dlrtp_1_125/a_817_48# sky130_fd_sc_hs__dlrtp_1_125/a_568_392#
+ sky130_fd_sc_hs__dlrtp_1_125/a_363_74# sky130_fd_sc_hs__dlrtp_1_125/a_769_74# sky130_fd_sc_hs__dlrtp_1
Xsky130_fd_sc_hs__dlrtp_1_136 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__dlrtp_1_137/Q
+ sky130_fd_sc_hs__clkbuf_16_53/X sky130_fd_sc_hs__conb_1_135/HI sky130_fd_sc_hs__buf_2_145/X
+ sky130_fd_sc_hs__dlrtp_1_137/a_216_424# sky130_fd_sc_hs__dlrtp_1_137/a_759_508#
+ sky130_fd_sc_hs__dlrtp_1_137/a_565_74# sky130_fd_sc_hs__dlrtp_1_137/a_27_424# sky130_fd_sc_hs__dlrtp_1_137/a_1045_74#
+ sky130_fd_sc_hs__dlrtp_1_137/a_643_74# sky130_fd_sc_hs__dlrtp_1_137/a_817_48# sky130_fd_sc_hs__dlrtp_1_137/a_568_392#
+ sky130_fd_sc_hs__dlrtp_1_137/a_363_74# sky130_fd_sc_hs__dlrtp_1_137/a_769_74# sky130_fd_sc_hs__dlrtp_1
Xsky130_fd_sc_hs__dlrtp_1_147 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__dlrtp_1_147/Q
+ sky130_fd_sc_hs__clkbuf_16_53/X sky130_fd_sc_hs__conb_1_127/HI sky130_fd_sc_hs__inv_4_29/Y
+ sky130_fd_sc_hs__dlrtp_1_147/a_216_424# sky130_fd_sc_hs__dlrtp_1_147/a_759_508#
+ sky130_fd_sc_hs__dlrtp_1_147/a_565_74# sky130_fd_sc_hs__dlrtp_1_147/a_27_424# sky130_fd_sc_hs__dlrtp_1_147/a_1045_74#
+ sky130_fd_sc_hs__dlrtp_1_147/a_643_74# sky130_fd_sc_hs__dlrtp_1_147/a_817_48# sky130_fd_sc_hs__dlrtp_1_147/a_568_392#
+ sky130_fd_sc_hs__dlrtp_1_147/a_363_74# sky130_fd_sc_hs__dlrtp_1_147/a_769_74# sky130_fd_sc_hs__dlrtp_1
Xsky130_fd_sc_hs__dlrtp_1_158 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__buf_2_161/A
+ sky130_fd_sc_hs__clkbuf_16_53/X sky130_fd_sc_hs__conb_1_137/HI sky130_fd_sc_hs__buf_2_75/X
+ sky130_fd_sc_hs__dlrtp_1_159/a_216_424# sky130_fd_sc_hs__dlrtp_1_159/a_759_508#
+ sky130_fd_sc_hs__dlrtp_1_159/a_565_74# sky130_fd_sc_hs__dlrtp_1_159/a_27_424# sky130_fd_sc_hs__dlrtp_1_159/a_1045_74#
+ sky130_fd_sc_hs__dlrtp_1_159/a_643_74# sky130_fd_sc_hs__dlrtp_1_159/a_817_48# sky130_fd_sc_hs__dlrtp_1_159/a_568_392#
+ sky130_fd_sc_hs__dlrtp_1_159/a_363_74# sky130_fd_sc_hs__dlrtp_1_159/a_769_74# sky130_fd_sc_hs__dlrtp_1
Xsky130_fd_sc_hs__inv_4_6 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__inv_4_7/Y fine_control_avg_window_select[1]
+ sky130_fd_sc_hs__inv_4
Xsky130_fd_sc_hs__dlrtp_1_60 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__buf_2_31/A sky130_fd_sc_hs__clkbuf_16_53/A
+ sky130_fd_sc_hs__conb_1_125/HI sky130_fd_sc_hs__buf_2_59/X sky130_fd_sc_hs__dlrtp_1_61/a_216_424#
+ sky130_fd_sc_hs__dlrtp_1_61/a_759_508# sky130_fd_sc_hs__dlrtp_1_61/a_565_74# sky130_fd_sc_hs__dlrtp_1_61/a_27_424#
+ sky130_fd_sc_hs__dlrtp_1_61/a_1045_74# sky130_fd_sc_hs__dlrtp_1_61/a_643_74# sky130_fd_sc_hs__dlrtp_1_61/a_817_48#
+ sky130_fd_sc_hs__dlrtp_1_61/a_568_392# sky130_fd_sc_hs__dlrtp_1_61/a_363_74# sky130_fd_sc_hs__dlrtp_1_61/a_769_74#
+ sky130_fd_sc_hs__dlrtp_1
Xsky130_fd_sc_hs__dlrtp_1_71 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__dlrtp_1_71/Q
+ sky130_fd_sc_hs__clkbuf_16_53/A sky130_fd_sc_hs__conb_1_129/HI sky130_fd_sc_hs__dlrtp_1_71/D
+ sky130_fd_sc_hs__dlrtp_1_71/a_216_424# sky130_fd_sc_hs__dlrtp_1_71/a_759_508# sky130_fd_sc_hs__dlrtp_1_71/a_565_74#
+ sky130_fd_sc_hs__dlrtp_1_71/a_27_424# sky130_fd_sc_hs__dlrtp_1_71/a_1045_74# sky130_fd_sc_hs__dlrtp_1_71/a_643_74#
+ sky130_fd_sc_hs__dlrtp_1_71/a_817_48# sky130_fd_sc_hs__dlrtp_1_71/a_568_392# sky130_fd_sc_hs__dlrtp_1_71/a_363_74#
+ sky130_fd_sc_hs__dlrtp_1_71/a_769_74# sky130_fd_sc_hs__dlrtp_1
Xsky130_fd_sc_hs__dlrtp_1_82 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__buf_2_63/A sky130_fd_sc_hs__clkbuf_16_53/X
+ sky130_fd_sc_hs__conb_1_137/HI sky130_fd_sc_hs__o21ai_2_17/Y sky130_fd_sc_hs__dlrtp_1_83/a_216_424#
+ sky130_fd_sc_hs__dlrtp_1_83/a_759_508# sky130_fd_sc_hs__dlrtp_1_83/a_565_74# sky130_fd_sc_hs__dlrtp_1_83/a_27_424#
+ sky130_fd_sc_hs__dlrtp_1_83/a_1045_74# sky130_fd_sc_hs__dlrtp_1_83/a_643_74# sky130_fd_sc_hs__dlrtp_1_83/a_817_48#
+ sky130_fd_sc_hs__dlrtp_1_83/a_568_392# sky130_fd_sc_hs__dlrtp_1_83/a_363_74# sky130_fd_sc_hs__dlrtp_1_83/a_769_74#
+ sky130_fd_sc_hs__dlrtp_1
Xsky130_fd_sc_hs__dlrtp_1_93 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__buf_2_93/A sky130_fd_sc_hs__dlrtp_1_9/GATE
+ sky130_fd_sc_hs__conb_1_95/HI sky130_fd_sc_hs__buf_2_107/X sky130_fd_sc_hs__dlrtp_1_93/a_216_424#
+ sky130_fd_sc_hs__dlrtp_1_93/a_759_508# sky130_fd_sc_hs__dlrtp_1_93/a_565_74# sky130_fd_sc_hs__dlrtp_1_93/a_27_424#
+ sky130_fd_sc_hs__dlrtp_1_93/a_1045_74# sky130_fd_sc_hs__dlrtp_1_93/a_643_74# sky130_fd_sc_hs__dlrtp_1_93/a_817_48#
+ sky130_fd_sc_hs__dlrtp_1_93/a_568_392# sky130_fd_sc_hs__dlrtp_1_93/a_363_74# sky130_fd_sc_hs__dlrtp_1_93/a_769_74#
+ sky130_fd_sc_hs__dlrtp_1
Xsky130_fd_sc_hs__clkbuf_2_1 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__dlrtp_1_27/D
+ sky130_fd_sc_hs__o21bai_4_3/Y sky130_fd_sc_hs__clkbuf_2_1/a_43_192# sky130_fd_sc_hs__clkbuf_2
Xsky130_fd_sc_hs__clkbuf_2_12 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__dlrtp_1_71/D
+ sky130_fd_sc_hs__o21bai_2_13/Y sky130_fd_sc_hs__clkbuf_2_13/a_43_192# sky130_fd_sc_hs__clkbuf_2
Xsky130_fd_sc_hs__clkbuf_2_23 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__dlrtp_1_157/D
+ sky130_fd_sc_hs__o21ai_2_25/Y sky130_fd_sc_hs__clkbuf_2_23/a_43_192# sky130_fd_sc_hs__clkbuf_2
Xsky130_fd_sc_hs__clkbuf_2_34 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__dlrtp_1_103/D
+ sky130_fd_sc_hs__o21ai_4_1/Y sky130_fd_sc_hs__clkbuf_2_35/a_43_192# sky130_fd_sc_hs__clkbuf_2
Xsky130_fd_sc_hs__clkbuf_2_45 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__dlrtp_1_19/D
+ sky130_fd_sc_hs__o21bai_2_37/Y sky130_fd_sc_hs__clkbuf_2_45/a_43_192# sky130_fd_sc_hs__clkbuf_2
Xsky130_fd_sc_hs__clkbuf_2_56 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__buf_2_131/A
+ sky130_fd_sc_hs__nor4_2_1/Y sky130_fd_sc_hs__clkbuf_2_57/a_43_192# sky130_fd_sc_hs__clkbuf_2
Xsky130_fd_sc_hs__clkbuf_2_67 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__dlrtp_1_143/D
+ sky130_fd_sc_hs__buf_2_147/X sky130_fd_sc_hs__clkbuf_2_67/a_43_192# sky130_fd_sc_hs__clkbuf_2
Xsky130_fd_sc_hs__clkinv_2_1 DVSS: DVDD: DVDD: DVSS: test_mux_clk_I sky130_fd_sc_hs__buf_2_3/X
+ sky130_fd_sc_hs__clkinv_2
Xsky130_fd_sc_hs__buf_2_3 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__buf_2_3/A sky130_fd_sc_hs__buf_2_3/X
+ sky130_fd_sc_hs__buf_2_3/a_21_260# sky130_fd_sc_hs__buf_2
Xsky130_fd_sc_hs__dlrtp_1_5 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__dlrtp_1_5/Q sky130_fd_sc_hs__dlrtp_1_9/GATE
+ sky130_fd_sc_hs__conb_1_117/HI sky130_fd_sc_hs__buf_2_87/A sky130_fd_sc_hs__dlrtp_1_5/a_216_424#
+ sky130_fd_sc_hs__dlrtp_1_5/a_759_508# sky130_fd_sc_hs__dlrtp_1_5/a_565_74# sky130_fd_sc_hs__dlrtp_1_5/a_27_424#
+ sky130_fd_sc_hs__dlrtp_1_5/a_1045_74# sky130_fd_sc_hs__dlrtp_1_5/a_643_74# sky130_fd_sc_hs__dlrtp_1_5/a_817_48#
+ sky130_fd_sc_hs__dlrtp_1_5/a_568_392# sky130_fd_sc_hs__dlrtp_1_5/a_363_74# sky130_fd_sc_hs__dlrtp_1_5/a_769_74#
+ sky130_fd_sc_hs__dlrtp_1
Xsky130_fd_sc_hs__buf_2_30 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__buf_2_30/A sky130_fd_sc_hs__buf_2_30/X
+ sky130_fd_sc_hs__buf_2_30/a_21_260# sky130_fd_sc_hs__buf_2
Xsky130_fd_sc_hs__buf_2_41 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__buf_2_41/A sky130_fd_sc_hs__buf_2_41/X
+ sky130_fd_sc_hs__buf_2_41/a_21_260# sky130_fd_sc_hs__buf_2
Xsky130_fd_sc_hs__buf_2_52 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__buf_2_61/X sky130_fd_sc_hs__buf_2_53/X
+ sky130_fd_sc_hs__buf_2_53/a_21_260# sky130_fd_sc_hs__buf_2
Xsky130_fd_sc_hs__buf_2_63 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__buf_2_63/A sky130_fd_sc_hs__buf_2_63/X
+ sky130_fd_sc_hs__buf_2_63/a_21_260# sky130_fd_sc_hs__buf_2
Xsky130_fd_sc_hs__buf_2_74 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__buf_2_75/A sky130_fd_sc_hs__buf_2_75/X
+ sky130_fd_sc_hs__buf_2_75/a_21_260# sky130_fd_sc_hs__buf_2
Xsky130_fd_sc_hs__buf_2_85 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__buf_2_85/A sky130_fd_sc_hs__buf_2_85/X
+ sky130_fd_sc_hs__buf_2_85/a_21_260# sky130_fd_sc_hs__buf_2
Xsky130_fd_sc_hs__buf_2_96 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__buf_2_98/A sky130_fd_sc_hs__buf_2_98/X
+ sky130_fd_sc_hs__buf_2_98/a_21_260# sky130_fd_sc_hs__buf_2
Xsky130_fd_sc_hs__o21bai_2_10 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__inv_8_1/Y sky130_fd_sc_hs__nand2_2_11/B
+ sky130_fd_sc_hs__dlrtp_1_69/D sky130_fd_sc_hs__buf_2_61/A sky130_fd_sc_hs__o21bai_2_11/a_27_74#
+ sky130_fd_sc_hs__o21bai_2_11/a_225_74# sky130_fd_sc_hs__o21bai_2_11/a_507_368# sky130_fd_sc_hs__o21bai_2
Xsky130_fd_sc_hs__o21bai_2_21 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__buf_8_3/X sky130_fd_sc_hs__o21bai_4_3/A2
+ sky130_fd_sc_hs__dlrtp_1_9/D sky130_fd_sc_hs__dlrtp_1_8/D sky130_fd_sc_hs__o21bai_2_21/a_27_74#
+ sky130_fd_sc_hs__o21bai_2_21/a_225_74# sky130_fd_sc_hs__o21bai_2_21/a_507_368# sky130_fd_sc_hs__o21bai_2
Xsky130_fd_sc_hs__o21bai_2_32 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__clkinv_4_3/Y
+ sky130_fd_sc_hs__or2b_2_3/A sky130_fd_sc_hs__dlrtp_1_99/D sky130_fd_sc_hs__buf_2_111/A
+ sky130_fd_sc_hs__o21bai_2_33/a_27_74# sky130_fd_sc_hs__o21bai_2_33/a_225_74# sky130_fd_sc_hs__o21bai_2_33/a_507_368#
+ sky130_fd_sc_hs__o21bai_2
Xsky130_fd_sc_hs__o21bai_2_43 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__nand2_2_15/B
+ sky130_fd_sc_hs__clkbuf_4_81/X sky130_fd_sc_hs__dlrtp_1_115/D sky130_fd_sc_hs__o21bai_2_43/Y
+ sky130_fd_sc_hs__o21bai_2_43/a_27_74# sky130_fd_sc_hs__o21bai_2_43/a_225_74# sky130_fd_sc_hs__o21bai_2_43/a_507_368#
+ sky130_fd_sc_hs__o21bai_2
Xsky130_fd_sc_hs__o21bai_2_54 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__o21bai_4_3/A2
+ sky130_fd_sc_hs__nand2_2_21/B sky130_fd_sc_hs__dlrtp_1_35/D sky130_fd_sc_hs__buf_2_133/A
+ sky130_fd_sc_hs__o21bai_2_55/a_27_74# sky130_fd_sc_hs__o21bai_2_55/a_225_74# sky130_fd_sc_hs__o21bai_2_55/a_507_368#
+ sky130_fd_sc_hs__o21bai_2
Xsky130_fd_sc_hs__o21bai_2_65 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__o21bai_2_5/A1
+ sky130_fd_sc_hs__nand2_2_9/B sky130_fd_sc_hs__buf_2_47/X sky130_fd_sc_hs__o21bai_2_67/Y
+ sky130_fd_sc_hs__o21bai_2_67/a_27_74# sky130_fd_sc_hs__o21bai_2_67/a_225_74# sky130_fd_sc_hs__o21bai_2_67/a_507_368#
+ sky130_fd_sc_hs__o21bai_2
Xsky130_fd_sc_hs__conb_1_230 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__conb_1_231/LO
+ sky130_fd_sc_hs__conb_1_231/HI sky130_fd_sc_hs__conb_1_231/a_165_290# sky130_fd_sc_hs__conb_1_231/a_21_290#
+ sky130_fd_sc_hs__conb_1
Xsky130_fd_sc_hs__conb_1_241 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__conb_1_241/LO
+ sky130_fd_sc_hs__conb_1_241/HI sky130_fd_sc_hs__conb_1_241/a_165_290# sky130_fd_sc_hs__conb_1_241/a_21_290#
+ sky130_fd_sc_hs__conb_1
Xsky130_fd_sc_hs__conb_1_252 DVSS: DVDD: DVDD: DVSS: prbs_generator_syn_27/eqn[30]
+ sky130_fd_sc_hs__conb_1_253/HI sky130_fd_sc_hs__conb_1_253/a_165_290# sky130_fd_sc_hs__conb_1_253/a_21_290#
+ sky130_fd_sc_hs__conb_1
Xsky130_fd_sc_hs__conb_1_263 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__conb_1_263/LO
+ sky130_fd_sc_hs__conb_1_263/HI sky130_fd_sc_hs__conb_1_263/a_165_290# sky130_fd_sc_hs__conb_1_263/a_21_290#
+ sky130_fd_sc_hs__conb_1
Xsky130_fd_sc_hs__clkbuf_8_11 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__clkbuf_8_11/X
+ sky130_fd_sc_hs__clkbuf_4_1/X sky130_fd_sc_hs__clkbuf_8_11/a_125_368# sky130_fd_sc_hs__clkbuf_8
Xsky130_fd_sc_hs__clkbuf_8_22 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__clkbuf_8_23/X
+ sky130_fd_sc_hs__clkbuf_8_23/A sky130_fd_sc_hs__clkbuf_8_23/a_125_368# sky130_fd_sc_hs__clkbuf_8
Xsky130_fd_sc_hs__clkbuf_8_33 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__nand2_2_11/B
+ sky130_fd_sc_hs__buf_2_77/X sky130_fd_sc_hs__clkbuf_8_33/a_125_368# sky130_fd_sc_hs__clkbuf_8
Xsky130_fd_sc_hs__clkbuf_8_44 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__clkbuf_2_3/A
+ sky130_fd_sc_hs__nand2_2_27/Y sky130_fd_sc_hs__clkbuf_8_45/a_125_368# sky130_fd_sc_hs__clkbuf_8
Xsky130_fd_sc_hs__clkbuf_8_55 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__inv_4_29/A
+ sky130_fd_sc_hs__or4_2_1/X sky130_fd_sc_hs__clkbuf_8_55/a_125_368# sky130_fd_sc_hs__clkbuf_8
Xsky130_fd_sc_hs__clkbuf_8_66 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__or4_2_1/B sky130_fd_sc_hs__clkbuf_8_67/A
+ sky130_fd_sc_hs__clkbuf_8_67/a_125_368# sky130_fd_sc_hs__clkbuf_8
Xsky130_fd_sc_hs__clkbuf_8_77 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__clkbuf_8_77/X
+ sky130_fd_sc_hs__clkbuf_8_77/A sky130_fd_sc_hs__clkbuf_8_77/a_125_368# sky130_fd_sc_hs__clkbuf_8
Xsky130_fd_sc_hs__clkbuf_8_88 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__einvp_8_7/TE
+ test_mux_select[3] sky130_fd_sc_hs__clkbuf_8_89/a_125_368# sky130_fd_sc_hs__clkbuf_8
Xsky130_fd_sc_hs__clkbuf_8_99 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__clkbuf_8_99/X
+ CTL_BUF_N[0] sky130_fd_sc_hs__clkbuf_8_99/a_125_368# sky130_fd_sc_hs__clkbuf_8
Xsky130_fd_sc_hs__nor2_4_3 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__nor2_4_3/Y sky130_fd_sc_hs__nor2_4_3/A
+ sky130_fd_sc_hs__nor2_4_3/B sky130_fd_sc_hs__nor2_4_3/a_27_368# sky130_fd_sc_hs__nor2_4
Xsky130_fd_sc_hs__einvp_8_8 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__inv_4_39/A sky130_fd_sc_hs__einvp_8_9/TE
+ fine_freq_track_1/out_star sky130_fd_sc_hs__einvp_8_9/a_802_323# sky130_fd_sc_hs__einvp_8_9/a_27_74#
+ sky130_fd_sc_hs__einvp_8_9/a_27_368# sky130_fd_sc_hs__einvp_8
Xsky130_fd_sc_hs__nand2_2_4 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__nand2_2_5/Y sky130_fd_sc_hs__nand2_2_5/B
+ sky130_fd_sc_hs__inv_4_29/A sky130_fd_sc_hs__nand2_2_5/a_27_74# sky130_fd_sc_hs__nand2_2
Xsky130_fd_sc_hs__or2b_4_0 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__or2b_4_1/A sky130_fd_sc_hs__nor4_2_1/A
+ sky130_fd_sc_hs__or2b_4_1/X sky130_fd_sc_hs__or2b_4_1/a_676_48# sky130_fd_sc_hs__or2b_4_1/a_489_392#
+ sky130_fd_sc_hs__or2b_4_1/a_81_296# sky130_fd_sc_hs__or2b_4
Xsky130_fd_sc_hs__clkbuf_4_5 DVSS: DVDD: DVDD: DVSS: pi3_con[2] sky130_fd_sc_hs__clkbuf_8_7/A
+ sky130_fd_sc_hs__clkbuf_4_5/a_83_270# sky130_fd_sc_hs__clkbuf_4
Xsky130_fd_sc_hs__einvp_2_60 DVSS: DVDD: DVDD: DVSS: dout_p sky130_fd_sc_hs__einvp_2_97/A
+ sky130_fd_sc_hs__dlrtp_1_51/Q sky130_fd_sc_hs__einvp_2_61/a_263_323# sky130_fd_sc_hs__einvp_2_61/a_36_74#
+ sky130_fd_sc_hs__einvp_2_61/a_27_368# sky130_fd_sc_hs__einvp_2
Xsky130_fd_sc_hs__einvp_2_71 DVSS: DVDD: DVDD: DVSS: dout_p sky130_fd_sc_hs__einvp_2_97/A
+ sky130_fd_sc_hs__dlrtp_1_58/Q sky130_fd_sc_hs__einvp_2_71/a_263_323# sky130_fd_sc_hs__einvp_2_71/a_36_74#
+ sky130_fd_sc_hs__einvp_2_71/a_27_368# sky130_fd_sc_hs__einvp_2
Xsky130_fd_sc_hs__einvp_2_82 DVSS: DVDD: DVDD: DVSS: dout_p sky130_fd_sc_hs__einvp_2_99/A
+ sky130_fd_sc_hs__buf_2_31/X sky130_fd_sc_hs__einvp_2_83/a_263_323# sky130_fd_sc_hs__einvp_2_83/a_36_74#
+ sky130_fd_sc_hs__einvp_2_83/a_27_368# sky130_fd_sc_hs__einvp_2
Xsky130_fd_sc_hs__einvp_2_93 DVSS: DVDD: DVDD: DVSS: dout_p sky130_fd_sc_hs__einvp_2_97/A
+ sky130_fd_sc_hs__dlrtp_1_77/Q sky130_fd_sc_hs__einvp_2_93/a_263_323# sky130_fd_sc_hs__einvp_2_93/a_36_74#
+ sky130_fd_sc_hs__einvp_2_93/a_27_368# sky130_fd_sc_hs__einvp_2
Xsky130_fd_sc_hs__clkinv_4_5 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__clkinv_4_5/Y
+ sky130_fd_sc_hs__nor4_2_1/A sky130_fd_sc_hs__clkinv_4
Xsky130_fd_sc_hs__conb_1_70 DVSS: DVDD: DVDD: DVSS: prbs_generator_syn_7/eqn[31] prbs_generator_syn_7/cke
+ sky130_fd_sc_hs__conb_1_71/a_165_290# sky130_fd_sc_hs__conb_1_71/a_21_290# sky130_fd_sc_hs__conb_1
Xsky130_fd_sc_hs__conb_1_81 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__conb_1_81/LO
+ prbs_generator_syn_11/cke sky130_fd_sc_hs__conb_1_81/a_165_290# sky130_fd_sc_hs__conb_1_81/a_21_290#
+ sky130_fd_sc_hs__conb_1
Xsky130_fd_sc_hs__conb_1_92 DVSS: DVDD: DVDD: DVSS: qr_4t1_mux_top_1/din_3_dummy sky130_fd_sc_hs__conb_1_93/HI
+ sky130_fd_sc_hs__conb_1_93/a_165_290# sky130_fd_sc_hs__conb_1_93/a_21_290# sky130_fd_sc_hs__conb_1
Xsky130_fd_sc_hs__dlrtp_1_104 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__dlrtp_1_105/Q
+ sky130_fd_sc_hs__dlrtp_1_9/GATE sky130_fd_sc_hs__conb_1_133/HI sky130_fd_sc_hs__o21bai_2_31/Y
+ sky130_fd_sc_hs__dlrtp_1_105/a_216_424# sky130_fd_sc_hs__dlrtp_1_105/a_759_508#
+ sky130_fd_sc_hs__dlrtp_1_105/a_565_74# sky130_fd_sc_hs__dlrtp_1_105/a_27_424# sky130_fd_sc_hs__dlrtp_1_105/a_1045_74#
+ sky130_fd_sc_hs__dlrtp_1_105/a_643_74# sky130_fd_sc_hs__dlrtp_1_105/a_817_48# sky130_fd_sc_hs__dlrtp_1_105/a_568_392#
+ sky130_fd_sc_hs__dlrtp_1_105/a_363_74# sky130_fd_sc_hs__dlrtp_1_105/a_769_74# sky130_fd_sc_hs__dlrtp_1
Xsky130_fd_sc_hs__dlrtp_1_115 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__buf_2_125/A
+ sky130_fd_sc_hs__dlrtp_1_9/GATE sky130_fd_sc_hs__conb_1_131/HI sky130_fd_sc_hs__dlrtp_1_115/D
+ sky130_fd_sc_hs__dlrtp_1_115/a_216_424# sky130_fd_sc_hs__dlrtp_1_115/a_759_508#
+ sky130_fd_sc_hs__dlrtp_1_115/a_565_74# sky130_fd_sc_hs__dlrtp_1_115/a_27_424# sky130_fd_sc_hs__dlrtp_1_115/a_1045_74#
+ sky130_fd_sc_hs__dlrtp_1_115/a_643_74# sky130_fd_sc_hs__dlrtp_1_115/a_817_48# sky130_fd_sc_hs__dlrtp_1_115/a_568_392#
+ sky130_fd_sc_hs__dlrtp_1_115/a_363_74# sky130_fd_sc_hs__dlrtp_1_115/a_769_74# sky130_fd_sc_hs__dlrtp_1
Xsky130_fd_sc_hs__dlrtp_1_126 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__dlrtp_1_127/Q
+ sky130_fd_sc_hs__clkbuf_2_3/A sky130_fd_sc_hs__conb_1_135/HI sky130_fd_sc_hs__buf_2_139/X
+ sky130_fd_sc_hs__dlrtp_1_127/a_216_424# sky130_fd_sc_hs__dlrtp_1_127/a_759_508#
+ sky130_fd_sc_hs__dlrtp_1_127/a_565_74# sky130_fd_sc_hs__dlrtp_1_127/a_27_424# sky130_fd_sc_hs__dlrtp_1_127/a_1045_74#
+ sky130_fd_sc_hs__dlrtp_1_127/a_643_74# sky130_fd_sc_hs__dlrtp_1_127/a_817_48# sky130_fd_sc_hs__dlrtp_1_127/a_568_392#
+ sky130_fd_sc_hs__dlrtp_1_127/a_363_74# sky130_fd_sc_hs__dlrtp_1_127/a_769_74# sky130_fd_sc_hs__dlrtp_1
Xsky130_fd_sc_hs__dlrtp_1_137 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__dlrtp_1_137/Q
+ sky130_fd_sc_hs__clkbuf_16_53/X sky130_fd_sc_hs__conb_1_135/HI sky130_fd_sc_hs__buf_2_145/X
+ sky130_fd_sc_hs__dlrtp_1_137/a_216_424# sky130_fd_sc_hs__dlrtp_1_137/a_759_508#
+ sky130_fd_sc_hs__dlrtp_1_137/a_565_74# sky130_fd_sc_hs__dlrtp_1_137/a_27_424# sky130_fd_sc_hs__dlrtp_1_137/a_1045_74#
+ sky130_fd_sc_hs__dlrtp_1_137/a_643_74# sky130_fd_sc_hs__dlrtp_1_137/a_817_48# sky130_fd_sc_hs__dlrtp_1_137/a_568_392#
+ sky130_fd_sc_hs__dlrtp_1_137/a_363_74# sky130_fd_sc_hs__dlrtp_1_137/a_769_74# sky130_fd_sc_hs__dlrtp_1
Xsky130_fd_sc_hs__dlrtp_1_148 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__dlrtp_1_149/Q
+ sky130_fd_sc_hs__clkbuf_16_53/X sky130_fd_sc_hs__conb_1_127/HI sky130_fd_sc_hs__buf_2_157/X
+ sky130_fd_sc_hs__dlrtp_1_149/a_216_424# sky130_fd_sc_hs__dlrtp_1_149/a_759_508#
+ sky130_fd_sc_hs__dlrtp_1_149/a_565_74# sky130_fd_sc_hs__dlrtp_1_149/a_27_424# sky130_fd_sc_hs__dlrtp_1_149/a_1045_74#
+ sky130_fd_sc_hs__dlrtp_1_149/a_643_74# sky130_fd_sc_hs__dlrtp_1_149/a_817_48# sky130_fd_sc_hs__dlrtp_1_149/a_568_392#
+ sky130_fd_sc_hs__dlrtp_1_149/a_363_74# sky130_fd_sc_hs__dlrtp_1_149/a_769_74# sky130_fd_sc_hs__dlrtp_1
Xsky130_fd_sc_hs__dlrtp_1_159 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__buf_2_161/A
+ sky130_fd_sc_hs__clkbuf_16_53/X sky130_fd_sc_hs__conb_1_137/HI sky130_fd_sc_hs__buf_2_75/X
+ sky130_fd_sc_hs__dlrtp_1_159/a_216_424# sky130_fd_sc_hs__dlrtp_1_159/a_759_508#
+ sky130_fd_sc_hs__dlrtp_1_159/a_565_74# sky130_fd_sc_hs__dlrtp_1_159/a_27_424# sky130_fd_sc_hs__dlrtp_1_159/a_1045_74#
+ sky130_fd_sc_hs__dlrtp_1_159/a_643_74# sky130_fd_sc_hs__dlrtp_1_159/a_817_48# sky130_fd_sc_hs__dlrtp_1_159/a_568_392#
+ sky130_fd_sc_hs__dlrtp_1_159/a_363_74# sky130_fd_sc_hs__dlrtp_1_159/a_769_74# sky130_fd_sc_hs__dlrtp_1
Xsky130_fd_sc_hs__inv_4_7 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__inv_4_7/Y fine_control_avg_window_select[1]
+ sky130_fd_sc_hs__inv_4
Xsky130_fd_sc_hs__dlrtp_1_50 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__dlrtp_1_51/Q
+ sky130_fd_sc_hs__clkbuf_16_53/A sky130_fd_sc_hs__conb_1_123/HI sky130_fd_sc_hs__inv_4_11/A
+ sky130_fd_sc_hs__dlrtp_1_51/a_216_424# sky130_fd_sc_hs__dlrtp_1_51/a_759_508# sky130_fd_sc_hs__dlrtp_1_51/a_565_74#
+ sky130_fd_sc_hs__dlrtp_1_51/a_27_424# sky130_fd_sc_hs__dlrtp_1_51/a_1045_74# sky130_fd_sc_hs__dlrtp_1_51/a_643_74#
+ sky130_fd_sc_hs__dlrtp_1_51/a_817_48# sky130_fd_sc_hs__dlrtp_1_51/a_568_392# sky130_fd_sc_hs__dlrtp_1_51/a_363_74#
+ sky130_fd_sc_hs__dlrtp_1_51/a_769_74# sky130_fd_sc_hs__dlrtp_1
Xsky130_fd_sc_hs__dlrtp_1_61 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__buf_2_31/A sky130_fd_sc_hs__clkbuf_16_53/A
+ sky130_fd_sc_hs__conb_1_125/HI sky130_fd_sc_hs__buf_2_59/X sky130_fd_sc_hs__dlrtp_1_61/a_216_424#
+ sky130_fd_sc_hs__dlrtp_1_61/a_759_508# sky130_fd_sc_hs__dlrtp_1_61/a_565_74# sky130_fd_sc_hs__dlrtp_1_61/a_27_424#
+ sky130_fd_sc_hs__dlrtp_1_61/a_1045_74# sky130_fd_sc_hs__dlrtp_1_61/a_643_74# sky130_fd_sc_hs__dlrtp_1_61/a_817_48#
+ sky130_fd_sc_hs__dlrtp_1_61/a_568_392# sky130_fd_sc_hs__dlrtp_1_61/a_363_74# sky130_fd_sc_hs__dlrtp_1_61/a_769_74#
+ sky130_fd_sc_hs__dlrtp_1
Xsky130_fd_sc_hs__dlrtp_1_72 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__dlrtp_1_74/Q
+ sky130_fd_sc_hs__clkbuf_16_53/X sky130_fd_sc_hs__conb_1_129/HI sky130_fd_sc_hs__dlrtp_1_74/D
+ sky130_fd_sc_hs__dlrtp_1_74/a_216_424# sky130_fd_sc_hs__dlrtp_1_74/a_759_508# sky130_fd_sc_hs__dlrtp_1_74/a_565_74#
+ sky130_fd_sc_hs__dlrtp_1_74/a_27_424# sky130_fd_sc_hs__dlrtp_1_74/a_1045_74# sky130_fd_sc_hs__dlrtp_1_74/a_643_74#
+ sky130_fd_sc_hs__dlrtp_1_74/a_817_48# sky130_fd_sc_hs__dlrtp_1_74/a_568_392# sky130_fd_sc_hs__dlrtp_1_74/a_363_74#
+ sky130_fd_sc_hs__dlrtp_1_74/a_769_74# sky130_fd_sc_hs__dlrtp_1
Xsky130_fd_sc_hs__dlrtp_1_83 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__buf_2_63/A sky130_fd_sc_hs__clkbuf_16_53/X
+ sky130_fd_sc_hs__conb_1_137/HI sky130_fd_sc_hs__o21ai_2_17/Y sky130_fd_sc_hs__dlrtp_1_83/a_216_424#
+ sky130_fd_sc_hs__dlrtp_1_83/a_759_508# sky130_fd_sc_hs__dlrtp_1_83/a_565_74# sky130_fd_sc_hs__dlrtp_1_83/a_27_424#
+ sky130_fd_sc_hs__dlrtp_1_83/a_1045_74# sky130_fd_sc_hs__dlrtp_1_83/a_643_74# sky130_fd_sc_hs__dlrtp_1_83/a_817_48#
+ sky130_fd_sc_hs__dlrtp_1_83/a_568_392# sky130_fd_sc_hs__dlrtp_1_83/a_363_74# sky130_fd_sc_hs__dlrtp_1_83/a_769_74#
+ sky130_fd_sc_hs__dlrtp_1
Xsky130_fd_sc_hs__dlrtp_1_94 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__dlrtp_1_95/Q
+ sky130_fd_sc_hs__dlrtp_1_9/GATE sky130_fd_sc_hs__conb_1_133/HI sky130_fd_sc_hs__buf_2_101/X
+ sky130_fd_sc_hs__dlrtp_1_95/a_216_424# sky130_fd_sc_hs__dlrtp_1_95/a_759_508# sky130_fd_sc_hs__dlrtp_1_95/a_565_74#
+ sky130_fd_sc_hs__dlrtp_1_95/a_27_424# sky130_fd_sc_hs__dlrtp_1_95/a_1045_74# sky130_fd_sc_hs__dlrtp_1_95/a_643_74#
+ sky130_fd_sc_hs__dlrtp_1_95/a_817_48# sky130_fd_sc_hs__dlrtp_1_95/a_568_392# sky130_fd_sc_hs__dlrtp_1_95/a_363_74#
+ sky130_fd_sc_hs__dlrtp_1_95/a_769_74# sky130_fd_sc_hs__dlrtp_1
Xsky130_fd_sc_hs__clkbuf_2_2 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__clkbuf_2_3/X
+ sky130_fd_sc_hs__clkbuf_2_3/A sky130_fd_sc_hs__clkbuf_2_3/a_43_192# sky130_fd_sc_hs__clkbuf_2
Xsky130_fd_sc_hs__clkbuf_2_13 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__dlrtp_1_71/D
+ sky130_fd_sc_hs__o21bai_2_13/Y sky130_fd_sc_hs__clkbuf_2_13/a_43_192# sky130_fd_sc_hs__clkbuf_2
Xsky130_fd_sc_hs__clkbuf_2_24 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__dlrtp_1_89/D
+ sky130_fd_sc_hs__o21ai_2_21/Y sky130_fd_sc_hs__clkbuf_2_25/a_43_192# sky130_fd_sc_hs__clkbuf_2
Xsky130_fd_sc_hs__clkbuf_2_35 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__dlrtp_1_103/D
+ sky130_fd_sc_hs__o21ai_4_1/Y sky130_fd_sc_hs__clkbuf_2_35/a_43_192# sky130_fd_sc_hs__clkbuf_2
Xsky130_fd_sc_hs__clkbuf_2_46 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__dlrtp_1_17/D
+ sky130_fd_sc_hs__o21bai_2_41/Y sky130_fd_sc_hs__clkbuf_2_47/a_43_192# sky130_fd_sc_hs__clkbuf_2
Xsky130_fd_sc_hs__clkbuf_2_57 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__buf_2_131/A
+ sky130_fd_sc_hs__nor4_2_1/Y sky130_fd_sc_hs__clkbuf_2_57/a_43_192# sky130_fd_sc_hs__clkbuf_2
Xsky130_fd_sc_hs__clkbuf_2_68 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__dlrtp_1_153/D
+ sky130_fd_sc_hs__o21bai_2_67/Y sky130_fd_sc_hs__clkbuf_2_69/a_43_192# sky130_fd_sc_hs__clkbuf_2
Xsky130_fd_sc_hs__clkinv_2_2 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__clkinv_2_3/Y
+ sky130_fd_sc_hs__inv_4_7/Y sky130_fd_sc_hs__clkinv_2
Xsky130_fd_sc_hs__buf_2_4 DVSS: DVDD: DVDD: DVSS: manual_control_osc[8] sky130_fd_sc_hs__buf_2_5/X
+ sky130_fd_sc_hs__buf_2_5/a_21_260# sky130_fd_sc_hs__buf_2
Xsky130_fd_sc_hs__dlrtp_1_6 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__dlrtp_1_7/Q sky130_fd_sc_hs__dlrtp_1_9/GATE
+ sky130_fd_sc_hs__conb_1_117/HI sky130_fd_sc_hs__inv_4_21/A sky130_fd_sc_hs__dlrtp_1_7/a_216_424#
+ sky130_fd_sc_hs__dlrtp_1_7/a_759_508# sky130_fd_sc_hs__dlrtp_1_7/a_565_74# sky130_fd_sc_hs__dlrtp_1_7/a_27_424#
+ sky130_fd_sc_hs__dlrtp_1_7/a_1045_74# sky130_fd_sc_hs__dlrtp_1_7/a_643_74# sky130_fd_sc_hs__dlrtp_1_7/a_817_48#
+ sky130_fd_sc_hs__dlrtp_1_7/a_568_392# sky130_fd_sc_hs__dlrtp_1_7/a_363_74# sky130_fd_sc_hs__dlrtp_1_7/a_769_74#
+ sky130_fd_sc_hs__dlrtp_1
Xsky130_fd_sc_hs__buf_2_20 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__buf_2_25/X sky130_fd_sc_hs__buf_2_21/X
+ sky130_fd_sc_hs__buf_2_21/a_21_260# sky130_fd_sc_hs__buf_2
Xsky130_fd_sc_hs__buf_2_31 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__buf_2_31/A sky130_fd_sc_hs__buf_2_31/X
+ sky130_fd_sc_hs__buf_2_31/a_21_260# sky130_fd_sc_hs__buf_2
Xsky130_fd_sc_hs__buf_2_42 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__buf_2_43/A sky130_fd_sc_hs__buf_2_55/A
+ sky130_fd_sc_hs__buf_2_43/a_21_260# sky130_fd_sc_hs__buf_2
Xsky130_fd_sc_hs__buf_2_53 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__buf_2_61/X sky130_fd_sc_hs__buf_2_53/X
+ sky130_fd_sc_hs__buf_2_53/a_21_260# sky130_fd_sc_hs__buf_2
Xsky130_fd_sc_hs__buf_2_64 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__inv_4_11/Y sky130_fd_sc_hs__buf_2_65/X
+ sky130_fd_sc_hs__buf_2_65/a_21_260# sky130_fd_sc_hs__buf_2
Xsky130_fd_sc_hs__buf_2_75 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__buf_2_75/A sky130_fd_sc_hs__buf_2_75/X
+ sky130_fd_sc_hs__buf_2_75/a_21_260# sky130_fd_sc_hs__buf_2
Xsky130_fd_sc_hs__buf_2_86 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__buf_2_87/A sky130_fd_sc_hs__inv_4_19/A
+ sky130_fd_sc_hs__buf_2_87/a_21_260# sky130_fd_sc_hs__buf_2
Xsky130_fd_sc_hs__buf_2_97 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__buf_2_99/A sky130_fd_sc_hs__buf_2_99/X
+ sky130_fd_sc_hs__buf_2_99/a_21_260# sky130_fd_sc_hs__buf_2
Xsky130_fd_sc_hs__o21bai_2_11 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__inv_8_1/Y sky130_fd_sc_hs__nand2_2_11/B
+ sky130_fd_sc_hs__dlrtp_1_69/D sky130_fd_sc_hs__buf_2_61/A sky130_fd_sc_hs__o21bai_2_11/a_27_74#
+ sky130_fd_sc_hs__o21bai_2_11/a_225_74# sky130_fd_sc_hs__o21bai_2_11/a_507_368# sky130_fd_sc_hs__o21bai_2
Xsky130_fd_sc_hs__o21bai_2_22 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__clkinv_4_3/Y
+ sky130_fd_sc_hs__buf_8_3/X sky130_fd_sc_hs__buf_2_101/X sky130_fd_sc_hs__buf_2_103/A
+ sky130_fd_sc_hs__o21bai_2_23/a_27_74# sky130_fd_sc_hs__o21bai_2_23/a_225_74# sky130_fd_sc_hs__o21bai_2_23/a_507_368#
+ sky130_fd_sc_hs__o21bai_2
Xsky130_fd_sc_hs__o21bai_2_33 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__clkinv_4_3/Y
+ sky130_fd_sc_hs__or2b_2_3/A sky130_fd_sc_hs__dlrtp_1_99/D sky130_fd_sc_hs__buf_2_111/A
+ sky130_fd_sc_hs__o21bai_2_33/a_27_74# sky130_fd_sc_hs__o21bai_2_33/a_225_74# sky130_fd_sc_hs__o21bai_2_33/a_507_368#
+ sky130_fd_sc_hs__o21bai_2
Xsky130_fd_sc_hs__o21bai_2_44 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__clkinv_4_5/Y
+ sky130_fd_sc_hs__nand2_2_15/B sky130_fd_sc_hs__buf_2_121/X sky130_fd_sc_hs__buf_2_117/A
+ sky130_fd_sc_hs__o21bai_2_45/a_27_74# sky130_fd_sc_hs__o21bai_2_45/a_225_74# sky130_fd_sc_hs__o21bai_2_45/a_507_368#
+ sky130_fd_sc_hs__o21bai_2
Xsky130_fd_sc_hs__o21bai_2_55 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__o21bai_4_3/A2
+ sky130_fd_sc_hs__nand2_2_21/B sky130_fd_sc_hs__dlrtp_1_35/D sky130_fd_sc_hs__buf_2_133/A
+ sky130_fd_sc_hs__o21bai_2_55/a_27_74# sky130_fd_sc_hs__o21bai_2_55/a_225_74# sky130_fd_sc_hs__o21bai_2_55/a_507_368#
+ sky130_fd_sc_hs__o21bai_2
Xsky130_fd_sc_hs__o21bai_2_66 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__nand2_2_9/B
+ sky130_fd_sc_hs__o21bai_4_7/A1 sky130_fd_sc_hs__buf_2_47/X sky130_fd_sc_hs__dlrtp_1_74/D
+ sky130_fd_sc_hs__o21bai_2_66/a_27_74# sky130_fd_sc_hs__o21bai_2_66/a_225_74# sky130_fd_sc_hs__o21bai_2_66/a_507_368#
+ sky130_fd_sc_hs__o21bai_2
Xsky130_fd_sc_hs__o21bai_4_0 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__buf_2_30/A sky130_fd_sc_hs__inv_8_1/Y
+ sky130_fd_sc_hs__nand2_2_3/B sky130_fd_sc_hs__buf_2_49/X sky130_fd_sc_hs__o21bai_4_1/a_28_368#
+ sky130_fd_sc_hs__o21bai_4_1/a_27_74# sky130_fd_sc_hs__o21bai_4_1/a_828_48# sky130_fd_sc_hs__o21bai_4
Xsky130_fd_sc_hs__conb_1_220 DVSS: DVDD: DVDD: DVSS: prbs_generator_syn_25/eqn[31]
+ prbs_generator_syn_25/cke sky130_fd_sc_hs__conb_1_221/a_165_290# sky130_fd_sc_hs__conb_1_221/a_21_290#
+ sky130_fd_sc_hs__conb_1
Xsky130_fd_sc_hs__conb_1_231 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__conb_1_231/LO
+ sky130_fd_sc_hs__conb_1_231/HI sky130_fd_sc_hs__conb_1_231/a_165_290# sky130_fd_sc_hs__conb_1_231/a_21_290#
+ sky130_fd_sc_hs__conb_1
Xsky130_fd_sc_hs__conb_1_242 DVSS: DVDD: DVDD: DVSS: prbs_generator_syn_31/eqn[9]
+ sky130_fd_sc_hs__conb_1_243/HI sky130_fd_sc_hs__conb_1_243/a_165_290# sky130_fd_sc_hs__conb_1_243/a_21_290#
+ sky130_fd_sc_hs__conb_1
Xsky130_fd_sc_hs__conb_1_253 DVSS: DVDD: DVDD: DVSS: prbs_generator_syn_27/eqn[30]
+ sky130_fd_sc_hs__conb_1_253/HI sky130_fd_sc_hs__conb_1_253/a_165_290# sky130_fd_sc_hs__conb_1_253/a_21_290#
+ sky130_fd_sc_hs__conb_1
Xsky130_fd_sc_hs__conb_1_264 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__conb_1_265/LO
+ sky130_fd_sc_hs__conb_1_265/HI sky130_fd_sc_hs__conb_1_265/a_165_290# sky130_fd_sc_hs__conb_1_265/a_21_290#
+ sky130_fd_sc_hs__conb_1
Xsky130_fd_sc_hs__clkbuf_8_12 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__clkbuf_8_13/X
+ sky130_fd_sc_hs__clkbuf_8_13/A sky130_fd_sc_hs__clkbuf_8_13/a_125_368# sky130_fd_sc_hs__clkbuf_8
Xsky130_fd_sc_hs__clkbuf_8_23 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__clkbuf_8_23/X
+ sky130_fd_sc_hs__clkbuf_8_23/A sky130_fd_sc_hs__clkbuf_8_23/a_125_368# sky130_fd_sc_hs__clkbuf_8
Xsky130_fd_sc_hs__clkbuf_8_34 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__clkbuf_8_35/X
+ sky130_fd_sc_hs__clkbuf_8_35/A sky130_fd_sc_hs__clkbuf_8_35/a_125_368# sky130_fd_sc_hs__clkbuf_8
Xsky130_fd_sc_hs__clkbuf_8_45 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__clkbuf_2_3/A
+ sky130_fd_sc_hs__nand2_2_27/Y sky130_fd_sc_hs__clkbuf_8_45/a_125_368# sky130_fd_sc_hs__clkbuf_8
Xsky130_fd_sc_hs__clkbuf_8_56 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__o21bai_2_3/A2
+ sky130_fd_sc_hs__nand2_2_33/Y sky130_fd_sc_hs__clkbuf_8_57/a_125_368# sky130_fd_sc_hs__clkbuf_8
Xsky130_fd_sc_hs__clkbuf_8_67 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__or4_2_1/B sky130_fd_sc_hs__clkbuf_8_67/A
+ sky130_fd_sc_hs__clkbuf_8_67/a_125_368# sky130_fd_sc_hs__clkbuf_8
Xsky130_fd_sc_hs__clkbuf_8_78 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__clkbuf_8_79/X
+ sky130_fd_sc_hs__clkbuf_8_79/A sky130_fd_sc_hs__clkbuf_8_79/a_125_368# sky130_fd_sc_hs__clkbuf_8
Xsky130_fd_sc_hs__clkbuf_8_89 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__einvp_8_7/TE
+ test_mux_select[3] sky130_fd_sc_hs__clkbuf_8_89/a_125_368# sky130_fd_sc_hs__clkbuf_8
Xsky130_fd_sc_hs__einvp_8_9 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__inv_4_39/A sky130_fd_sc_hs__einvp_8_9/TE
+ fine_freq_track_1/out_star sky130_fd_sc_hs__einvp_8_9/a_802_323# sky130_fd_sc_hs__einvp_8_9/a_27_74#
+ sky130_fd_sc_hs__einvp_8_9/a_27_368# sky130_fd_sc_hs__einvp_8
Xsky130_fd_sc_hs__nand2_2_5 DVSS: DVDD: DVDD: DVSS: sky130_fd_sc_hs__nand2_2_5/Y sky130_fd_sc_hs__nand2_2_5/B
+ sky130_fd_sc_hs__inv_4_29/A sky130_fd_sc_hs__nand2_2_5/a_27_74# sky130_fd_sc_hs__nand2_2
.ends

